magic
tech sky130A
magscale 1 2
timestamp 1757045633
<< nwell >>
rect 14815 19209 17501 19733
rect 8225 17041 8749 18633
rect 9012 16642 9868 18636
rect 10125 16111 10981 18633
rect 15445 16111 16301 18633
rect 16558 17248 17082 18630
rect 17345 17041 17869 18633
rect 10398 11580 13128 11860
rect 13428 11580 16158 11860
rect 19298 11490 22738 12800
rect 22995 11913 23519 13323
rect 11498 10020 15058 10700
rect 15358 10220 16128 10500
rect 11508 9420 13148 9700
rect 13408 9420 15048 9700
rect 22995 9449 23519 10803
rect 13128 6470 18108 7710
rect 19388 6500 22608 7080
rect 12318 3390 22768 3600
rect 23048 3340 25358 5570
<< pwell >>
rect 13238 18810 13318 19090
rect 11248 18657 12588 18810
rect 11248 17623 11401 18657
rect 12435 17623 12588 18657
rect 11248 17470 12588 17623
rect 12608 18657 13948 18810
rect 12608 17623 12761 18657
rect 13795 17623 13948 18657
rect 12608 17470 13948 17623
rect 13968 18657 15308 18810
rect 13968 17623 14121 18657
rect 15155 17623 15308 18657
rect 13968 17470 15308 17623
rect 11248 17297 12588 17450
rect 11248 16263 11401 17297
rect 12435 16263 12588 17297
rect 11248 16110 12588 16263
rect 12608 17297 13948 17450
rect 12608 16263 12761 17297
rect 13795 16263 13948 17297
rect 12608 16110 13948 16263
rect 13968 17297 15308 17450
rect 13968 16263 14121 17297
rect 15155 16263 15308 17297
rect 13968 16110 15308 16263
rect 11248 15937 12588 16090
rect 11248 14903 11401 15937
rect 12435 14903 12588 15937
rect 11248 14750 12588 14903
rect 12608 15937 13948 16090
rect 12608 14903 12761 15937
rect 13795 14903 13948 15937
rect 12608 14750 13948 14903
rect 13968 15937 15308 16090
rect 13968 14903 14121 15937
rect 15155 14903 15308 15937
rect 13968 14750 15308 14903
rect 23048 1840 25168 3260
<< nbase >>
rect 11401 17623 12435 18657
rect 12761 17623 13795 18657
rect 14121 17623 15155 18657
rect 11401 16263 12435 17297
rect 12761 16263 13795 17297
rect 14121 16263 15155 17297
rect 11401 14903 12435 15937
rect 12761 14903 13795 15937
rect 14121 14903 15155 15937
<< nmos >>
rect 11238 14080 13238 14280
rect 13318 14080 15318 14280
rect 10818 13170 11818 13670
rect 12058 13170 13058 13670
rect 13498 13170 14498 13670
rect 14738 13170 15738 13670
rect 11438 12560 11478 12660
rect 11558 12560 11598 12660
rect 11678 12560 11718 12660
rect 11798 12560 11838 12660
rect 11918 12560 11958 12660
rect 12038 12560 12078 12660
rect 12158 12560 12198 12660
rect 12278 12560 12318 12660
rect 12398 12560 12438 12660
rect 12518 12560 12558 12660
rect 13998 12560 14038 12660
rect 14118 12560 14158 12660
rect 14238 12560 14278 12660
rect 14358 12560 14398 12660
rect 14478 12560 14518 12660
rect 14598 12560 14638 12660
rect 14718 12560 14758 12660
rect 14838 12560 14878 12660
rect 14958 12560 14998 12660
rect 15078 12560 15118 12660
rect 19538 10960 19568 11060
rect 19668 10960 19698 11060
rect 19798 10960 19828 11060
rect 19928 10960 19958 11060
rect 20058 10960 20088 11060
rect 20188 10960 20218 11060
rect 20678 10960 20708 11060
rect 20808 10960 20838 11060
rect 20938 10960 20968 11060
rect 21068 10960 21098 11060
rect 21198 10960 21228 11060
rect 21328 10960 21358 11060
rect 21818 10960 21848 11060
rect 21948 10960 21978 11060
rect 22078 10960 22108 11060
rect 22208 10960 22238 11060
rect 22338 10960 22368 11060
rect 22468 10960 22498 11060
rect 19488 10270 19588 10520
rect 19688 10270 19788 10520
rect 19888 10270 19988 10520
rect 20088 10270 20188 10520
rect 20288 10270 20388 10520
rect 20488 10270 20588 10520
rect 20688 10270 20788 10520
rect 20888 10270 20988 10520
rect 21088 10270 21188 10520
rect 21288 10270 21388 10520
rect 13328 7890 13358 8090
rect 13438 7890 13468 8090
rect 13848 7890 13878 8090
rect 13958 7890 13988 8090
rect 14228 7890 14258 8090
rect 14338 7890 14368 8090
rect 14748 7890 14778 8090
rect 14858 7890 14888 8090
rect 15258 7890 15288 8090
rect 15588 7890 15618 8090
rect 15918 7890 15948 8090
rect 16478 7890 16508 8090
rect 16868 7890 16898 8090
rect 17258 7890 17288 8090
rect 17548 7890 17578 8090
rect 17938 7890 17968 8090
rect 19428 7640 19548 8040
rect 19648 7640 19768 8040
rect 19868 7640 19988 8040
rect 20088 7640 20208 8040
rect 20508 7640 20628 8040
rect 20728 7640 20848 8040
rect 20948 7640 21068 8040
rect 21168 7640 21288 8040
rect 21588 7640 21708 8040
rect 21808 7640 21928 8040
rect 22028 7640 22148 8040
rect 22248 7640 22368 8040
rect 13328 6090 13358 6290
rect 13438 6090 13468 6290
rect 13848 6090 13878 6290
rect 13958 6090 13988 6290
rect 14228 6090 14258 6290
rect 14338 6090 14368 6290
rect 14748 6090 14778 6290
rect 14858 6090 14888 6290
rect 15268 6090 15298 6290
rect 15378 6090 15408 6290
rect 15708 6090 15738 6290
rect 16038 6090 16068 6290
rect 16478 6090 16508 6290
rect 16868 6090 16898 6290
rect 17258 6090 17288 6290
rect 17548 6090 17578 6290
rect 12508 3110 12538 3210
rect 12618 3110 12648 3210
rect 12728 3110 12758 3210
rect 12838 3110 12868 3210
rect 13088 3110 13118 3210
rect 13198 3110 13228 3210
rect 13538 3110 13568 3210
rect 13648 3110 13678 3210
rect 13758 3110 13788 3210
rect 13868 3110 13898 3210
rect 14198 3110 14228 3210
rect 14308 3110 14338 3210
rect 14418 3110 14448 3210
rect 14528 3110 14558 3210
rect 14878 3110 14908 3210
rect 14988 3110 15018 3210
rect 15098 3110 15128 3210
rect 15208 3110 15238 3210
rect 15458 3110 15488 3210
rect 15568 3110 15598 3210
rect 16018 3110 16048 3210
rect 16378 3110 16408 3210
rect 16628 3110 16658 3210
rect 16738 3110 16768 3210
rect 16848 3110 16878 3210
rect 16958 3110 16988 3210
rect 17288 3110 17318 3210
rect 17398 3110 17428 3210
rect 17508 3110 17538 3210
rect 17838 3110 17868 3210
rect 17948 3110 17978 3210
rect 18058 3110 18088 3210
rect 18168 3110 18198 3210
rect 18498 3110 18528 3210
rect 18608 3110 18638 3210
rect 18718 3110 18748 3210
rect 19138 3020 19168 3120
rect 19248 3020 19278 3120
rect 19358 3020 19388 3120
rect 19468 3020 19498 3120
rect 19798 3020 19828 3120
rect 19908 3020 19938 3120
rect 20018 3020 20048 3120
rect 20438 3020 20468 3120
rect 20548 3020 20578 3120
rect 20658 3020 20688 3120
rect 20768 3020 20798 3120
rect 21098 3020 21128 3120
rect 21208 3020 21238 3120
rect 21318 3020 21348 3120
rect 21738 3020 21768 3120
rect 21848 3020 21878 3120
rect 21958 3020 21988 3120
rect 22068 3020 22098 3120
rect 22398 3020 22428 3120
rect 22508 3020 22538 3120
rect 22618 3020 22648 3120
rect 23276 2840 23308 3040
rect 23796 2840 23828 3040
rect 24316 2840 24348 3040
rect 23278 2360 23308 2660
rect 23798 2360 23828 2660
rect 24318 2360 24348 2660
rect 23278 1980 23308 2180
rect 23798 1980 23828 2180
rect 24318 1980 24348 2180
rect 24918 1980 24948 2180
<< pmos >>
rect 19608 12190 19708 12690
rect 19808 12190 19908 12690
rect 20008 12190 20108 12690
rect 20208 12190 20308 12690
rect 20408 12190 20508 12690
rect 20608 12190 20708 12690
rect 20808 12190 20908 12690
rect 21008 12190 21108 12690
rect 21208 12190 21308 12690
rect 21408 12190 21508 12690
rect 10598 11620 10638 11820
rect 10718 11620 10758 11820
rect 10838 11620 10878 11820
rect 10958 11620 10998 11820
rect 11078 11620 11118 11820
rect 11198 11620 11238 11820
rect 11318 11620 11358 11820
rect 11438 11620 11478 11820
rect 11558 11620 11598 11820
rect 11678 11620 11718 11820
rect 11798 11620 11838 11820
rect 11918 11620 11958 11820
rect 12038 11620 12078 11820
rect 12158 11620 12198 11820
rect 12278 11620 12318 11820
rect 12398 11620 12438 11820
rect 12518 11620 12558 11820
rect 12638 11620 12678 11820
rect 12758 11620 12798 11820
rect 12878 11620 12918 11820
rect 13638 11620 13678 11820
rect 13758 11620 13798 11820
rect 13878 11620 13918 11820
rect 13998 11620 14038 11820
rect 14118 11620 14158 11820
rect 14238 11620 14278 11820
rect 14358 11620 14398 11820
rect 14478 11620 14518 11820
rect 14598 11620 14638 11820
rect 14718 11620 14758 11820
rect 14838 11620 14878 11820
rect 14958 11620 14998 11820
rect 15078 11620 15118 11820
rect 15198 11620 15238 11820
rect 15318 11620 15358 11820
rect 15438 11620 15478 11820
rect 15558 11620 15598 11820
rect 15678 11620 15718 11820
rect 15798 11620 15838 11820
rect 15918 11620 15958 11820
rect 19538 11540 19568 11740
rect 19668 11540 19698 11740
rect 19798 11540 19828 11740
rect 19928 11540 19958 11740
rect 20058 11540 20088 11740
rect 20188 11540 20218 11740
rect 20678 11540 20708 11740
rect 20808 11540 20838 11740
rect 20938 11540 20968 11740
rect 21068 11540 21098 11740
rect 21198 11540 21228 11740
rect 21328 11540 21358 11740
rect 21818 11540 21848 11740
rect 21948 11540 21978 11740
rect 22078 11540 22108 11740
rect 22208 11540 22238 11740
rect 22338 11540 22368 11740
rect 22468 11540 22498 11740
rect 11698 10060 11798 10660
rect 11878 10060 11978 10660
rect 12058 10060 12158 10660
rect 12238 10060 12338 10660
rect 12418 10060 12518 10660
rect 12598 10060 12698 10660
rect 12778 10060 12878 10660
rect 12958 10060 13058 10660
rect 13138 10060 13238 10660
rect 13318 10060 13418 10660
rect 13498 10060 13598 10660
rect 13678 10060 13778 10660
rect 13858 10060 13958 10660
rect 14038 10060 14138 10660
rect 14218 10060 14318 10660
rect 14398 10060 14498 10660
rect 14578 10060 14678 10660
rect 14758 10060 14858 10660
rect 15568 10260 15598 10460
rect 15678 10260 15708 10460
rect 15788 10260 15818 10460
rect 15898 10260 15928 10460
rect 11708 9460 11738 9660
rect 11818 9460 11848 9660
rect 11928 9460 11958 9660
rect 12038 9460 12068 9660
rect 12148 9460 12178 9660
rect 12258 9460 12288 9660
rect 12368 9460 12398 9660
rect 12478 9460 12508 9660
rect 12588 9460 12618 9660
rect 12698 9460 12728 9660
rect 12808 9460 12838 9660
rect 12918 9460 12948 9660
rect 13608 9460 13638 9660
rect 13718 9460 13748 9660
rect 13828 9460 13858 9660
rect 13938 9460 13968 9660
rect 14048 9460 14078 9660
rect 14158 9460 14188 9660
rect 14268 9460 14298 9660
rect 14378 9460 14408 9660
rect 14488 9460 14518 9660
rect 14598 9460 14628 9660
rect 14708 9460 14738 9660
rect 14818 9460 14848 9660
rect 13328 7270 13358 7670
rect 13438 7270 13468 7670
rect 13848 7270 13878 7670
rect 13958 7270 13988 7670
rect 14228 7270 14258 7670
rect 14338 7270 14368 7670
rect 14748 7270 14778 7670
rect 14858 7270 14888 7670
rect 15258 7270 15288 7670
rect 15588 7270 15618 7670
rect 15918 7270 15948 7670
rect 16478 7270 16508 7670
rect 16868 7270 16898 7670
rect 17258 7270 17288 7670
rect 17548 7270 17578 7670
rect 13328 6510 13358 6910
rect 13438 6510 13468 6910
rect 13848 6510 13878 6910
rect 13958 6510 13988 6910
rect 14228 6510 14258 6910
rect 14338 6510 14368 6910
rect 14748 6510 14778 6910
rect 14858 6510 14888 6910
rect 15268 6510 15298 6910
rect 15378 6510 15408 6910
rect 15708 6510 15738 6910
rect 16038 6510 16068 6910
rect 16478 6510 16508 6910
rect 16868 6510 16898 6910
rect 17258 6510 17288 6910
rect 17548 6510 17578 6910
rect 17938 6510 17968 6910
rect 19628 6540 19748 6940
rect 19848 6540 19968 6940
rect 20068 6540 20188 6940
rect 20288 6540 20408 6940
rect 20508 6540 20628 6940
rect 20728 6540 20848 6940
rect 21148 6540 21268 6940
rect 21368 6540 21488 6940
rect 21588 6540 21708 6940
rect 21808 6540 21928 6940
rect 22028 6540 22148 6940
rect 22248 6540 22368 6940
rect 23278 5030 23578 5430
rect 23798 5030 24098 5430
rect 24318 5030 24618 5430
rect 24838 5030 25138 5430
rect 12668 3430 12698 3530
rect 13088 3430 13118 3530
rect 13198 3430 13228 3530
rect 13758 3430 13788 3530
rect 13868 3430 13898 3530
rect 14198 3430 14228 3530
rect 14308 3430 14338 3530
rect 14418 3430 14448 3530
rect 15038 3430 15068 3530
rect 15458 3430 15488 3530
rect 15568 3430 15598 3530
rect 15908 3430 15938 3530
rect 16018 3430 16048 3530
rect 16268 3430 16298 3530
rect 16378 3430 16408 3530
rect 16848 3430 16878 3530
rect 16958 3430 16988 3530
rect 17288 3430 17318 3530
rect 17398 3430 17428 3530
rect 17908 3430 17938 3530
rect 18248 3430 18278 3530
rect 18358 3430 18388 3530
rect 18608 3430 18638 3530
rect 18718 3430 18748 3530
rect 19208 3430 19238 3530
rect 19548 3430 19578 3530
rect 19658 3430 19688 3530
rect 19908 3430 19938 3530
rect 20018 3430 20048 3530
rect 20508 3430 20538 3530
rect 20848 3430 20878 3530
rect 20958 3430 20988 3530
rect 21208 3430 21238 3530
rect 21318 3430 21348 3530
rect 21808 3430 21838 3530
rect 22148 3430 22178 3530
rect 22258 3430 22288 3530
rect 22508 3430 22538 3530
rect 22618 3430 22648 3530
rect 23278 4140 23308 4740
rect 23798 4140 23828 4740
rect 24318 4140 24348 4740
rect 23276 3560 23308 3960
rect 23796 3560 23828 3960
rect 24316 3560 24348 3960
<< ndiff >>
rect 11158 14250 11238 14280
rect 11158 14210 11178 14250
rect 11218 14210 11238 14250
rect 11158 14150 11238 14210
rect 11158 14110 11178 14150
rect 11218 14110 11238 14150
rect 11158 14080 11238 14110
rect 13238 14250 13318 14280
rect 13238 14210 13258 14250
rect 13298 14210 13318 14250
rect 13238 14150 13318 14210
rect 13238 14110 13258 14150
rect 13298 14110 13318 14150
rect 13238 14080 13318 14110
rect 15318 14250 15398 14280
rect 15318 14210 15338 14250
rect 15378 14210 15398 14250
rect 15318 14150 15398 14210
rect 15318 14110 15338 14150
rect 15378 14110 15398 14150
rect 15318 14080 15398 14110
rect 10738 13640 10818 13670
rect 10738 13600 10758 13640
rect 10798 13600 10818 13640
rect 10738 13540 10818 13600
rect 10738 13500 10758 13540
rect 10798 13500 10818 13540
rect 10738 13440 10818 13500
rect 10738 13400 10758 13440
rect 10798 13400 10818 13440
rect 10738 13340 10818 13400
rect 10738 13300 10758 13340
rect 10798 13300 10818 13340
rect 10738 13240 10818 13300
rect 10738 13200 10758 13240
rect 10798 13200 10818 13240
rect 10738 13170 10818 13200
rect 11818 13640 11898 13670
rect 11978 13640 12058 13670
rect 11818 13600 11838 13640
rect 11878 13600 11898 13640
rect 11978 13600 11998 13640
rect 12038 13600 12058 13640
rect 11818 13540 11898 13600
rect 11978 13540 12058 13600
rect 11818 13500 11838 13540
rect 11878 13500 11898 13540
rect 11978 13500 11998 13540
rect 12038 13500 12058 13540
rect 11818 13440 11898 13500
rect 11978 13440 12058 13500
rect 11818 13400 11838 13440
rect 11878 13400 11898 13440
rect 11978 13400 11998 13440
rect 12038 13400 12058 13440
rect 11818 13340 11898 13400
rect 11978 13340 12058 13400
rect 11818 13300 11838 13340
rect 11878 13300 11898 13340
rect 11978 13300 11998 13340
rect 12038 13300 12058 13340
rect 11818 13240 11898 13300
rect 11978 13240 12058 13300
rect 11818 13200 11838 13240
rect 11878 13200 11898 13240
rect 11978 13200 11998 13240
rect 12038 13200 12058 13240
rect 11818 13170 11898 13200
rect 11978 13170 12058 13200
rect 13058 13640 13138 13670
rect 13058 13600 13078 13640
rect 13118 13600 13138 13640
rect 13058 13540 13138 13600
rect 13058 13500 13078 13540
rect 13118 13500 13138 13540
rect 13058 13440 13138 13500
rect 13058 13400 13078 13440
rect 13118 13400 13138 13440
rect 13058 13340 13138 13400
rect 13058 13300 13078 13340
rect 13118 13300 13138 13340
rect 13058 13240 13138 13300
rect 13058 13200 13078 13240
rect 13118 13200 13138 13240
rect 13058 13170 13138 13200
rect 13418 13640 13498 13670
rect 13418 13600 13438 13640
rect 13478 13600 13498 13640
rect 13418 13540 13498 13600
rect 13418 13500 13438 13540
rect 13478 13500 13498 13540
rect 13418 13440 13498 13500
rect 13418 13400 13438 13440
rect 13478 13400 13498 13440
rect 13418 13340 13498 13400
rect 13418 13300 13438 13340
rect 13478 13300 13498 13340
rect 13418 13240 13498 13300
rect 13418 13200 13438 13240
rect 13478 13200 13498 13240
rect 13418 13170 13498 13200
rect 14498 13660 14738 13670
rect 14498 13640 14578 13660
rect 14658 13640 14738 13660
rect 14498 13600 14518 13640
rect 14558 13600 14578 13640
rect 14658 13600 14678 13640
rect 14718 13600 14738 13640
rect 14498 13540 14578 13600
rect 14658 13540 14738 13600
rect 14498 13500 14518 13540
rect 14558 13500 14578 13540
rect 14658 13500 14678 13540
rect 14718 13500 14738 13540
rect 14498 13440 14578 13500
rect 14658 13440 14738 13500
rect 14498 13400 14518 13440
rect 14558 13400 14578 13440
rect 14658 13400 14678 13440
rect 14718 13400 14738 13440
rect 14498 13340 14578 13400
rect 14658 13340 14738 13400
rect 14498 13300 14518 13340
rect 14558 13300 14578 13340
rect 14658 13300 14678 13340
rect 14718 13300 14738 13340
rect 14498 13240 14578 13300
rect 14658 13240 14738 13300
rect 14498 13200 14518 13240
rect 14558 13200 14578 13240
rect 14658 13200 14678 13240
rect 14718 13200 14738 13240
rect 14498 13170 14578 13200
rect 14658 13170 14738 13200
rect 15738 13640 15818 13670
rect 15738 13600 15758 13640
rect 15798 13600 15818 13640
rect 15738 13540 15818 13600
rect 15738 13500 15758 13540
rect 15798 13500 15818 13540
rect 15738 13440 15818 13500
rect 15738 13400 15758 13440
rect 15798 13400 15818 13440
rect 15738 13340 15818 13400
rect 15738 13300 15758 13340
rect 15798 13300 15818 13340
rect 15738 13240 15818 13300
rect 15738 13200 15758 13240
rect 15798 13200 15818 13240
rect 15738 13170 15818 13200
rect 11358 12630 11438 12660
rect 11358 12590 11378 12630
rect 11418 12590 11438 12630
rect 11358 12560 11438 12590
rect 11478 12630 11558 12660
rect 11478 12590 11498 12630
rect 11538 12590 11558 12630
rect 11478 12560 11558 12590
rect 11598 12630 11678 12660
rect 11598 12590 11618 12630
rect 11658 12590 11678 12630
rect 11598 12560 11678 12590
rect 11718 12630 11798 12660
rect 11718 12590 11738 12630
rect 11778 12590 11798 12630
rect 11718 12560 11798 12590
rect 11838 12630 11918 12660
rect 11838 12590 11858 12630
rect 11898 12590 11918 12630
rect 11838 12560 11918 12590
rect 11958 12630 12038 12660
rect 11958 12590 11978 12630
rect 12018 12590 12038 12630
rect 11958 12560 12038 12590
rect 12078 12630 12158 12660
rect 12078 12590 12098 12630
rect 12138 12590 12158 12630
rect 12078 12560 12158 12590
rect 12198 12630 12278 12660
rect 12198 12590 12218 12630
rect 12258 12590 12278 12630
rect 12198 12560 12278 12590
rect 12318 12630 12398 12660
rect 12318 12590 12338 12630
rect 12378 12590 12398 12630
rect 12318 12560 12398 12590
rect 12438 12630 12518 12660
rect 12438 12590 12458 12630
rect 12498 12590 12518 12630
rect 12438 12560 12518 12590
rect 12558 12630 12638 12660
rect 12558 12590 12578 12630
rect 12618 12590 12638 12630
rect 12558 12560 12638 12590
rect 13918 12630 13998 12660
rect 13918 12590 13938 12630
rect 13978 12590 13998 12630
rect 13918 12560 13998 12590
rect 14038 12630 14118 12660
rect 14038 12590 14058 12630
rect 14098 12590 14118 12630
rect 14038 12560 14118 12590
rect 14158 12630 14238 12660
rect 14158 12590 14178 12630
rect 14218 12590 14238 12630
rect 14158 12560 14238 12590
rect 14278 12630 14358 12660
rect 14278 12590 14298 12630
rect 14338 12590 14358 12630
rect 14278 12560 14358 12590
rect 14398 12630 14478 12660
rect 14398 12590 14418 12630
rect 14458 12590 14478 12630
rect 14398 12560 14478 12590
rect 14518 12630 14598 12660
rect 14518 12590 14538 12630
rect 14578 12590 14598 12630
rect 14518 12560 14598 12590
rect 14638 12630 14718 12660
rect 14638 12590 14658 12630
rect 14698 12590 14718 12630
rect 14638 12560 14718 12590
rect 14758 12630 14838 12660
rect 14758 12590 14778 12630
rect 14818 12590 14838 12630
rect 14758 12560 14838 12590
rect 14878 12630 14958 12660
rect 14878 12590 14898 12630
rect 14938 12590 14958 12630
rect 14878 12560 14958 12590
rect 14998 12630 15078 12660
rect 14998 12590 15018 12630
rect 15058 12590 15078 12630
rect 14998 12560 15078 12590
rect 15118 12630 15198 12660
rect 15118 12590 15138 12630
rect 15178 12590 15198 12630
rect 15118 12560 15198 12590
rect 19438 11030 19538 11060
rect 19438 10990 19468 11030
rect 19508 10990 19538 11030
rect 19438 10960 19538 10990
rect 19568 11030 19668 11060
rect 19568 10990 19598 11030
rect 19638 10990 19668 11030
rect 19568 10960 19668 10990
rect 19698 11030 19798 11060
rect 19698 10990 19728 11030
rect 19768 10990 19798 11030
rect 19698 10960 19798 10990
rect 19828 11030 19928 11060
rect 19828 10990 19858 11030
rect 19898 10990 19928 11030
rect 19828 10960 19928 10990
rect 19958 11030 20058 11060
rect 19958 10990 19988 11030
rect 20028 10990 20058 11030
rect 19958 10960 20058 10990
rect 20088 11030 20188 11060
rect 20088 10990 20118 11030
rect 20158 10990 20188 11030
rect 20088 10960 20188 10990
rect 20218 11030 20318 11060
rect 20218 10990 20248 11030
rect 20288 10990 20318 11030
rect 20218 10960 20318 10990
rect 20578 11030 20678 11060
rect 20578 10990 20608 11030
rect 20648 10990 20678 11030
rect 20578 10960 20678 10990
rect 20708 11030 20808 11060
rect 20708 10990 20738 11030
rect 20778 10990 20808 11030
rect 20708 10960 20808 10990
rect 20838 11030 20938 11060
rect 20838 10990 20868 11030
rect 20908 10990 20938 11030
rect 20838 10960 20938 10990
rect 20968 11030 21068 11060
rect 20968 10990 20998 11030
rect 21038 10990 21068 11030
rect 20968 10960 21068 10990
rect 21098 11030 21198 11060
rect 21098 10990 21128 11030
rect 21168 10990 21198 11030
rect 21098 10960 21198 10990
rect 21228 11030 21328 11060
rect 21228 10990 21258 11030
rect 21298 10990 21328 11030
rect 21228 10960 21328 10990
rect 21358 11030 21458 11060
rect 21358 10990 21388 11030
rect 21428 10990 21458 11030
rect 21358 10960 21458 10990
rect 21718 11030 21818 11060
rect 21718 10990 21748 11030
rect 21788 10990 21818 11030
rect 21718 10960 21818 10990
rect 21848 11030 21948 11060
rect 21848 10990 21878 11030
rect 21918 10990 21948 11030
rect 21848 10960 21948 10990
rect 21978 11030 22078 11060
rect 21978 10990 22008 11030
rect 22048 10990 22078 11030
rect 21978 10960 22078 10990
rect 22108 11030 22208 11060
rect 22108 10990 22138 11030
rect 22178 10990 22208 11030
rect 22108 10960 22208 10990
rect 22238 11030 22338 11060
rect 22238 10990 22268 11030
rect 22308 10990 22338 11030
rect 22238 10960 22338 10990
rect 22368 11030 22468 11060
rect 22368 10990 22398 11030
rect 22438 10990 22468 11030
rect 22368 10960 22468 10990
rect 22498 11030 22598 11060
rect 22498 10990 22528 11030
rect 22568 10990 22598 11030
rect 22498 10960 22598 10990
rect 19388 10490 19488 10520
rect 19388 10440 19418 10490
rect 19458 10440 19488 10490
rect 19388 10350 19488 10440
rect 19388 10300 19418 10350
rect 19458 10300 19488 10350
rect 19388 10270 19488 10300
rect 19588 10490 19688 10520
rect 19588 10440 19618 10490
rect 19658 10440 19688 10490
rect 19588 10350 19688 10440
rect 19588 10300 19618 10350
rect 19658 10300 19688 10350
rect 19588 10270 19688 10300
rect 19788 10490 19888 10520
rect 19788 10440 19818 10490
rect 19858 10440 19888 10490
rect 19788 10350 19888 10440
rect 19788 10300 19818 10350
rect 19858 10300 19888 10350
rect 19788 10270 19888 10300
rect 19988 10490 20088 10520
rect 19988 10440 20018 10490
rect 20058 10440 20088 10490
rect 19988 10350 20088 10440
rect 19988 10300 20018 10350
rect 20058 10300 20088 10350
rect 19988 10270 20088 10300
rect 20188 10490 20288 10520
rect 20188 10440 20218 10490
rect 20258 10440 20288 10490
rect 20188 10350 20288 10440
rect 20188 10300 20218 10350
rect 20258 10300 20288 10350
rect 20188 10270 20288 10300
rect 20388 10490 20488 10520
rect 20388 10440 20418 10490
rect 20458 10440 20488 10490
rect 20388 10350 20488 10440
rect 20388 10300 20418 10350
rect 20458 10300 20488 10350
rect 20388 10270 20488 10300
rect 20588 10490 20688 10520
rect 20588 10440 20618 10490
rect 20658 10440 20688 10490
rect 20588 10350 20688 10440
rect 20588 10300 20618 10350
rect 20658 10300 20688 10350
rect 20588 10270 20688 10300
rect 20788 10490 20888 10520
rect 20788 10440 20818 10490
rect 20858 10440 20888 10490
rect 20788 10350 20888 10440
rect 20788 10300 20818 10350
rect 20858 10300 20888 10350
rect 20788 10270 20888 10300
rect 20988 10490 21088 10520
rect 20988 10440 21018 10490
rect 21058 10440 21088 10490
rect 20988 10350 21088 10440
rect 20988 10300 21018 10350
rect 21058 10300 21088 10350
rect 20988 10270 21088 10300
rect 21188 10490 21288 10520
rect 21188 10440 21218 10490
rect 21258 10440 21288 10490
rect 21188 10350 21288 10440
rect 21188 10300 21218 10350
rect 21258 10300 21288 10350
rect 21188 10270 21288 10300
rect 21388 10490 21488 10520
rect 21388 10440 21418 10490
rect 21458 10440 21488 10490
rect 21388 10350 21488 10440
rect 21388 10300 21418 10350
rect 21458 10300 21488 10350
rect 21388 10270 21488 10300
rect 13248 8060 13328 8090
rect 13248 8020 13268 8060
rect 13308 8020 13328 8060
rect 13248 7960 13328 8020
rect 13248 7920 13268 7960
rect 13308 7920 13328 7960
rect 13248 7890 13328 7920
rect 13358 8060 13438 8090
rect 13358 8020 13378 8060
rect 13418 8020 13438 8060
rect 13358 7960 13438 8020
rect 13358 7920 13378 7960
rect 13418 7920 13438 7960
rect 13358 7890 13438 7920
rect 13468 8060 13548 8090
rect 13468 8020 13488 8060
rect 13528 8020 13548 8060
rect 13468 7960 13548 8020
rect 13468 7920 13488 7960
rect 13528 7920 13548 7960
rect 13468 7890 13548 7920
rect 13768 8060 13848 8090
rect 13768 8020 13788 8060
rect 13828 8020 13848 8060
rect 13768 7960 13848 8020
rect 13768 7920 13788 7960
rect 13828 7920 13848 7960
rect 13768 7890 13848 7920
rect 13878 8060 13958 8090
rect 13878 8020 13898 8060
rect 13938 8020 13958 8060
rect 13878 7960 13958 8020
rect 13878 7920 13898 7960
rect 13938 7920 13958 7960
rect 13878 7890 13958 7920
rect 13988 8060 14068 8090
rect 14148 8060 14228 8090
rect 13988 8020 14008 8060
rect 14048 8020 14068 8060
rect 14148 8020 14168 8060
rect 14208 8020 14228 8060
rect 13988 7960 14068 8020
rect 14148 7960 14228 8020
rect 13988 7920 14008 7960
rect 14048 7920 14068 7960
rect 14148 7920 14168 7960
rect 14208 7920 14228 7960
rect 13988 7890 14068 7920
rect 14148 7890 14228 7920
rect 14258 8060 14338 8090
rect 14258 8020 14278 8060
rect 14318 8020 14338 8060
rect 14258 7960 14338 8020
rect 14258 7920 14278 7960
rect 14318 7920 14338 7960
rect 14258 7890 14338 7920
rect 14368 8060 14448 8090
rect 14368 8020 14388 8060
rect 14428 8020 14448 8060
rect 14368 7960 14448 8020
rect 14368 7920 14388 7960
rect 14428 7920 14448 7960
rect 14368 7890 14448 7920
rect 14668 8060 14748 8090
rect 14668 8020 14688 8060
rect 14728 8020 14748 8060
rect 14668 7960 14748 8020
rect 14668 7920 14688 7960
rect 14728 7920 14748 7960
rect 14668 7890 14748 7920
rect 14778 8060 14858 8090
rect 14778 8020 14798 8060
rect 14838 8020 14858 8060
rect 14778 7960 14858 8020
rect 14778 7920 14798 7960
rect 14838 7920 14858 7960
rect 14778 7890 14858 7920
rect 14888 8060 14968 8090
rect 14888 8020 14908 8060
rect 14948 8020 14968 8060
rect 14888 7960 14968 8020
rect 14888 7920 14908 7960
rect 14948 7920 14968 7960
rect 14888 7890 14968 7920
rect 15178 8060 15258 8090
rect 15178 8020 15198 8060
rect 15238 8020 15258 8060
rect 15178 7960 15258 8020
rect 15178 7920 15198 7960
rect 15238 7920 15258 7960
rect 15178 7890 15258 7920
rect 15288 8060 15368 8090
rect 15288 8020 15308 8060
rect 15348 8020 15368 8060
rect 15288 7960 15368 8020
rect 15288 7920 15308 7960
rect 15348 7920 15368 7960
rect 15288 7890 15368 7920
rect 15508 8060 15588 8090
rect 15508 8020 15528 8060
rect 15568 8020 15588 8060
rect 15508 7960 15588 8020
rect 15508 7920 15528 7960
rect 15568 7920 15588 7960
rect 15508 7890 15588 7920
rect 15618 8060 15698 8090
rect 15618 8020 15638 8060
rect 15678 8020 15698 8060
rect 15618 7960 15698 8020
rect 15618 7920 15638 7960
rect 15678 7920 15698 7960
rect 15618 7890 15698 7920
rect 15838 8060 15918 8090
rect 15838 8020 15858 8060
rect 15898 8020 15918 8060
rect 15838 7960 15918 8020
rect 15838 7920 15858 7960
rect 15898 7920 15918 7960
rect 15838 7890 15918 7920
rect 15948 8060 16028 8090
rect 15948 8020 15968 8060
rect 16008 8020 16028 8060
rect 15948 7960 16028 8020
rect 15948 7920 15968 7960
rect 16008 7920 16028 7960
rect 15948 7890 16028 7920
rect 16378 8060 16478 8090
rect 16378 8020 16408 8060
rect 16448 8020 16478 8060
rect 16378 7960 16478 8020
rect 16378 7920 16408 7960
rect 16448 7920 16478 7960
rect 16378 7890 16478 7920
rect 16508 8060 16608 8090
rect 16508 8020 16538 8060
rect 16578 8020 16608 8060
rect 16508 7960 16608 8020
rect 16508 7920 16538 7960
rect 16578 7920 16608 7960
rect 16508 7890 16608 7920
rect 16768 8060 16868 8090
rect 16768 8020 16798 8060
rect 16838 8020 16868 8060
rect 16768 7960 16868 8020
rect 16768 7920 16798 7960
rect 16838 7920 16868 7960
rect 16768 7890 16868 7920
rect 16898 8060 16998 8090
rect 16898 8020 16928 8060
rect 16968 8020 16998 8060
rect 16898 7960 16998 8020
rect 16898 7920 16928 7960
rect 16968 7920 16998 7960
rect 16898 7890 16998 7920
rect 17158 8060 17258 8090
rect 17158 8020 17188 8060
rect 17228 8020 17258 8060
rect 17158 7960 17258 8020
rect 17158 7920 17188 7960
rect 17228 7920 17258 7960
rect 17158 7890 17258 7920
rect 17288 8060 17388 8090
rect 17288 8020 17318 8060
rect 17358 8020 17388 8060
rect 17288 7960 17388 8020
rect 17288 7920 17318 7960
rect 17358 7920 17388 7960
rect 17288 7890 17388 7920
rect 17448 8060 17548 8090
rect 17448 8020 17478 8060
rect 17518 8020 17548 8060
rect 17448 7960 17548 8020
rect 17448 7920 17478 7960
rect 17518 7920 17548 7960
rect 17448 7890 17548 7920
rect 17578 8060 17678 8090
rect 17578 8020 17608 8060
rect 17648 8020 17678 8060
rect 17578 7960 17678 8020
rect 17578 7920 17608 7960
rect 17648 7920 17678 7960
rect 17578 7890 17678 7920
rect 17838 8060 17938 8090
rect 17838 8020 17868 8060
rect 17908 8020 17938 8060
rect 17838 7960 17938 8020
rect 17838 7920 17868 7960
rect 17908 7920 17938 7960
rect 17838 7890 17938 7920
rect 17968 8060 18068 8090
rect 17968 8020 17998 8060
rect 18038 8020 18068 8060
rect 17968 7960 18068 8020
rect 17968 7920 17998 7960
rect 18038 7920 18068 7960
rect 17968 7890 18068 7920
rect 19328 8010 19428 8040
rect 19328 7970 19358 8010
rect 19398 7970 19428 8010
rect 19328 7910 19428 7970
rect 19328 7870 19358 7910
rect 19398 7870 19428 7910
rect 19328 7810 19428 7870
rect 19328 7770 19358 7810
rect 19398 7770 19428 7810
rect 19328 7710 19428 7770
rect 19328 7670 19358 7710
rect 19398 7670 19428 7710
rect 19328 7640 19428 7670
rect 19548 8010 19648 8040
rect 19548 7970 19578 8010
rect 19618 7970 19648 8010
rect 19548 7910 19648 7970
rect 19548 7870 19578 7910
rect 19618 7870 19648 7910
rect 19548 7810 19648 7870
rect 19548 7770 19578 7810
rect 19618 7770 19648 7810
rect 19548 7710 19648 7770
rect 19548 7670 19578 7710
rect 19618 7670 19648 7710
rect 19548 7640 19648 7670
rect 19768 8010 19868 8040
rect 19768 7970 19798 8010
rect 19838 7970 19868 8010
rect 19768 7910 19868 7970
rect 19768 7870 19798 7910
rect 19838 7870 19868 7910
rect 19768 7810 19868 7870
rect 19768 7770 19798 7810
rect 19838 7770 19868 7810
rect 19768 7710 19868 7770
rect 19768 7670 19798 7710
rect 19838 7670 19868 7710
rect 19768 7640 19868 7670
rect 19988 8010 20088 8040
rect 19988 7970 20018 8010
rect 20058 7970 20088 8010
rect 19988 7910 20088 7970
rect 19988 7870 20018 7910
rect 20058 7870 20088 7910
rect 19988 7810 20088 7870
rect 19988 7770 20018 7810
rect 20058 7770 20088 7810
rect 19988 7710 20088 7770
rect 19988 7670 20018 7710
rect 20058 7670 20088 7710
rect 19988 7640 20088 7670
rect 20208 8010 20308 8040
rect 20408 8010 20508 8040
rect 20208 7970 20238 8010
rect 20278 7970 20308 8010
rect 20408 7970 20438 8010
rect 20478 7970 20508 8010
rect 20208 7910 20308 7970
rect 20408 7910 20508 7970
rect 20208 7870 20238 7910
rect 20278 7870 20308 7910
rect 20408 7870 20438 7910
rect 20478 7870 20508 7910
rect 20208 7810 20308 7870
rect 20408 7810 20508 7870
rect 20208 7770 20238 7810
rect 20278 7770 20308 7810
rect 20408 7770 20438 7810
rect 20478 7770 20508 7810
rect 20208 7710 20308 7770
rect 20408 7710 20508 7770
rect 20208 7670 20238 7710
rect 20278 7670 20308 7710
rect 20408 7670 20438 7710
rect 20478 7670 20508 7710
rect 20208 7640 20308 7670
rect 20408 7640 20508 7670
rect 20628 8010 20728 8040
rect 20628 7970 20658 8010
rect 20698 7970 20728 8010
rect 20628 7910 20728 7970
rect 20628 7870 20658 7910
rect 20698 7870 20728 7910
rect 20628 7810 20728 7870
rect 20628 7770 20658 7810
rect 20698 7770 20728 7810
rect 20628 7710 20728 7770
rect 20628 7670 20658 7710
rect 20698 7670 20728 7710
rect 20628 7640 20728 7670
rect 20848 8010 20948 8040
rect 20848 7970 20878 8010
rect 20918 7970 20948 8010
rect 20848 7910 20948 7970
rect 20848 7870 20878 7910
rect 20918 7870 20948 7910
rect 20848 7810 20948 7870
rect 20848 7770 20878 7810
rect 20918 7770 20948 7810
rect 20848 7710 20948 7770
rect 20848 7670 20878 7710
rect 20918 7670 20948 7710
rect 20848 7640 20948 7670
rect 21068 8010 21168 8040
rect 21068 7970 21098 8010
rect 21138 7970 21168 8010
rect 21068 7910 21168 7970
rect 21068 7870 21098 7910
rect 21138 7870 21168 7910
rect 21068 7810 21168 7870
rect 21068 7770 21098 7810
rect 21138 7770 21168 7810
rect 21068 7710 21168 7770
rect 21068 7670 21098 7710
rect 21138 7670 21168 7710
rect 21068 7640 21168 7670
rect 21288 8010 21388 8040
rect 21488 8010 21588 8040
rect 21288 7970 21318 8010
rect 21358 7970 21388 8010
rect 21488 7970 21518 8010
rect 21558 7970 21588 8010
rect 21288 7910 21388 7970
rect 21488 7910 21588 7970
rect 21288 7870 21318 7910
rect 21358 7870 21388 7910
rect 21488 7870 21518 7910
rect 21558 7870 21588 7910
rect 21288 7810 21388 7870
rect 21488 7810 21588 7870
rect 21288 7770 21318 7810
rect 21358 7770 21388 7810
rect 21488 7770 21518 7810
rect 21558 7770 21588 7810
rect 21288 7710 21388 7770
rect 21488 7710 21588 7770
rect 21288 7670 21318 7710
rect 21358 7670 21388 7710
rect 21488 7670 21518 7710
rect 21558 7670 21588 7710
rect 21288 7640 21388 7670
rect 21488 7640 21588 7670
rect 21708 8010 21808 8040
rect 21708 7970 21738 8010
rect 21778 7970 21808 8010
rect 21708 7910 21808 7970
rect 21708 7870 21738 7910
rect 21778 7870 21808 7910
rect 21708 7810 21808 7870
rect 21708 7770 21738 7810
rect 21778 7770 21808 7810
rect 21708 7710 21808 7770
rect 21708 7670 21738 7710
rect 21778 7670 21808 7710
rect 21708 7640 21808 7670
rect 21928 8010 22028 8040
rect 21928 7970 21958 8010
rect 21998 7970 22028 8010
rect 21928 7910 22028 7970
rect 21928 7870 21958 7910
rect 21998 7870 22028 7910
rect 21928 7810 22028 7870
rect 21928 7770 21958 7810
rect 21998 7770 22028 7810
rect 21928 7710 22028 7770
rect 21928 7670 21958 7710
rect 21998 7670 22028 7710
rect 21928 7640 22028 7670
rect 22148 8010 22248 8040
rect 22148 7970 22178 8010
rect 22218 7970 22248 8010
rect 22148 7910 22248 7970
rect 22148 7870 22178 7910
rect 22218 7870 22248 7910
rect 22148 7810 22248 7870
rect 22148 7770 22178 7810
rect 22218 7770 22248 7810
rect 22148 7710 22248 7770
rect 22148 7670 22178 7710
rect 22218 7670 22248 7710
rect 22148 7640 22248 7670
rect 22368 8010 22468 8040
rect 22368 7970 22398 8010
rect 22438 7970 22468 8010
rect 22368 7910 22468 7970
rect 22368 7870 22398 7910
rect 22438 7870 22468 7910
rect 22368 7810 22468 7870
rect 22368 7770 22398 7810
rect 22438 7770 22468 7810
rect 22368 7710 22468 7770
rect 22368 7670 22398 7710
rect 22438 7670 22468 7710
rect 22368 7640 22468 7670
rect 13248 6260 13328 6290
rect 13248 6220 13268 6260
rect 13308 6220 13328 6260
rect 13248 6160 13328 6220
rect 13248 6120 13268 6160
rect 13308 6120 13328 6160
rect 13248 6090 13328 6120
rect 13358 6260 13438 6290
rect 13358 6220 13378 6260
rect 13418 6220 13438 6260
rect 13358 6160 13438 6220
rect 13358 6120 13378 6160
rect 13418 6120 13438 6160
rect 13358 6090 13438 6120
rect 13468 6260 13548 6290
rect 13468 6220 13488 6260
rect 13528 6220 13548 6260
rect 13468 6160 13548 6220
rect 13468 6120 13488 6160
rect 13528 6120 13548 6160
rect 13468 6090 13548 6120
rect 13768 6260 13848 6290
rect 13768 6220 13788 6260
rect 13828 6220 13848 6260
rect 13768 6160 13848 6220
rect 13768 6120 13788 6160
rect 13828 6120 13848 6160
rect 13768 6090 13848 6120
rect 13878 6260 13958 6290
rect 13878 6220 13898 6260
rect 13938 6220 13958 6260
rect 13878 6160 13958 6220
rect 13878 6120 13898 6160
rect 13938 6120 13958 6160
rect 13878 6090 13958 6120
rect 13988 6260 14068 6290
rect 14148 6260 14228 6290
rect 13988 6220 14008 6260
rect 14048 6220 14068 6260
rect 14148 6220 14168 6260
rect 14208 6220 14228 6260
rect 13988 6160 14068 6220
rect 14148 6160 14228 6220
rect 13988 6120 14008 6160
rect 14048 6120 14068 6160
rect 14148 6120 14168 6160
rect 14208 6120 14228 6160
rect 13988 6090 14068 6120
rect 14148 6090 14228 6120
rect 14258 6260 14338 6290
rect 14258 6220 14278 6260
rect 14318 6220 14338 6260
rect 14258 6160 14338 6220
rect 14258 6120 14278 6160
rect 14318 6120 14338 6160
rect 14258 6090 14338 6120
rect 14368 6260 14448 6290
rect 14368 6220 14388 6260
rect 14428 6220 14448 6260
rect 14368 6160 14448 6220
rect 14368 6120 14388 6160
rect 14428 6120 14448 6160
rect 14368 6090 14448 6120
rect 14668 6260 14748 6290
rect 14668 6220 14688 6260
rect 14728 6220 14748 6260
rect 14668 6160 14748 6220
rect 14668 6120 14688 6160
rect 14728 6120 14748 6160
rect 14668 6090 14748 6120
rect 14778 6260 14858 6290
rect 14778 6220 14798 6260
rect 14838 6220 14858 6260
rect 14778 6160 14858 6220
rect 14778 6120 14798 6160
rect 14838 6120 14858 6160
rect 14778 6090 14858 6120
rect 14888 6260 14968 6290
rect 14888 6220 14908 6260
rect 14948 6220 14968 6260
rect 14888 6160 14968 6220
rect 14888 6120 14908 6160
rect 14948 6120 14968 6160
rect 14888 6090 14968 6120
rect 15188 6260 15268 6290
rect 15188 6220 15208 6260
rect 15248 6220 15268 6260
rect 15188 6160 15268 6220
rect 15188 6120 15208 6160
rect 15248 6120 15268 6160
rect 15188 6090 15268 6120
rect 15298 6260 15378 6290
rect 15298 6220 15318 6260
rect 15358 6220 15378 6260
rect 15298 6160 15378 6220
rect 15298 6120 15318 6160
rect 15358 6120 15378 6160
rect 15298 6090 15378 6120
rect 15408 6260 15488 6290
rect 15408 6220 15428 6260
rect 15468 6220 15488 6260
rect 15408 6160 15488 6220
rect 15408 6120 15428 6160
rect 15468 6120 15488 6160
rect 15408 6090 15488 6120
rect 15628 6260 15708 6290
rect 15628 6220 15648 6260
rect 15688 6220 15708 6260
rect 15628 6160 15708 6220
rect 15628 6120 15648 6160
rect 15688 6120 15708 6160
rect 15628 6090 15708 6120
rect 15738 6260 15818 6290
rect 15738 6220 15758 6260
rect 15798 6220 15818 6260
rect 15738 6160 15818 6220
rect 15738 6120 15758 6160
rect 15798 6120 15818 6160
rect 15738 6090 15818 6120
rect 15958 6260 16038 6290
rect 15958 6220 15978 6260
rect 16018 6220 16038 6260
rect 15958 6160 16038 6220
rect 15958 6120 15978 6160
rect 16018 6120 16038 6160
rect 15958 6090 16038 6120
rect 16068 6260 16148 6290
rect 16068 6220 16088 6260
rect 16128 6220 16148 6260
rect 16068 6160 16148 6220
rect 16068 6120 16088 6160
rect 16128 6120 16148 6160
rect 16068 6090 16148 6120
rect 16378 6260 16478 6290
rect 16378 6220 16408 6260
rect 16448 6220 16478 6260
rect 16378 6160 16478 6220
rect 16378 6120 16408 6160
rect 16448 6120 16478 6160
rect 16378 6090 16478 6120
rect 16508 6260 16608 6290
rect 16508 6220 16538 6260
rect 16578 6220 16608 6260
rect 16508 6160 16608 6220
rect 16508 6120 16538 6160
rect 16578 6120 16608 6160
rect 16508 6090 16608 6120
rect 16768 6260 16868 6290
rect 16768 6220 16798 6260
rect 16838 6220 16868 6260
rect 16768 6160 16868 6220
rect 16768 6120 16798 6160
rect 16838 6120 16868 6160
rect 16768 6090 16868 6120
rect 16898 6260 16998 6290
rect 16898 6220 16928 6260
rect 16968 6220 16998 6260
rect 16898 6160 16998 6220
rect 16898 6120 16928 6160
rect 16968 6120 16998 6160
rect 16898 6090 16998 6120
rect 17158 6260 17258 6290
rect 17158 6220 17188 6260
rect 17228 6220 17258 6260
rect 17158 6160 17258 6220
rect 17158 6120 17188 6160
rect 17228 6120 17258 6160
rect 17158 6090 17258 6120
rect 17288 6260 17388 6290
rect 17288 6220 17318 6260
rect 17358 6220 17388 6260
rect 17288 6160 17388 6220
rect 17288 6120 17318 6160
rect 17358 6120 17388 6160
rect 17288 6090 17388 6120
rect 17448 6260 17548 6290
rect 17448 6220 17478 6260
rect 17518 6220 17548 6260
rect 17448 6160 17548 6220
rect 17448 6120 17478 6160
rect 17518 6120 17548 6160
rect 17448 6090 17548 6120
rect 17578 6260 17678 6290
rect 17578 6220 17608 6260
rect 17648 6220 17678 6260
rect 17578 6160 17678 6220
rect 17578 6120 17608 6160
rect 17648 6120 17678 6160
rect 17578 6090 17678 6120
rect 12428 3180 12508 3210
rect 12428 3140 12448 3180
rect 12488 3140 12508 3180
rect 12428 3110 12508 3140
rect 12538 3180 12618 3210
rect 12538 3140 12558 3180
rect 12598 3140 12618 3180
rect 12538 3110 12618 3140
rect 12648 3180 12728 3210
rect 12648 3140 12668 3180
rect 12708 3140 12728 3180
rect 12648 3110 12728 3140
rect 12758 3180 12838 3210
rect 12758 3140 12778 3180
rect 12818 3140 12838 3180
rect 12758 3110 12838 3140
rect 12868 3180 12948 3210
rect 12868 3140 12888 3180
rect 12928 3140 12948 3180
rect 12868 3110 12948 3140
rect 13008 3180 13088 3210
rect 13008 3140 13028 3180
rect 13068 3140 13088 3180
rect 13008 3110 13088 3140
rect 13118 3180 13198 3210
rect 13118 3140 13138 3180
rect 13178 3140 13198 3180
rect 13118 3110 13198 3140
rect 13228 3180 13308 3210
rect 13228 3140 13248 3180
rect 13288 3140 13308 3180
rect 13228 3110 13308 3140
rect 13458 3180 13538 3210
rect 13458 3140 13478 3180
rect 13518 3140 13538 3180
rect 13458 3110 13538 3140
rect 13568 3180 13648 3210
rect 13568 3140 13588 3180
rect 13628 3140 13648 3180
rect 13568 3110 13648 3140
rect 13678 3180 13758 3210
rect 13678 3140 13698 3180
rect 13738 3140 13758 3180
rect 13678 3110 13758 3140
rect 13788 3180 13868 3210
rect 13788 3140 13808 3180
rect 13848 3140 13868 3180
rect 13788 3110 13868 3140
rect 13898 3180 13978 3210
rect 13898 3140 13918 3180
rect 13958 3140 13978 3180
rect 13898 3110 13978 3140
rect 14118 3180 14198 3210
rect 14118 3140 14138 3180
rect 14178 3140 14198 3180
rect 14118 3110 14198 3140
rect 14228 3180 14308 3210
rect 14228 3140 14248 3180
rect 14288 3140 14308 3180
rect 14228 3110 14308 3140
rect 14338 3180 14418 3210
rect 14338 3140 14358 3180
rect 14398 3140 14418 3180
rect 14338 3110 14418 3140
rect 14448 3180 14528 3210
rect 14448 3140 14468 3180
rect 14508 3140 14528 3180
rect 14448 3110 14528 3140
rect 14558 3180 14638 3210
rect 14558 3140 14578 3180
rect 14618 3140 14638 3180
rect 14558 3110 14638 3140
rect 14798 3180 14878 3210
rect 14798 3140 14818 3180
rect 14858 3140 14878 3180
rect 14798 3110 14878 3140
rect 14908 3180 14988 3210
rect 14908 3140 14928 3180
rect 14968 3140 14988 3180
rect 14908 3110 14988 3140
rect 15018 3180 15098 3210
rect 15018 3140 15038 3180
rect 15078 3140 15098 3180
rect 15018 3110 15098 3140
rect 15128 3180 15208 3210
rect 15128 3140 15148 3180
rect 15188 3140 15208 3180
rect 15128 3110 15208 3140
rect 15238 3180 15318 3210
rect 15238 3140 15258 3180
rect 15298 3140 15318 3180
rect 15238 3110 15318 3140
rect 15378 3180 15458 3210
rect 15378 3140 15398 3180
rect 15438 3140 15458 3180
rect 15378 3110 15458 3140
rect 15488 3180 15568 3210
rect 15488 3140 15508 3180
rect 15548 3140 15568 3180
rect 15488 3110 15568 3140
rect 15598 3180 15678 3210
rect 15598 3140 15618 3180
rect 15658 3140 15678 3180
rect 15598 3110 15678 3140
rect 15938 3180 16018 3210
rect 15938 3140 15958 3180
rect 15998 3140 16018 3180
rect 15938 3110 16018 3140
rect 16048 3180 16128 3210
rect 16048 3140 16068 3180
rect 16108 3140 16128 3180
rect 16048 3110 16128 3140
rect 16298 3180 16378 3210
rect 16298 3140 16318 3180
rect 16358 3140 16378 3180
rect 16298 3110 16378 3140
rect 16408 3180 16488 3210
rect 16408 3140 16428 3180
rect 16468 3140 16488 3180
rect 16408 3110 16488 3140
rect 16548 3180 16628 3210
rect 16548 3140 16568 3180
rect 16608 3140 16628 3180
rect 16548 3110 16628 3140
rect 16658 3180 16738 3210
rect 16658 3140 16678 3180
rect 16718 3140 16738 3180
rect 16658 3110 16738 3140
rect 16768 3180 16848 3210
rect 16768 3140 16788 3180
rect 16828 3140 16848 3180
rect 16768 3110 16848 3140
rect 16878 3180 16958 3210
rect 16878 3140 16898 3180
rect 16938 3140 16958 3180
rect 16878 3110 16958 3140
rect 16988 3180 17068 3210
rect 16988 3140 17008 3180
rect 17048 3140 17068 3180
rect 16988 3110 17068 3140
rect 17208 3180 17288 3210
rect 17208 3140 17228 3180
rect 17268 3140 17288 3180
rect 17208 3110 17288 3140
rect 17318 3180 17398 3210
rect 17318 3140 17338 3180
rect 17378 3140 17398 3180
rect 17318 3110 17398 3140
rect 17428 3180 17508 3210
rect 17428 3140 17448 3180
rect 17488 3140 17508 3180
rect 17428 3110 17508 3140
rect 17538 3180 17618 3210
rect 17538 3140 17558 3180
rect 17598 3140 17618 3180
rect 17538 3110 17618 3140
rect 17758 3180 17838 3210
rect 17758 3140 17778 3180
rect 17818 3140 17838 3180
rect 17758 3110 17838 3140
rect 17868 3180 17948 3210
rect 17868 3140 17888 3180
rect 17928 3140 17948 3180
rect 17868 3110 17948 3140
rect 17978 3180 18058 3210
rect 17978 3140 17998 3180
rect 18038 3140 18058 3180
rect 17978 3110 18058 3140
rect 18088 3180 18168 3210
rect 18088 3140 18108 3180
rect 18148 3140 18168 3180
rect 18088 3110 18168 3140
rect 18198 3180 18278 3210
rect 18198 3140 18218 3180
rect 18258 3140 18278 3180
rect 18198 3110 18278 3140
rect 18418 3180 18498 3210
rect 18418 3140 18438 3180
rect 18478 3140 18498 3180
rect 18418 3110 18498 3140
rect 18528 3180 18608 3210
rect 18528 3140 18548 3180
rect 18588 3140 18608 3180
rect 18528 3110 18608 3140
rect 18638 3180 18718 3210
rect 18638 3140 18658 3180
rect 18698 3140 18718 3180
rect 18638 3110 18718 3140
rect 18748 3180 18828 3210
rect 18748 3140 18768 3180
rect 18808 3140 18828 3180
rect 18748 3110 18828 3140
rect 19058 3090 19138 3120
rect 19058 3050 19078 3090
rect 19118 3050 19138 3090
rect 19058 3020 19138 3050
rect 19168 3090 19248 3120
rect 19168 3050 19188 3090
rect 19228 3050 19248 3090
rect 19168 3020 19248 3050
rect 19278 3090 19358 3120
rect 19278 3050 19298 3090
rect 19338 3050 19358 3090
rect 19278 3020 19358 3050
rect 19388 3090 19468 3120
rect 19388 3050 19408 3090
rect 19448 3050 19468 3090
rect 19388 3020 19468 3050
rect 19498 3090 19578 3120
rect 19498 3050 19518 3090
rect 19558 3050 19578 3090
rect 19498 3020 19578 3050
rect 19718 3090 19798 3120
rect 19718 3050 19738 3090
rect 19778 3050 19798 3090
rect 19718 3020 19798 3050
rect 19828 3090 19908 3120
rect 19828 3050 19848 3090
rect 19888 3050 19908 3090
rect 19828 3020 19908 3050
rect 19938 3090 20018 3120
rect 19938 3050 19958 3090
rect 19998 3050 20018 3090
rect 19938 3020 20018 3050
rect 20048 3090 20128 3120
rect 20048 3050 20068 3090
rect 20108 3050 20128 3090
rect 20048 3020 20128 3050
rect 20358 3090 20438 3120
rect 20358 3050 20378 3090
rect 20418 3050 20438 3090
rect 20358 3020 20438 3050
rect 20468 3090 20548 3120
rect 20468 3050 20488 3090
rect 20528 3050 20548 3090
rect 20468 3020 20548 3050
rect 20578 3090 20658 3120
rect 20578 3050 20598 3090
rect 20638 3050 20658 3090
rect 20578 3020 20658 3050
rect 20688 3090 20768 3120
rect 20688 3050 20708 3090
rect 20748 3050 20768 3090
rect 20688 3020 20768 3050
rect 20798 3090 20878 3120
rect 20798 3050 20818 3090
rect 20858 3050 20878 3090
rect 20798 3020 20878 3050
rect 21018 3090 21098 3120
rect 21018 3050 21038 3090
rect 21078 3050 21098 3090
rect 21018 3020 21098 3050
rect 21128 3090 21208 3120
rect 21128 3050 21148 3090
rect 21188 3050 21208 3090
rect 21128 3020 21208 3050
rect 21238 3090 21318 3120
rect 21238 3050 21258 3090
rect 21298 3050 21318 3090
rect 21238 3020 21318 3050
rect 21348 3090 21428 3120
rect 21348 3050 21368 3090
rect 21408 3050 21428 3090
rect 21348 3020 21428 3050
rect 21658 3090 21738 3120
rect 21658 3050 21678 3090
rect 21718 3050 21738 3090
rect 21658 3020 21738 3050
rect 21768 3090 21848 3120
rect 21768 3050 21788 3090
rect 21828 3050 21848 3090
rect 21768 3020 21848 3050
rect 21878 3090 21958 3120
rect 21878 3050 21898 3090
rect 21938 3050 21958 3090
rect 21878 3020 21958 3050
rect 21988 3090 22068 3120
rect 21988 3050 22008 3090
rect 22048 3050 22068 3090
rect 21988 3020 22068 3050
rect 22098 3090 22178 3120
rect 22098 3050 22118 3090
rect 22158 3050 22178 3090
rect 22098 3020 22178 3050
rect 22318 3090 22398 3120
rect 22318 3050 22338 3090
rect 22378 3050 22398 3090
rect 22318 3020 22398 3050
rect 22428 3090 22508 3120
rect 22428 3050 22448 3090
rect 22488 3050 22508 3090
rect 22428 3020 22508 3050
rect 22538 3090 22618 3120
rect 22538 3050 22558 3090
rect 22598 3050 22618 3090
rect 22538 3020 22618 3050
rect 22648 3090 22728 3120
rect 22648 3050 22668 3090
rect 22708 3050 22728 3090
rect 22648 3020 22728 3050
rect 23196 3010 23276 3040
rect 23196 2970 23216 3010
rect 23256 2970 23276 3010
rect 23196 2910 23276 2970
rect 23196 2870 23216 2910
rect 23256 2870 23276 2910
rect 23196 2840 23276 2870
rect 23308 3010 23388 3040
rect 23308 2970 23328 3010
rect 23368 2970 23388 3010
rect 23308 2910 23388 2970
rect 23308 2870 23328 2910
rect 23368 2870 23388 2910
rect 23308 2840 23388 2870
rect 23716 3010 23796 3040
rect 23716 2970 23736 3010
rect 23776 2970 23796 3010
rect 23716 2910 23796 2970
rect 23716 2870 23736 2910
rect 23776 2870 23796 2910
rect 23716 2840 23796 2870
rect 23828 3010 23908 3040
rect 23828 2970 23848 3010
rect 23888 2970 23908 3010
rect 23828 2910 23908 2970
rect 23828 2870 23848 2910
rect 23888 2870 23908 2910
rect 23828 2840 23908 2870
rect 24236 3010 24316 3040
rect 24236 2970 24256 3010
rect 24296 2970 24316 3010
rect 24236 2910 24316 2970
rect 24236 2870 24256 2910
rect 24296 2870 24316 2910
rect 24236 2840 24316 2870
rect 24348 3010 24428 3040
rect 24348 2970 24368 3010
rect 24408 2970 24428 3010
rect 24348 2910 24428 2970
rect 24348 2870 24368 2910
rect 24408 2870 24428 2910
rect 24348 2840 24428 2870
rect 23198 2630 23278 2660
rect 23198 2590 23218 2630
rect 23258 2590 23278 2630
rect 23198 2530 23278 2590
rect 23198 2490 23218 2530
rect 23258 2490 23278 2530
rect 23198 2430 23278 2490
rect 23198 2390 23218 2430
rect 23258 2390 23278 2430
rect 23198 2360 23278 2390
rect 23308 2630 23388 2660
rect 23308 2590 23328 2630
rect 23368 2590 23388 2630
rect 23308 2530 23388 2590
rect 23308 2490 23328 2530
rect 23368 2490 23388 2530
rect 23308 2430 23388 2490
rect 23308 2390 23328 2430
rect 23368 2390 23388 2430
rect 23308 2360 23388 2390
rect 23718 2630 23798 2660
rect 23718 2590 23738 2630
rect 23778 2590 23798 2630
rect 23718 2530 23798 2590
rect 23718 2490 23738 2530
rect 23778 2490 23798 2530
rect 23718 2430 23798 2490
rect 23718 2390 23738 2430
rect 23778 2390 23798 2430
rect 23718 2360 23798 2390
rect 23828 2630 23908 2660
rect 23828 2590 23848 2630
rect 23888 2590 23908 2630
rect 23828 2530 23908 2590
rect 23828 2490 23848 2530
rect 23888 2490 23908 2530
rect 23828 2430 23908 2490
rect 23828 2390 23848 2430
rect 23888 2390 23908 2430
rect 23828 2360 23908 2390
rect 24238 2630 24318 2660
rect 24238 2590 24258 2630
rect 24298 2590 24318 2630
rect 24238 2530 24318 2590
rect 24238 2490 24258 2530
rect 24298 2490 24318 2530
rect 24238 2430 24318 2490
rect 24238 2390 24258 2430
rect 24298 2390 24318 2430
rect 24238 2360 24318 2390
rect 24348 2630 24428 2660
rect 24348 2590 24368 2630
rect 24408 2590 24428 2630
rect 24348 2530 24428 2590
rect 24348 2490 24368 2530
rect 24408 2490 24428 2530
rect 24348 2430 24428 2490
rect 24348 2390 24368 2430
rect 24408 2390 24428 2430
rect 24348 2360 24428 2390
rect 23198 2150 23278 2180
rect 23198 2110 23218 2150
rect 23258 2110 23278 2150
rect 23198 2050 23278 2110
rect 23198 2010 23218 2050
rect 23258 2010 23278 2050
rect 23198 1980 23278 2010
rect 23308 2150 23388 2180
rect 23308 2110 23328 2150
rect 23368 2110 23388 2150
rect 23308 2050 23388 2110
rect 23308 2010 23328 2050
rect 23368 2010 23388 2050
rect 23308 1980 23388 2010
rect 23718 2150 23798 2180
rect 23718 2110 23738 2150
rect 23778 2110 23798 2150
rect 23718 2050 23798 2110
rect 23718 2010 23738 2050
rect 23778 2010 23798 2050
rect 23718 1980 23798 2010
rect 23828 2150 23908 2180
rect 23828 2110 23848 2150
rect 23888 2110 23908 2150
rect 23828 2050 23908 2110
rect 23828 2010 23848 2050
rect 23888 2010 23908 2050
rect 23828 1980 23908 2010
rect 24238 2150 24318 2180
rect 24238 2110 24258 2150
rect 24298 2110 24318 2150
rect 24238 2050 24318 2110
rect 24238 2010 24258 2050
rect 24298 2010 24318 2050
rect 24238 1980 24318 2010
rect 24348 2150 24428 2180
rect 24348 2110 24368 2150
rect 24408 2110 24428 2150
rect 24348 2050 24428 2110
rect 24348 2010 24368 2050
rect 24408 2010 24428 2050
rect 24348 1980 24428 2010
rect 24838 2150 24918 2180
rect 24838 2110 24858 2150
rect 24898 2110 24918 2150
rect 24838 2050 24918 2110
rect 24838 2010 24858 2050
rect 24898 2010 24918 2050
rect 24838 1980 24918 2010
rect 24948 2150 25028 2180
rect 24948 2110 24968 2150
rect 25008 2110 25028 2150
rect 24948 2050 25028 2110
rect 24948 2010 24968 2050
rect 25008 2010 25028 2050
rect 24948 1980 25028 2010
<< pdiff >>
rect 11578 18426 12258 18480
rect 11578 18392 11630 18426
rect 11664 18392 11720 18426
rect 11754 18392 11810 18426
rect 11844 18392 11900 18426
rect 11934 18392 11990 18426
rect 12024 18392 12080 18426
rect 12114 18392 12170 18426
rect 12204 18392 12258 18426
rect 11578 18336 12258 18392
rect 11578 18302 11630 18336
rect 11664 18302 11720 18336
rect 11754 18302 11810 18336
rect 11844 18302 11900 18336
rect 11934 18302 11990 18336
rect 12024 18302 12080 18336
rect 12114 18302 12170 18336
rect 12204 18302 12258 18336
rect 11578 18246 12258 18302
rect 11578 18212 11630 18246
rect 11664 18212 11720 18246
rect 11754 18212 11810 18246
rect 11844 18212 11900 18246
rect 11934 18212 11990 18246
rect 12024 18212 12080 18246
rect 12114 18212 12170 18246
rect 12204 18212 12258 18246
rect 11578 18156 12258 18212
rect 11578 18122 11630 18156
rect 11664 18122 11720 18156
rect 11754 18122 11810 18156
rect 11844 18122 11900 18156
rect 11934 18122 11990 18156
rect 12024 18122 12080 18156
rect 12114 18122 12170 18156
rect 12204 18122 12258 18156
rect 11578 18066 12258 18122
rect 11578 18032 11630 18066
rect 11664 18032 11720 18066
rect 11754 18032 11810 18066
rect 11844 18032 11900 18066
rect 11934 18032 11990 18066
rect 12024 18032 12080 18066
rect 12114 18032 12170 18066
rect 12204 18032 12258 18066
rect 11578 17976 12258 18032
rect 11578 17942 11630 17976
rect 11664 17942 11720 17976
rect 11754 17942 11810 17976
rect 11844 17942 11900 17976
rect 11934 17942 11990 17976
rect 12024 17942 12080 17976
rect 12114 17942 12170 17976
rect 12204 17942 12258 17976
rect 11578 17886 12258 17942
rect 11578 17852 11630 17886
rect 11664 17852 11720 17886
rect 11754 17852 11810 17886
rect 11844 17852 11900 17886
rect 11934 17852 11990 17886
rect 12024 17852 12080 17886
rect 12114 17852 12170 17886
rect 12204 17852 12258 17886
rect 11578 17800 12258 17852
rect 12938 18426 13618 18480
rect 12938 18392 12990 18426
rect 13024 18392 13080 18426
rect 13114 18392 13170 18426
rect 13204 18392 13260 18426
rect 13294 18392 13350 18426
rect 13384 18392 13440 18426
rect 13474 18392 13530 18426
rect 13564 18392 13618 18426
rect 12938 18336 13618 18392
rect 12938 18302 12990 18336
rect 13024 18302 13080 18336
rect 13114 18302 13170 18336
rect 13204 18302 13260 18336
rect 13294 18302 13350 18336
rect 13384 18302 13440 18336
rect 13474 18302 13530 18336
rect 13564 18302 13618 18336
rect 12938 18246 13618 18302
rect 12938 18212 12990 18246
rect 13024 18212 13080 18246
rect 13114 18212 13170 18246
rect 13204 18212 13260 18246
rect 13294 18212 13350 18246
rect 13384 18212 13440 18246
rect 13474 18212 13530 18246
rect 13564 18212 13618 18246
rect 12938 18156 13618 18212
rect 12938 18122 12990 18156
rect 13024 18122 13080 18156
rect 13114 18122 13170 18156
rect 13204 18122 13260 18156
rect 13294 18122 13350 18156
rect 13384 18122 13440 18156
rect 13474 18122 13530 18156
rect 13564 18122 13618 18156
rect 12938 18066 13618 18122
rect 12938 18032 12990 18066
rect 13024 18032 13080 18066
rect 13114 18032 13170 18066
rect 13204 18032 13260 18066
rect 13294 18032 13350 18066
rect 13384 18032 13440 18066
rect 13474 18032 13530 18066
rect 13564 18032 13618 18066
rect 12938 17976 13618 18032
rect 12938 17942 12990 17976
rect 13024 17942 13080 17976
rect 13114 17942 13170 17976
rect 13204 17942 13260 17976
rect 13294 17942 13350 17976
rect 13384 17942 13440 17976
rect 13474 17942 13530 17976
rect 13564 17942 13618 17976
rect 12938 17886 13618 17942
rect 12938 17852 12990 17886
rect 13024 17852 13080 17886
rect 13114 17852 13170 17886
rect 13204 17852 13260 17886
rect 13294 17852 13350 17886
rect 13384 17852 13440 17886
rect 13474 17852 13530 17886
rect 13564 17852 13618 17886
rect 12938 17800 13618 17852
rect 14298 18426 14978 18480
rect 14298 18392 14350 18426
rect 14384 18392 14440 18426
rect 14474 18392 14530 18426
rect 14564 18392 14620 18426
rect 14654 18392 14710 18426
rect 14744 18392 14800 18426
rect 14834 18392 14890 18426
rect 14924 18392 14978 18426
rect 14298 18336 14978 18392
rect 14298 18302 14350 18336
rect 14384 18302 14440 18336
rect 14474 18302 14530 18336
rect 14564 18302 14620 18336
rect 14654 18302 14710 18336
rect 14744 18302 14800 18336
rect 14834 18302 14890 18336
rect 14924 18302 14978 18336
rect 14298 18246 14978 18302
rect 14298 18212 14350 18246
rect 14384 18212 14440 18246
rect 14474 18212 14530 18246
rect 14564 18212 14620 18246
rect 14654 18212 14710 18246
rect 14744 18212 14800 18246
rect 14834 18212 14890 18246
rect 14924 18212 14978 18246
rect 14298 18156 14978 18212
rect 14298 18122 14350 18156
rect 14384 18122 14440 18156
rect 14474 18122 14530 18156
rect 14564 18122 14620 18156
rect 14654 18122 14710 18156
rect 14744 18122 14800 18156
rect 14834 18122 14890 18156
rect 14924 18122 14978 18156
rect 14298 18066 14978 18122
rect 14298 18032 14350 18066
rect 14384 18032 14440 18066
rect 14474 18032 14530 18066
rect 14564 18032 14620 18066
rect 14654 18032 14710 18066
rect 14744 18032 14800 18066
rect 14834 18032 14890 18066
rect 14924 18032 14978 18066
rect 14298 17976 14978 18032
rect 14298 17942 14350 17976
rect 14384 17942 14440 17976
rect 14474 17942 14530 17976
rect 14564 17942 14620 17976
rect 14654 17942 14710 17976
rect 14744 17942 14800 17976
rect 14834 17942 14890 17976
rect 14924 17942 14978 17976
rect 14298 17886 14978 17942
rect 14298 17852 14350 17886
rect 14384 17852 14440 17886
rect 14474 17852 14530 17886
rect 14564 17852 14620 17886
rect 14654 17852 14710 17886
rect 14744 17852 14800 17886
rect 14834 17852 14890 17886
rect 14924 17852 14978 17886
rect 14298 17800 14978 17852
rect 11578 17066 12258 17120
rect 11578 17032 11630 17066
rect 11664 17032 11720 17066
rect 11754 17032 11810 17066
rect 11844 17032 11900 17066
rect 11934 17032 11990 17066
rect 12024 17032 12080 17066
rect 12114 17032 12170 17066
rect 12204 17032 12258 17066
rect 11578 16976 12258 17032
rect 11578 16942 11630 16976
rect 11664 16942 11720 16976
rect 11754 16942 11810 16976
rect 11844 16942 11900 16976
rect 11934 16942 11990 16976
rect 12024 16942 12080 16976
rect 12114 16942 12170 16976
rect 12204 16942 12258 16976
rect 11578 16886 12258 16942
rect 11578 16852 11630 16886
rect 11664 16852 11720 16886
rect 11754 16852 11810 16886
rect 11844 16852 11900 16886
rect 11934 16852 11990 16886
rect 12024 16852 12080 16886
rect 12114 16852 12170 16886
rect 12204 16852 12258 16886
rect 11578 16796 12258 16852
rect 11578 16762 11630 16796
rect 11664 16762 11720 16796
rect 11754 16762 11810 16796
rect 11844 16762 11900 16796
rect 11934 16762 11990 16796
rect 12024 16762 12080 16796
rect 12114 16762 12170 16796
rect 12204 16762 12258 16796
rect 11578 16706 12258 16762
rect 11578 16672 11630 16706
rect 11664 16672 11720 16706
rect 11754 16672 11810 16706
rect 11844 16672 11900 16706
rect 11934 16672 11990 16706
rect 12024 16672 12080 16706
rect 12114 16672 12170 16706
rect 12204 16672 12258 16706
rect 11578 16616 12258 16672
rect 11578 16582 11630 16616
rect 11664 16582 11720 16616
rect 11754 16582 11810 16616
rect 11844 16582 11900 16616
rect 11934 16582 11990 16616
rect 12024 16582 12080 16616
rect 12114 16582 12170 16616
rect 12204 16582 12258 16616
rect 11578 16526 12258 16582
rect 11578 16492 11630 16526
rect 11664 16492 11720 16526
rect 11754 16492 11810 16526
rect 11844 16492 11900 16526
rect 11934 16492 11990 16526
rect 12024 16492 12080 16526
rect 12114 16492 12170 16526
rect 12204 16492 12258 16526
rect 11578 16440 12258 16492
rect 12938 17066 13618 17120
rect 12938 17032 12990 17066
rect 13024 17032 13080 17066
rect 13114 17032 13170 17066
rect 13204 17032 13260 17066
rect 13294 17032 13350 17066
rect 13384 17032 13440 17066
rect 13474 17032 13530 17066
rect 13564 17032 13618 17066
rect 12938 16976 13618 17032
rect 12938 16942 12990 16976
rect 13024 16942 13080 16976
rect 13114 16942 13170 16976
rect 13204 16942 13260 16976
rect 13294 16942 13350 16976
rect 13384 16942 13440 16976
rect 13474 16942 13530 16976
rect 13564 16942 13618 16976
rect 12938 16886 13618 16942
rect 12938 16852 12990 16886
rect 13024 16852 13080 16886
rect 13114 16852 13170 16886
rect 13204 16852 13260 16886
rect 13294 16852 13350 16886
rect 13384 16852 13440 16886
rect 13474 16852 13530 16886
rect 13564 16852 13618 16886
rect 12938 16796 13618 16852
rect 12938 16762 12990 16796
rect 13024 16762 13080 16796
rect 13114 16762 13170 16796
rect 13204 16762 13260 16796
rect 13294 16762 13350 16796
rect 13384 16762 13440 16796
rect 13474 16762 13530 16796
rect 13564 16762 13618 16796
rect 12938 16706 13618 16762
rect 12938 16672 12990 16706
rect 13024 16672 13080 16706
rect 13114 16672 13170 16706
rect 13204 16672 13260 16706
rect 13294 16672 13350 16706
rect 13384 16672 13440 16706
rect 13474 16672 13530 16706
rect 13564 16672 13618 16706
rect 12938 16616 13618 16672
rect 12938 16582 12990 16616
rect 13024 16582 13080 16616
rect 13114 16582 13170 16616
rect 13204 16582 13260 16616
rect 13294 16582 13350 16616
rect 13384 16582 13440 16616
rect 13474 16582 13530 16616
rect 13564 16582 13618 16616
rect 12938 16526 13618 16582
rect 12938 16492 12990 16526
rect 13024 16492 13080 16526
rect 13114 16492 13170 16526
rect 13204 16492 13260 16526
rect 13294 16492 13350 16526
rect 13384 16492 13440 16526
rect 13474 16492 13530 16526
rect 13564 16492 13618 16526
rect 12938 16440 13618 16492
rect 14298 17066 14978 17120
rect 14298 17032 14350 17066
rect 14384 17032 14440 17066
rect 14474 17032 14530 17066
rect 14564 17032 14620 17066
rect 14654 17032 14710 17066
rect 14744 17032 14800 17066
rect 14834 17032 14890 17066
rect 14924 17032 14978 17066
rect 14298 16976 14978 17032
rect 14298 16942 14350 16976
rect 14384 16942 14440 16976
rect 14474 16942 14530 16976
rect 14564 16942 14620 16976
rect 14654 16942 14710 16976
rect 14744 16942 14800 16976
rect 14834 16942 14890 16976
rect 14924 16942 14978 16976
rect 14298 16886 14978 16942
rect 14298 16852 14350 16886
rect 14384 16852 14440 16886
rect 14474 16852 14530 16886
rect 14564 16852 14620 16886
rect 14654 16852 14710 16886
rect 14744 16852 14800 16886
rect 14834 16852 14890 16886
rect 14924 16852 14978 16886
rect 14298 16796 14978 16852
rect 14298 16762 14350 16796
rect 14384 16762 14440 16796
rect 14474 16762 14530 16796
rect 14564 16762 14620 16796
rect 14654 16762 14710 16796
rect 14744 16762 14800 16796
rect 14834 16762 14890 16796
rect 14924 16762 14978 16796
rect 14298 16706 14978 16762
rect 14298 16672 14350 16706
rect 14384 16672 14440 16706
rect 14474 16672 14530 16706
rect 14564 16672 14620 16706
rect 14654 16672 14710 16706
rect 14744 16672 14800 16706
rect 14834 16672 14890 16706
rect 14924 16672 14978 16706
rect 14298 16616 14978 16672
rect 14298 16582 14350 16616
rect 14384 16582 14440 16616
rect 14474 16582 14530 16616
rect 14564 16582 14620 16616
rect 14654 16582 14710 16616
rect 14744 16582 14800 16616
rect 14834 16582 14890 16616
rect 14924 16582 14978 16616
rect 14298 16526 14978 16582
rect 14298 16492 14350 16526
rect 14384 16492 14440 16526
rect 14474 16492 14530 16526
rect 14564 16492 14620 16526
rect 14654 16492 14710 16526
rect 14744 16492 14800 16526
rect 14834 16492 14890 16526
rect 14924 16492 14978 16526
rect 14298 16440 14978 16492
rect 11578 15706 12258 15760
rect 11578 15672 11630 15706
rect 11664 15672 11720 15706
rect 11754 15672 11810 15706
rect 11844 15672 11900 15706
rect 11934 15672 11990 15706
rect 12024 15672 12080 15706
rect 12114 15672 12170 15706
rect 12204 15672 12258 15706
rect 11578 15616 12258 15672
rect 11578 15582 11630 15616
rect 11664 15582 11720 15616
rect 11754 15582 11810 15616
rect 11844 15582 11900 15616
rect 11934 15582 11990 15616
rect 12024 15582 12080 15616
rect 12114 15582 12170 15616
rect 12204 15582 12258 15616
rect 11578 15526 12258 15582
rect 11578 15492 11630 15526
rect 11664 15492 11720 15526
rect 11754 15492 11810 15526
rect 11844 15492 11900 15526
rect 11934 15492 11990 15526
rect 12024 15492 12080 15526
rect 12114 15492 12170 15526
rect 12204 15492 12258 15526
rect 11578 15436 12258 15492
rect 11578 15402 11630 15436
rect 11664 15402 11720 15436
rect 11754 15402 11810 15436
rect 11844 15402 11900 15436
rect 11934 15402 11990 15436
rect 12024 15402 12080 15436
rect 12114 15402 12170 15436
rect 12204 15402 12258 15436
rect 11578 15346 12258 15402
rect 11578 15312 11630 15346
rect 11664 15312 11720 15346
rect 11754 15312 11810 15346
rect 11844 15312 11900 15346
rect 11934 15312 11990 15346
rect 12024 15312 12080 15346
rect 12114 15312 12170 15346
rect 12204 15312 12258 15346
rect 11578 15256 12258 15312
rect 11578 15222 11630 15256
rect 11664 15222 11720 15256
rect 11754 15222 11810 15256
rect 11844 15222 11900 15256
rect 11934 15222 11990 15256
rect 12024 15222 12080 15256
rect 12114 15222 12170 15256
rect 12204 15222 12258 15256
rect 11578 15166 12258 15222
rect 11578 15132 11630 15166
rect 11664 15132 11720 15166
rect 11754 15132 11810 15166
rect 11844 15132 11900 15166
rect 11934 15132 11990 15166
rect 12024 15132 12080 15166
rect 12114 15132 12170 15166
rect 12204 15132 12258 15166
rect 11578 15080 12258 15132
rect 12938 15706 13618 15760
rect 12938 15672 12990 15706
rect 13024 15672 13080 15706
rect 13114 15672 13170 15706
rect 13204 15672 13260 15706
rect 13294 15672 13350 15706
rect 13384 15672 13440 15706
rect 13474 15672 13530 15706
rect 13564 15672 13618 15706
rect 12938 15616 13618 15672
rect 12938 15582 12990 15616
rect 13024 15582 13080 15616
rect 13114 15582 13170 15616
rect 13204 15582 13260 15616
rect 13294 15582 13350 15616
rect 13384 15582 13440 15616
rect 13474 15582 13530 15616
rect 13564 15582 13618 15616
rect 12938 15526 13618 15582
rect 12938 15492 12990 15526
rect 13024 15492 13080 15526
rect 13114 15492 13170 15526
rect 13204 15492 13260 15526
rect 13294 15492 13350 15526
rect 13384 15492 13440 15526
rect 13474 15492 13530 15526
rect 13564 15492 13618 15526
rect 12938 15436 13618 15492
rect 12938 15402 12990 15436
rect 13024 15402 13080 15436
rect 13114 15402 13170 15436
rect 13204 15402 13260 15436
rect 13294 15402 13350 15436
rect 13384 15402 13440 15436
rect 13474 15402 13530 15436
rect 13564 15402 13618 15436
rect 12938 15346 13618 15402
rect 12938 15312 12990 15346
rect 13024 15312 13080 15346
rect 13114 15312 13170 15346
rect 13204 15312 13260 15346
rect 13294 15312 13350 15346
rect 13384 15312 13440 15346
rect 13474 15312 13530 15346
rect 13564 15312 13618 15346
rect 12938 15256 13618 15312
rect 12938 15222 12990 15256
rect 13024 15222 13080 15256
rect 13114 15222 13170 15256
rect 13204 15222 13260 15256
rect 13294 15222 13350 15256
rect 13384 15222 13440 15256
rect 13474 15222 13530 15256
rect 13564 15222 13618 15256
rect 12938 15166 13618 15222
rect 12938 15132 12990 15166
rect 13024 15132 13080 15166
rect 13114 15132 13170 15166
rect 13204 15132 13260 15166
rect 13294 15132 13350 15166
rect 13384 15132 13440 15166
rect 13474 15132 13530 15166
rect 13564 15132 13618 15166
rect 12938 15080 13618 15132
rect 14298 15706 14978 15760
rect 14298 15672 14350 15706
rect 14384 15672 14440 15706
rect 14474 15672 14530 15706
rect 14564 15672 14620 15706
rect 14654 15672 14710 15706
rect 14744 15672 14800 15706
rect 14834 15672 14890 15706
rect 14924 15672 14978 15706
rect 14298 15616 14978 15672
rect 14298 15582 14350 15616
rect 14384 15582 14440 15616
rect 14474 15582 14530 15616
rect 14564 15582 14620 15616
rect 14654 15582 14710 15616
rect 14744 15582 14800 15616
rect 14834 15582 14890 15616
rect 14924 15582 14978 15616
rect 14298 15526 14978 15582
rect 14298 15492 14350 15526
rect 14384 15492 14440 15526
rect 14474 15492 14530 15526
rect 14564 15492 14620 15526
rect 14654 15492 14710 15526
rect 14744 15492 14800 15526
rect 14834 15492 14890 15526
rect 14924 15492 14978 15526
rect 14298 15436 14978 15492
rect 14298 15402 14350 15436
rect 14384 15402 14440 15436
rect 14474 15402 14530 15436
rect 14564 15402 14620 15436
rect 14654 15402 14710 15436
rect 14744 15402 14800 15436
rect 14834 15402 14890 15436
rect 14924 15402 14978 15436
rect 14298 15346 14978 15402
rect 14298 15312 14350 15346
rect 14384 15312 14440 15346
rect 14474 15312 14530 15346
rect 14564 15312 14620 15346
rect 14654 15312 14710 15346
rect 14744 15312 14800 15346
rect 14834 15312 14890 15346
rect 14924 15312 14978 15346
rect 14298 15256 14978 15312
rect 14298 15222 14350 15256
rect 14384 15222 14440 15256
rect 14474 15222 14530 15256
rect 14564 15222 14620 15256
rect 14654 15222 14710 15256
rect 14744 15222 14800 15256
rect 14834 15222 14890 15256
rect 14924 15222 14978 15256
rect 14298 15166 14978 15222
rect 14298 15132 14350 15166
rect 14384 15132 14440 15166
rect 14474 15132 14530 15166
rect 14564 15132 14620 15166
rect 14654 15132 14710 15166
rect 14744 15132 14800 15166
rect 14834 15132 14890 15166
rect 14924 15132 14978 15166
rect 14298 15080 14978 15132
rect 19508 12660 19608 12690
rect 19508 12620 19538 12660
rect 19578 12620 19608 12660
rect 19508 12560 19608 12620
rect 19508 12520 19538 12560
rect 19578 12520 19608 12560
rect 19508 12460 19608 12520
rect 19508 12420 19538 12460
rect 19578 12420 19608 12460
rect 19508 12360 19608 12420
rect 19508 12320 19538 12360
rect 19578 12320 19608 12360
rect 19508 12260 19608 12320
rect 19508 12220 19538 12260
rect 19578 12220 19608 12260
rect 19508 12190 19608 12220
rect 19708 12660 19808 12690
rect 19708 12620 19738 12660
rect 19778 12620 19808 12660
rect 19708 12560 19808 12620
rect 19708 12520 19738 12560
rect 19778 12520 19808 12560
rect 19708 12460 19808 12520
rect 19708 12420 19738 12460
rect 19778 12420 19808 12460
rect 19708 12360 19808 12420
rect 19708 12320 19738 12360
rect 19778 12320 19808 12360
rect 19708 12260 19808 12320
rect 19708 12220 19738 12260
rect 19778 12220 19808 12260
rect 19708 12190 19808 12220
rect 19908 12660 20008 12690
rect 19908 12620 19938 12660
rect 19978 12620 20008 12660
rect 19908 12560 20008 12620
rect 19908 12520 19938 12560
rect 19978 12520 20008 12560
rect 19908 12460 20008 12520
rect 19908 12420 19938 12460
rect 19978 12420 20008 12460
rect 19908 12360 20008 12420
rect 19908 12320 19938 12360
rect 19978 12320 20008 12360
rect 19908 12260 20008 12320
rect 19908 12220 19938 12260
rect 19978 12220 20008 12260
rect 19908 12190 20008 12220
rect 20108 12660 20208 12690
rect 20108 12620 20138 12660
rect 20178 12620 20208 12660
rect 20108 12560 20208 12620
rect 20108 12520 20138 12560
rect 20178 12520 20208 12560
rect 20108 12460 20208 12520
rect 20108 12420 20138 12460
rect 20178 12420 20208 12460
rect 20108 12360 20208 12420
rect 20108 12320 20138 12360
rect 20178 12320 20208 12360
rect 20108 12260 20208 12320
rect 20108 12220 20138 12260
rect 20178 12220 20208 12260
rect 20108 12190 20208 12220
rect 20308 12660 20408 12690
rect 20308 12620 20338 12660
rect 20378 12620 20408 12660
rect 20308 12560 20408 12620
rect 20308 12520 20338 12560
rect 20378 12520 20408 12560
rect 20308 12460 20408 12520
rect 20308 12420 20338 12460
rect 20378 12420 20408 12460
rect 20308 12360 20408 12420
rect 20308 12320 20338 12360
rect 20378 12320 20408 12360
rect 20308 12260 20408 12320
rect 20308 12220 20338 12260
rect 20378 12220 20408 12260
rect 20308 12190 20408 12220
rect 20508 12660 20608 12690
rect 20508 12620 20538 12660
rect 20578 12620 20608 12660
rect 20508 12560 20608 12620
rect 20508 12520 20538 12560
rect 20578 12520 20608 12560
rect 20508 12460 20608 12520
rect 20508 12420 20538 12460
rect 20578 12420 20608 12460
rect 20508 12360 20608 12420
rect 20508 12320 20538 12360
rect 20578 12320 20608 12360
rect 20508 12260 20608 12320
rect 20508 12220 20538 12260
rect 20578 12220 20608 12260
rect 20508 12190 20608 12220
rect 20708 12660 20808 12690
rect 20708 12620 20738 12660
rect 20778 12620 20808 12660
rect 20708 12560 20808 12620
rect 20708 12520 20738 12560
rect 20778 12520 20808 12560
rect 20708 12460 20808 12520
rect 20708 12420 20738 12460
rect 20778 12420 20808 12460
rect 20708 12360 20808 12420
rect 20708 12320 20738 12360
rect 20778 12320 20808 12360
rect 20708 12260 20808 12320
rect 20708 12220 20738 12260
rect 20778 12220 20808 12260
rect 20708 12190 20808 12220
rect 20908 12660 21008 12690
rect 20908 12620 20938 12660
rect 20978 12620 21008 12660
rect 20908 12560 21008 12620
rect 20908 12520 20938 12560
rect 20978 12520 21008 12560
rect 20908 12460 21008 12520
rect 20908 12420 20938 12460
rect 20978 12420 21008 12460
rect 20908 12360 21008 12420
rect 20908 12320 20938 12360
rect 20978 12320 21008 12360
rect 20908 12260 21008 12320
rect 20908 12220 20938 12260
rect 20978 12220 21008 12260
rect 20908 12190 21008 12220
rect 21108 12660 21208 12690
rect 21108 12620 21138 12660
rect 21178 12620 21208 12660
rect 21108 12560 21208 12620
rect 21108 12520 21138 12560
rect 21178 12520 21208 12560
rect 21108 12460 21208 12520
rect 21108 12420 21138 12460
rect 21178 12420 21208 12460
rect 21108 12360 21208 12420
rect 21108 12320 21138 12360
rect 21178 12320 21208 12360
rect 21108 12260 21208 12320
rect 21108 12220 21138 12260
rect 21178 12220 21208 12260
rect 21108 12190 21208 12220
rect 21308 12660 21408 12690
rect 21308 12620 21338 12660
rect 21378 12620 21408 12660
rect 21308 12560 21408 12620
rect 21308 12520 21338 12560
rect 21378 12520 21408 12560
rect 21308 12460 21408 12520
rect 21308 12420 21338 12460
rect 21378 12420 21408 12460
rect 21308 12360 21408 12420
rect 21308 12320 21338 12360
rect 21378 12320 21408 12360
rect 21308 12260 21408 12320
rect 21308 12220 21338 12260
rect 21378 12220 21408 12260
rect 21308 12190 21408 12220
rect 21508 12660 21608 12690
rect 21508 12620 21538 12660
rect 21578 12620 21608 12660
rect 21508 12560 21608 12620
rect 21508 12520 21538 12560
rect 21578 12520 21608 12560
rect 21508 12460 21608 12520
rect 21508 12420 21538 12460
rect 21578 12420 21608 12460
rect 21508 12360 21608 12420
rect 21508 12320 21538 12360
rect 21578 12320 21608 12360
rect 21508 12260 21608 12320
rect 21508 12220 21538 12260
rect 21578 12220 21608 12260
rect 21508 12190 21608 12220
rect 10518 11790 10598 11820
rect 10518 11750 10538 11790
rect 10578 11750 10598 11790
rect 10518 11690 10598 11750
rect 10518 11650 10538 11690
rect 10578 11650 10598 11690
rect 10518 11620 10598 11650
rect 10638 11790 10718 11820
rect 10638 11750 10658 11790
rect 10698 11750 10718 11790
rect 10638 11690 10718 11750
rect 10638 11650 10658 11690
rect 10698 11650 10718 11690
rect 10638 11620 10718 11650
rect 10758 11790 10838 11820
rect 10758 11750 10778 11790
rect 10818 11750 10838 11790
rect 10758 11690 10838 11750
rect 10758 11650 10778 11690
rect 10818 11650 10838 11690
rect 10758 11620 10838 11650
rect 10878 11790 10958 11820
rect 10878 11750 10898 11790
rect 10938 11750 10958 11790
rect 10878 11690 10958 11750
rect 10878 11650 10898 11690
rect 10938 11650 10958 11690
rect 10878 11620 10958 11650
rect 10998 11790 11078 11820
rect 10998 11750 11018 11790
rect 11058 11750 11078 11790
rect 10998 11690 11078 11750
rect 10998 11650 11018 11690
rect 11058 11650 11078 11690
rect 10998 11620 11078 11650
rect 11118 11790 11198 11820
rect 11118 11750 11138 11790
rect 11178 11750 11198 11790
rect 11118 11690 11198 11750
rect 11118 11650 11138 11690
rect 11178 11650 11198 11690
rect 11118 11620 11198 11650
rect 11238 11790 11318 11820
rect 11238 11750 11258 11790
rect 11298 11750 11318 11790
rect 11238 11690 11318 11750
rect 11238 11650 11258 11690
rect 11298 11650 11318 11690
rect 11238 11620 11318 11650
rect 11358 11790 11438 11820
rect 11358 11750 11378 11790
rect 11418 11750 11438 11790
rect 11358 11690 11438 11750
rect 11358 11650 11378 11690
rect 11418 11650 11438 11690
rect 11358 11620 11438 11650
rect 11478 11790 11558 11820
rect 11478 11750 11498 11790
rect 11538 11750 11558 11790
rect 11478 11690 11558 11750
rect 11478 11650 11498 11690
rect 11538 11650 11558 11690
rect 11478 11620 11558 11650
rect 11598 11790 11678 11820
rect 11598 11750 11618 11790
rect 11658 11750 11678 11790
rect 11598 11690 11678 11750
rect 11598 11650 11618 11690
rect 11658 11650 11678 11690
rect 11598 11620 11678 11650
rect 11718 11790 11798 11820
rect 11718 11750 11738 11790
rect 11778 11750 11798 11790
rect 11718 11690 11798 11750
rect 11718 11650 11738 11690
rect 11778 11650 11798 11690
rect 11718 11620 11798 11650
rect 11838 11790 11918 11820
rect 11838 11750 11858 11790
rect 11898 11750 11918 11790
rect 11838 11690 11918 11750
rect 11838 11650 11858 11690
rect 11898 11650 11918 11690
rect 11838 11620 11918 11650
rect 11958 11790 12038 11820
rect 11958 11750 11978 11790
rect 12018 11750 12038 11790
rect 11958 11690 12038 11750
rect 11958 11650 11978 11690
rect 12018 11650 12038 11690
rect 11958 11620 12038 11650
rect 12078 11790 12158 11820
rect 12078 11750 12098 11790
rect 12138 11750 12158 11790
rect 12078 11690 12158 11750
rect 12078 11650 12098 11690
rect 12138 11650 12158 11690
rect 12078 11620 12158 11650
rect 12198 11790 12278 11820
rect 12198 11750 12218 11790
rect 12258 11750 12278 11790
rect 12198 11690 12278 11750
rect 12198 11650 12218 11690
rect 12258 11650 12278 11690
rect 12198 11620 12278 11650
rect 12318 11790 12398 11820
rect 12318 11750 12338 11790
rect 12378 11750 12398 11790
rect 12318 11690 12398 11750
rect 12318 11650 12338 11690
rect 12378 11650 12398 11690
rect 12318 11620 12398 11650
rect 12438 11790 12518 11820
rect 12438 11750 12458 11790
rect 12498 11750 12518 11790
rect 12438 11690 12518 11750
rect 12438 11650 12458 11690
rect 12498 11650 12518 11690
rect 12438 11620 12518 11650
rect 12558 11790 12638 11820
rect 12558 11750 12578 11790
rect 12618 11750 12638 11790
rect 12558 11690 12638 11750
rect 12558 11650 12578 11690
rect 12618 11650 12638 11690
rect 12558 11620 12638 11650
rect 12678 11790 12758 11820
rect 12678 11750 12698 11790
rect 12738 11750 12758 11790
rect 12678 11690 12758 11750
rect 12678 11650 12698 11690
rect 12738 11650 12758 11690
rect 12678 11620 12758 11650
rect 12798 11790 12878 11820
rect 12798 11750 12818 11790
rect 12858 11750 12878 11790
rect 12798 11690 12878 11750
rect 12798 11650 12818 11690
rect 12858 11650 12878 11690
rect 12798 11620 12878 11650
rect 12918 11790 12998 11820
rect 12918 11750 12938 11790
rect 12978 11750 12998 11790
rect 12918 11690 12998 11750
rect 12918 11650 12938 11690
rect 12978 11650 12998 11690
rect 12918 11620 12998 11650
rect 13558 11790 13638 11820
rect 13558 11750 13578 11790
rect 13618 11750 13638 11790
rect 13558 11690 13638 11750
rect 13558 11650 13578 11690
rect 13618 11650 13638 11690
rect 13558 11620 13638 11650
rect 13678 11790 13758 11820
rect 13678 11750 13698 11790
rect 13738 11750 13758 11790
rect 13678 11690 13758 11750
rect 13678 11650 13698 11690
rect 13738 11650 13758 11690
rect 13678 11620 13758 11650
rect 13798 11790 13878 11820
rect 13798 11750 13818 11790
rect 13858 11750 13878 11790
rect 13798 11690 13878 11750
rect 13798 11650 13818 11690
rect 13858 11650 13878 11690
rect 13798 11620 13878 11650
rect 13918 11790 13998 11820
rect 13918 11750 13938 11790
rect 13978 11750 13998 11790
rect 13918 11690 13998 11750
rect 13918 11650 13938 11690
rect 13978 11650 13998 11690
rect 13918 11620 13998 11650
rect 14038 11790 14118 11820
rect 14038 11750 14058 11790
rect 14098 11750 14118 11790
rect 14038 11690 14118 11750
rect 14038 11650 14058 11690
rect 14098 11650 14118 11690
rect 14038 11620 14118 11650
rect 14158 11790 14238 11820
rect 14158 11750 14178 11790
rect 14218 11750 14238 11790
rect 14158 11690 14238 11750
rect 14158 11650 14178 11690
rect 14218 11650 14238 11690
rect 14158 11620 14238 11650
rect 14278 11790 14358 11820
rect 14278 11750 14298 11790
rect 14338 11750 14358 11790
rect 14278 11690 14358 11750
rect 14278 11650 14298 11690
rect 14338 11650 14358 11690
rect 14278 11620 14358 11650
rect 14398 11790 14478 11820
rect 14398 11750 14418 11790
rect 14458 11750 14478 11790
rect 14398 11690 14478 11750
rect 14398 11650 14418 11690
rect 14458 11650 14478 11690
rect 14398 11620 14478 11650
rect 14518 11790 14598 11820
rect 14518 11750 14538 11790
rect 14578 11750 14598 11790
rect 14518 11690 14598 11750
rect 14518 11650 14538 11690
rect 14578 11650 14598 11690
rect 14518 11620 14598 11650
rect 14638 11790 14718 11820
rect 14638 11750 14658 11790
rect 14698 11750 14718 11790
rect 14638 11690 14718 11750
rect 14638 11650 14658 11690
rect 14698 11650 14718 11690
rect 14638 11620 14718 11650
rect 14758 11790 14838 11820
rect 14758 11750 14778 11790
rect 14818 11750 14838 11790
rect 14758 11690 14838 11750
rect 14758 11650 14778 11690
rect 14818 11650 14838 11690
rect 14758 11620 14838 11650
rect 14878 11790 14958 11820
rect 14878 11750 14898 11790
rect 14938 11750 14958 11790
rect 14878 11690 14958 11750
rect 14878 11650 14898 11690
rect 14938 11650 14958 11690
rect 14878 11620 14958 11650
rect 14998 11790 15078 11820
rect 14998 11750 15018 11790
rect 15058 11750 15078 11790
rect 14998 11690 15078 11750
rect 14998 11650 15018 11690
rect 15058 11650 15078 11690
rect 14998 11620 15078 11650
rect 15118 11790 15198 11820
rect 15118 11750 15138 11790
rect 15178 11750 15198 11790
rect 15118 11690 15198 11750
rect 15118 11650 15138 11690
rect 15178 11650 15198 11690
rect 15118 11620 15198 11650
rect 15238 11790 15318 11820
rect 15238 11750 15258 11790
rect 15298 11750 15318 11790
rect 15238 11690 15318 11750
rect 15238 11650 15258 11690
rect 15298 11650 15318 11690
rect 15238 11620 15318 11650
rect 15358 11790 15438 11820
rect 15358 11750 15378 11790
rect 15418 11750 15438 11790
rect 15358 11690 15438 11750
rect 15358 11650 15378 11690
rect 15418 11650 15438 11690
rect 15358 11620 15438 11650
rect 15478 11790 15558 11820
rect 15478 11750 15498 11790
rect 15538 11750 15558 11790
rect 15478 11690 15558 11750
rect 15478 11650 15498 11690
rect 15538 11650 15558 11690
rect 15478 11620 15558 11650
rect 15598 11790 15678 11820
rect 15598 11750 15618 11790
rect 15658 11750 15678 11790
rect 15598 11690 15678 11750
rect 15598 11650 15618 11690
rect 15658 11650 15678 11690
rect 15598 11620 15678 11650
rect 15718 11790 15798 11820
rect 15718 11750 15738 11790
rect 15778 11750 15798 11790
rect 15718 11690 15798 11750
rect 15718 11650 15738 11690
rect 15778 11650 15798 11690
rect 15718 11620 15798 11650
rect 15838 11790 15918 11820
rect 15838 11750 15858 11790
rect 15898 11750 15918 11790
rect 15838 11690 15918 11750
rect 15838 11650 15858 11690
rect 15898 11650 15918 11690
rect 15838 11620 15918 11650
rect 15958 11790 16038 11820
rect 15958 11750 15978 11790
rect 16018 11750 16038 11790
rect 15958 11690 16038 11750
rect 15958 11650 15978 11690
rect 16018 11650 16038 11690
rect 15958 11620 16038 11650
rect 19438 11710 19538 11740
rect 19438 11670 19468 11710
rect 19508 11670 19538 11710
rect 19438 11610 19538 11670
rect 19438 11570 19468 11610
rect 19508 11570 19538 11610
rect 19438 11540 19538 11570
rect 19568 11710 19668 11740
rect 19568 11670 19598 11710
rect 19638 11670 19668 11710
rect 19568 11610 19668 11670
rect 19568 11570 19598 11610
rect 19638 11570 19668 11610
rect 19568 11540 19668 11570
rect 19698 11710 19798 11740
rect 19698 11670 19728 11710
rect 19768 11670 19798 11710
rect 19698 11610 19798 11670
rect 19698 11570 19728 11610
rect 19768 11570 19798 11610
rect 19698 11540 19798 11570
rect 19828 11710 19928 11740
rect 19828 11670 19858 11710
rect 19898 11670 19928 11710
rect 19828 11610 19928 11670
rect 19828 11570 19858 11610
rect 19898 11570 19928 11610
rect 19828 11540 19928 11570
rect 19958 11710 20058 11740
rect 19958 11670 19988 11710
rect 20028 11670 20058 11710
rect 19958 11610 20058 11670
rect 19958 11570 19988 11610
rect 20028 11570 20058 11610
rect 19958 11540 20058 11570
rect 20088 11710 20188 11740
rect 20088 11670 20118 11710
rect 20158 11670 20188 11710
rect 20088 11610 20188 11670
rect 20088 11570 20118 11610
rect 20158 11570 20188 11610
rect 20088 11540 20188 11570
rect 20218 11710 20318 11740
rect 20218 11670 20248 11710
rect 20288 11670 20318 11710
rect 20218 11610 20318 11670
rect 20218 11570 20248 11610
rect 20288 11570 20318 11610
rect 20218 11540 20318 11570
rect 20578 11710 20678 11740
rect 20578 11670 20608 11710
rect 20648 11670 20678 11710
rect 20578 11610 20678 11670
rect 20578 11570 20608 11610
rect 20648 11570 20678 11610
rect 20578 11540 20678 11570
rect 20708 11710 20808 11740
rect 20708 11670 20738 11710
rect 20778 11670 20808 11710
rect 20708 11610 20808 11670
rect 20708 11570 20738 11610
rect 20778 11570 20808 11610
rect 20708 11540 20808 11570
rect 20838 11710 20938 11740
rect 20838 11670 20868 11710
rect 20908 11670 20938 11710
rect 20838 11610 20938 11670
rect 20838 11570 20868 11610
rect 20908 11570 20938 11610
rect 20838 11540 20938 11570
rect 20968 11710 21068 11740
rect 20968 11670 20998 11710
rect 21038 11670 21068 11710
rect 20968 11610 21068 11670
rect 20968 11570 20998 11610
rect 21038 11570 21068 11610
rect 20968 11540 21068 11570
rect 21098 11710 21198 11740
rect 21098 11670 21128 11710
rect 21168 11670 21198 11710
rect 21098 11610 21198 11670
rect 21098 11570 21128 11610
rect 21168 11570 21198 11610
rect 21098 11540 21198 11570
rect 21228 11710 21328 11740
rect 21228 11670 21258 11710
rect 21298 11670 21328 11710
rect 21228 11610 21328 11670
rect 21228 11570 21258 11610
rect 21298 11570 21328 11610
rect 21228 11540 21328 11570
rect 21358 11710 21458 11740
rect 21358 11670 21388 11710
rect 21428 11670 21458 11710
rect 21358 11610 21458 11670
rect 21358 11570 21388 11610
rect 21428 11570 21458 11610
rect 21358 11540 21458 11570
rect 21718 11710 21818 11740
rect 21718 11670 21748 11710
rect 21788 11670 21818 11710
rect 21718 11610 21818 11670
rect 21718 11570 21748 11610
rect 21788 11570 21818 11610
rect 21718 11540 21818 11570
rect 21848 11710 21948 11740
rect 21848 11670 21878 11710
rect 21918 11670 21948 11710
rect 21848 11610 21948 11670
rect 21848 11570 21878 11610
rect 21918 11570 21948 11610
rect 21848 11540 21948 11570
rect 21978 11710 22078 11740
rect 21978 11670 22008 11710
rect 22048 11670 22078 11710
rect 21978 11610 22078 11670
rect 21978 11570 22008 11610
rect 22048 11570 22078 11610
rect 21978 11540 22078 11570
rect 22108 11710 22208 11740
rect 22108 11670 22138 11710
rect 22178 11670 22208 11710
rect 22108 11610 22208 11670
rect 22108 11570 22138 11610
rect 22178 11570 22208 11610
rect 22108 11540 22208 11570
rect 22238 11710 22338 11740
rect 22238 11670 22268 11710
rect 22308 11670 22338 11710
rect 22238 11610 22338 11670
rect 22238 11570 22268 11610
rect 22308 11570 22338 11610
rect 22238 11540 22338 11570
rect 22368 11710 22468 11740
rect 22368 11670 22398 11710
rect 22438 11670 22468 11710
rect 22368 11610 22468 11670
rect 22368 11570 22398 11610
rect 22438 11570 22468 11610
rect 22368 11540 22468 11570
rect 22498 11710 22598 11740
rect 22498 11670 22528 11710
rect 22568 11670 22598 11710
rect 22498 11610 22598 11670
rect 22498 11570 22528 11610
rect 22568 11570 22598 11610
rect 22498 11540 22598 11570
rect 11618 10630 11698 10660
rect 11618 10590 11638 10630
rect 11678 10590 11698 10630
rect 11618 10530 11698 10590
rect 11618 10490 11638 10530
rect 11678 10490 11698 10530
rect 11618 10430 11698 10490
rect 11618 10390 11638 10430
rect 11678 10390 11698 10430
rect 11618 10330 11698 10390
rect 11618 10290 11638 10330
rect 11678 10290 11698 10330
rect 11618 10230 11698 10290
rect 11618 10190 11638 10230
rect 11678 10190 11698 10230
rect 11618 10130 11698 10190
rect 11618 10090 11638 10130
rect 11678 10090 11698 10130
rect 11618 10060 11698 10090
rect 11798 10630 11878 10660
rect 11798 10590 11818 10630
rect 11858 10590 11878 10630
rect 11798 10530 11878 10590
rect 11798 10490 11818 10530
rect 11858 10490 11878 10530
rect 11798 10430 11878 10490
rect 11798 10390 11818 10430
rect 11858 10390 11878 10430
rect 11798 10330 11878 10390
rect 11798 10290 11818 10330
rect 11858 10290 11878 10330
rect 11798 10230 11878 10290
rect 11798 10190 11818 10230
rect 11858 10190 11878 10230
rect 11798 10130 11878 10190
rect 11798 10090 11818 10130
rect 11858 10090 11878 10130
rect 11798 10060 11878 10090
rect 11978 10630 12058 10660
rect 11978 10590 11998 10630
rect 12038 10590 12058 10630
rect 11978 10530 12058 10590
rect 11978 10490 11998 10530
rect 12038 10490 12058 10530
rect 11978 10430 12058 10490
rect 11978 10390 11998 10430
rect 12038 10390 12058 10430
rect 11978 10330 12058 10390
rect 11978 10290 11998 10330
rect 12038 10290 12058 10330
rect 11978 10230 12058 10290
rect 11978 10190 11998 10230
rect 12038 10190 12058 10230
rect 11978 10130 12058 10190
rect 11978 10090 11998 10130
rect 12038 10090 12058 10130
rect 11978 10060 12058 10090
rect 12158 10630 12238 10660
rect 12158 10590 12178 10630
rect 12218 10590 12238 10630
rect 12158 10530 12238 10590
rect 12158 10490 12178 10530
rect 12218 10490 12238 10530
rect 12158 10430 12238 10490
rect 12158 10390 12178 10430
rect 12218 10390 12238 10430
rect 12158 10330 12238 10390
rect 12158 10290 12178 10330
rect 12218 10290 12238 10330
rect 12158 10230 12238 10290
rect 12158 10190 12178 10230
rect 12218 10190 12238 10230
rect 12158 10130 12238 10190
rect 12158 10090 12178 10130
rect 12218 10090 12238 10130
rect 12158 10060 12238 10090
rect 12338 10630 12418 10660
rect 12338 10590 12358 10630
rect 12398 10590 12418 10630
rect 12338 10530 12418 10590
rect 12338 10490 12358 10530
rect 12398 10490 12418 10530
rect 12338 10430 12418 10490
rect 12338 10390 12358 10430
rect 12398 10390 12418 10430
rect 12338 10330 12418 10390
rect 12338 10290 12358 10330
rect 12398 10290 12418 10330
rect 12338 10230 12418 10290
rect 12338 10190 12358 10230
rect 12398 10190 12418 10230
rect 12338 10130 12418 10190
rect 12338 10090 12358 10130
rect 12398 10090 12418 10130
rect 12338 10060 12418 10090
rect 12518 10630 12598 10660
rect 12518 10590 12538 10630
rect 12578 10590 12598 10630
rect 12518 10530 12598 10590
rect 12518 10490 12538 10530
rect 12578 10490 12598 10530
rect 12518 10430 12598 10490
rect 12518 10390 12538 10430
rect 12578 10390 12598 10430
rect 12518 10330 12598 10390
rect 12518 10290 12538 10330
rect 12578 10290 12598 10330
rect 12518 10230 12598 10290
rect 12518 10190 12538 10230
rect 12578 10190 12598 10230
rect 12518 10130 12598 10190
rect 12518 10090 12538 10130
rect 12578 10090 12598 10130
rect 12518 10060 12598 10090
rect 12698 10630 12778 10660
rect 12698 10590 12718 10630
rect 12758 10590 12778 10630
rect 12698 10530 12778 10590
rect 12698 10490 12718 10530
rect 12758 10490 12778 10530
rect 12698 10430 12778 10490
rect 12698 10390 12718 10430
rect 12758 10390 12778 10430
rect 12698 10330 12778 10390
rect 12698 10290 12718 10330
rect 12758 10290 12778 10330
rect 12698 10230 12778 10290
rect 12698 10190 12718 10230
rect 12758 10190 12778 10230
rect 12698 10130 12778 10190
rect 12698 10090 12718 10130
rect 12758 10090 12778 10130
rect 12698 10060 12778 10090
rect 12878 10630 12958 10660
rect 12878 10590 12898 10630
rect 12938 10590 12958 10630
rect 12878 10530 12958 10590
rect 12878 10490 12898 10530
rect 12938 10490 12958 10530
rect 12878 10430 12958 10490
rect 12878 10390 12898 10430
rect 12938 10390 12958 10430
rect 12878 10330 12958 10390
rect 12878 10290 12898 10330
rect 12938 10290 12958 10330
rect 12878 10230 12958 10290
rect 12878 10190 12898 10230
rect 12938 10190 12958 10230
rect 12878 10130 12958 10190
rect 12878 10090 12898 10130
rect 12938 10090 12958 10130
rect 12878 10060 12958 10090
rect 13058 10630 13138 10660
rect 13058 10590 13078 10630
rect 13118 10590 13138 10630
rect 13058 10530 13138 10590
rect 13058 10490 13078 10530
rect 13118 10490 13138 10530
rect 13058 10430 13138 10490
rect 13058 10390 13078 10430
rect 13118 10390 13138 10430
rect 13058 10330 13138 10390
rect 13058 10290 13078 10330
rect 13118 10290 13138 10330
rect 13058 10230 13138 10290
rect 13058 10190 13078 10230
rect 13118 10190 13138 10230
rect 13058 10130 13138 10190
rect 13058 10090 13078 10130
rect 13118 10090 13138 10130
rect 13058 10060 13138 10090
rect 13238 10630 13318 10660
rect 13238 10590 13258 10630
rect 13298 10590 13318 10630
rect 13238 10530 13318 10590
rect 13238 10490 13258 10530
rect 13298 10490 13318 10530
rect 13238 10430 13318 10490
rect 13238 10390 13258 10430
rect 13298 10390 13318 10430
rect 13238 10330 13318 10390
rect 13238 10290 13258 10330
rect 13298 10290 13318 10330
rect 13238 10230 13318 10290
rect 13238 10190 13258 10230
rect 13298 10190 13318 10230
rect 13238 10130 13318 10190
rect 13238 10090 13258 10130
rect 13298 10090 13318 10130
rect 13238 10060 13318 10090
rect 13418 10630 13498 10660
rect 13418 10590 13438 10630
rect 13478 10590 13498 10630
rect 13418 10530 13498 10590
rect 13418 10490 13438 10530
rect 13478 10490 13498 10530
rect 13418 10430 13498 10490
rect 13418 10390 13438 10430
rect 13478 10390 13498 10430
rect 13418 10330 13498 10390
rect 13418 10290 13438 10330
rect 13478 10290 13498 10330
rect 13418 10230 13498 10290
rect 13418 10190 13438 10230
rect 13478 10190 13498 10230
rect 13418 10130 13498 10190
rect 13418 10090 13438 10130
rect 13478 10090 13498 10130
rect 13418 10060 13498 10090
rect 13598 10630 13678 10660
rect 13598 10590 13618 10630
rect 13658 10590 13678 10630
rect 13598 10530 13678 10590
rect 13598 10490 13618 10530
rect 13658 10490 13678 10530
rect 13598 10430 13678 10490
rect 13598 10390 13618 10430
rect 13658 10390 13678 10430
rect 13598 10330 13678 10390
rect 13598 10290 13618 10330
rect 13658 10290 13678 10330
rect 13598 10230 13678 10290
rect 13598 10190 13618 10230
rect 13658 10190 13678 10230
rect 13598 10130 13678 10190
rect 13598 10090 13618 10130
rect 13658 10090 13678 10130
rect 13598 10060 13678 10090
rect 13778 10630 13858 10660
rect 13778 10590 13798 10630
rect 13838 10590 13858 10630
rect 13778 10530 13858 10590
rect 13778 10490 13798 10530
rect 13838 10490 13858 10530
rect 13778 10430 13858 10490
rect 13778 10390 13798 10430
rect 13838 10390 13858 10430
rect 13778 10330 13858 10390
rect 13778 10290 13798 10330
rect 13838 10290 13858 10330
rect 13778 10230 13858 10290
rect 13778 10190 13798 10230
rect 13838 10190 13858 10230
rect 13778 10130 13858 10190
rect 13778 10090 13798 10130
rect 13838 10090 13858 10130
rect 13778 10060 13858 10090
rect 13958 10630 14038 10660
rect 13958 10590 13978 10630
rect 14018 10590 14038 10630
rect 13958 10530 14038 10590
rect 13958 10490 13978 10530
rect 14018 10490 14038 10530
rect 13958 10430 14038 10490
rect 13958 10390 13978 10430
rect 14018 10390 14038 10430
rect 13958 10330 14038 10390
rect 13958 10290 13978 10330
rect 14018 10290 14038 10330
rect 13958 10230 14038 10290
rect 13958 10190 13978 10230
rect 14018 10190 14038 10230
rect 13958 10130 14038 10190
rect 13958 10090 13978 10130
rect 14018 10090 14038 10130
rect 13958 10060 14038 10090
rect 14138 10630 14218 10660
rect 14138 10590 14158 10630
rect 14198 10590 14218 10630
rect 14138 10530 14218 10590
rect 14138 10490 14158 10530
rect 14198 10490 14218 10530
rect 14138 10430 14218 10490
rect 14138 10390 14158 10430
rect 14198 10390 14218 10430
rect 14138 10330 14218 10390
rect 14138 10290 14158 10330
rect 14198 10290 14218 10330
rect 14138 10230 14218 10290
rect 14138 10190 14158 10230
rect 14198 10190 14218 10230
rect 14138 10130 14218 10190
rect 14138 10090 14158 10130
rect 14198 10090 14218 10130
rect 14138 10060 14218 10090
rect 14318 10630 14398 10660
rect 14318 10590 14338 10630
rect 14378 10590 14398 10630
rect 14318 10530 14398 10590
rect 14318 10490 14338 10530
rect 14378 10490 14398 10530
rect 14318 10430 14398 10490
rect 14318 10390 14338 10430
rect 14378 10390 14398 10430
rect 14318 10330 14398 10390
rect 14318 10290 14338 10330
rect 14378 10290 14398 10330
rect 14318 10230 14398 10290
rect 14318 10190 14338 10230
rect 14378 10190 14398 10230
rect 14318 10130 14398 10190
rect 14318 10090 14338 10130
rect 14378 10090 14398 10130
rect 14318 10060 14398 10090
rect 14498 10630 14578 10660
rect 14498 10590 14518 10630
rect 14558 10590 14578 10630
rect 14498 10530 14578 10590
rect 14498 10490 14518 10530
rect 14558 10490 14578 10530
rect 14498 10430 14578 10490
rect 14498 10390 14518 10430
rect 14558 10390 14578 10430
rect 14498 10330 14578 10390
rect 14498 10290 14518 10330
rect 14558 10290 14578 10330
rect 14498 10230 14578 10290
rect 14498 10190 14518 10230
rect 14558 10190 14578 10230
rect 14498 10130 14578 10190
rect 14498 10090 14518 10130
rect 14558 10090 14578 10130
rect 14498 10060 14578 10090
rect 14678 10630 14758 10660
rect 14678 10590 14698 10630
rect 14738 10590 14758 10630
rect 14678 10530 14758 10590
rect 14678 10490 14698 10530
rect 14738 10490 14758 10530
rect 14678 10430 14758 10490
rect 14678 10390 14698 10430
rect 14738 10390 14758 10430
rect 14678 10330 14758 10390
rect 14678 10290 14698 10330
rect 14738 10290 14758 10330
rect 14678 10230 14758 10290
rect 14678 10190 14698 10230
rect 14738 10190 14758 10230
rect 14678 10130 14758 10190
rect 14678 10090 14698 10130
rect 14738 10090 14758 10130
rect 14678 10060 14758 10090
rect 14858 10630 14938 10660
rect 14858 10590 14878 10630
rect 14918 10590 14938 10630
rect 14858 10530 14938 10590
rect 14858 10490 14878 10530
rect 14918 10490 14938 10530
rect 14858 10430 14938 10490
rect 14858 10390 14878 10430
rect 14918 10390 14938 10430
rect 14858 10330 14938 10390
rect 14858 10290 14878 10330
rect 14918 10290 14938 10330
rect 14858 10230 14938 10290
rect 15478 10430 15568 10460
rect 15478 10390 15508 10430
rect 15548 10390 15568 10430
rect 15478 10330 15568 10390
rect 15478 10290 15508 10330
rect 15548 10290 15568 10330
rect 15478 10260 15568 10290
rect 15598 10430 15678 10460
rect 15598 10390 15618 10430
rect 15658 10390 15678 10430
rect 15598 10330 15678 10390
rect 15598 10290 15618 10330
rect 15658 10290 15678 10330
rect 15598 10260 15678 10290
rect 15708 10430 15788 10460
rect 15708 10390 15728 10430
rect 15768 10390 15788 10430
rect 15708 10330 15788 10390
rect 15708 10290 15728 10330
rect 15768 10290 15788 10330
rect 15708 10260 15788 10290
rect 15818 10430 15898 10460
rect 15818 10390 15838 10430
rect 15878 10390 15898 10430
rect 15818 10330 15898 10390
rect 15818 10290 15838 10330
rect 15878 10290 15898 10330
rect 15818 10260 15898 10290
rect 15928 10430 16008 10460
rect 15928 10390 15948 10430
rect 15988 10390 16008 10430
rect 15928 10330 16008 10390
rect 15928 10290 15948 10330
rect 15988 10290 16008 10330
rect 15928 10260 16008 10290
rect 14858 10190 14878 10230
rect 14918 10190 14938 10230
rect 14858 10130 14938 10190
rect 14858 10090 14878 10130
rect 14918 10090 14938 10130
rect 14858 10060 14938 10090
rect 11628 9630 11708 9660
rect 11628 9590 11648 9630
rect 11688 9590 11708 9630
rect 11628 9530 11708 9590
rect 11628 9490 11648 9530
rect 11688 9490 11708 9530
rect 11628 9460 11708 9490
rect 11738 9630 11818 9660
rect 11738 9590 11758 9630
rect 11798 9590 11818 9630
rect 11738 9530 11818 9590
rect 11738 9490 11758 9530
rect 11798 9490 11818 9530
rect 11738 9460 11818 9490
rect 11848 9630 11928 9660
rect 11848 9590 11868 9630
rect 11908 9590 11928 9630
rect 11848 9530 11928 9590
rect 11848 9490 11868 9530
rect 11908 9490 11928 9530
rect 11848 9460 11928 9490
rect 11958 9630 12038 9660
rect 11958 9590 11978 9630
rect 12018 9590 12038 9630
rect 11958 9530 12038 9590
rect 11958 9490 11978 9530
rect 12018 9490 12038 9530
rect 11958 9460 12038 9490
rect 12068 9630 12148 9660
rect 12068 9590 12088 9630
rect 12128 9590 12148 9630
rect 12068 9530 12148 9590
rect 12068 9490 12088 9530
rect 12128 9490 12148 9530
rect 12068 9460 12148 9490
rect 12178 9630 12258 9660
rect 12178 9590 12198 9630
rect 12238 9590 12258 9630
rect 12178 9530 12258 9590
rect 12178 9490 12198 9530
rect 12238 9490 12258 9530
rect 12178 9460 12258 9490
rect 12288 9630 12368 9660
rect 12288 9590 12308 9630
rect 12348 9590 12368 9630
rect 12288 9530 12368 9590
rect 12288 9490 12308 9530
rect 12348 9490 12368 9530
rect 12288 9460 12368 9490
rect 12398 9630 12478 9660
rect 12398 9590 12418 9630
rect 12458 9590 12478 9630
rect 12398 9530 12478 9590
rect 12398 9490 12418 9530
rect 12458 9490 12478 9530
rect 12398 9460 12478 9490
rect 12508 9630 12588 9660
rect 12508 9590 12528 9630
rect 12568 9590 12588 9630
rect 12508 9530 12588 9590
rect 12508 9490 12528 9530
rect 12568 9490 12588 9530
rect 12508 9460 12588 9490
rect 12618 9630 12698 9660
rect 12618 9590 12638 9630
rect 12678 9590 12698 9630
rect 12618 9530 12698 9590
rect 12618 9490 12638 9530
rect 12678 9490 12698 9530
rect 12618 9460 12698 9490
rect 12728 9630 12808 9660
rect 12728 9590 12748 9630
rect 12788 9590 12808 9630
rect 12728 9530 12808 9590
rect 12728 9490 12748 9530
rect 12788 9490 12808 9530
rect 12728 9460 12808 9490
rect 12838 9630 12918 9660
rect 12838 9590 12858 9630
rect 12898 9590 12918 9630
rect 12838 9530 12918 9590
rect 12838 9490 12858 9530
rect 12898 9490 12918 9530
rect 12838 9460 12918 9490
rect 12948 9630 13028 9660
rect 12948 9590 12968 9630
rect 13008 9590 13028 9630
rect 12948 9530 13028 9590
rect 12948 9490 12968 9530
rect 13008 9490 13028 9530
rect 12948 9460 13028 9490
rect 13528 9630 13608 9660
rect 13528 9590 13548 9630
rect 13588 9590 13608 9630
rect 13528 9530 13608 9590
rect 13528 9490 13548 9530
rect 13588 9490 13608 9530
rect 13528 9460 13608 9490
rect 13638 9630 13718 9660
rect 13638 9590 13658 9630
rect 13698 9590 13718 9630
rect 13638 9530 13718 9590
rect 13638 9490 13658 9530
rect 13698 9490 13718 9530
rect 13638 9460 13718 9490
rect 13748 9630 13828 9660
rect 13748 9590 13768 9630
rect 13808 9590 13828 9630
rect 13748 9530 13828 9590
rect 13748 9490 13768 9530
rect 13808 9490 13828 9530
rect 13748 9460 13828 9490
rect 13858 9630 13938 9660
rect 13858 9590 13878 9630
rect 13918 9590 13938 9630
rect 13858 9530 13938 9590
rect 13858 9490 13878 9530
rect 13918 9490 13938 9530
rect 13858 9460 13938 9490
rect 13968 9630 14048 9660
rect 13968 9590 13988 9630
rect 14028 9590 14048 9630
rect 13968 9530 14048 9590
rect 13968 9490 13988 9530
rect 14028 9490 14048 9530
rect 13968 9460 14048 9490
rect 14078 9630 14158 9660
rect 14078 9590 14098 9630
rect 14138 9590 14158 9630
rect 14078 9530 14158 9590
rect 14078 9490 14098 9530
rect 14138 9490 14158 9530
rect 14078 9460 14158 9490
rect 14188 9630 14268 9660
rect 14188 9590 14208 9630
rect 14248 9590 14268 9630
rect 14188 9530 14268 9590
rect 14188 9490 14208 9530
rect 14248 9490 14268 9530
rect 14188 9460 14268 9490
rect 14298 9630 14378 9660
rect 14298 9590 14318 9630
rect 14358 9590 14378 9630
rect 14298 9530 14378 9590
rect 14298 9490 14318 9530
rect 14358 9490 14378 9530
rect 14298 9460 14378 9490
rect 14408 9630 14488 9660
rect 14408 9590 14428 9630
rect 14468 9590 14488 9630
rect 14408 9530 14488 9590
rect 14408 9490 14428 9530
rect 14468 9490 14488 9530
rect 14408 9460 14488 9490
rect 14518 9630 14598 9660
rect 14518 9590 14538 9630
rect 14578 9590 14598 9630
rect 14518 9530 14598 9590
rect 14518 9490 14538 9530
rect 14578 9490 14598 9530
rect 14518 9460 14598 9490
rect 14628 9630 14708 9660
rect 14628 9590 14648 9630
rect 14688 9590 14708 9630
rect 14628 9530 14708 9590
rect 14628 9490 14648 9530
rect 14688 9490 14708 9530
rect 14628 9460 14708 9490
rect 14738 9630 14818 9660
rect 14738 9590 14758 9630
rect 14798 9590 14818 9630
rect 14738 9530 14818 9590
rect 14738 9490 14758 9530
rect 14798 9490 14818 9530
rect 14738 9460 14818 9490
rect 14848 9630 14928 9660
rect 14848 9590 14868 9630
rect 14908 9590 14928 9630
rect 14848 9530 14928 9590
rect 14848 9490 14868 9530
rect 14908 9490 14928 9530
rect 14848 9460 14928 9490
rect 13248 7640 13328 7670
rect 13248 7600 13268 7640
rect 13308 7600 13328 7640
rect 13248 7540 13328 7600
rect 13248 7500 13268 7540
rect 13308 7500 13328 7540
rect 13248 7440 13328 7500
rect 13248 7400 13268 7440
rect 13308 7400 13328 7440
rect 13248 7340 13328 7400
rect 13248 7300 13268 7340
rect 13308 7300 13328 7340
rect 13248 7270 13328 7300
rect 13358 7640 13438 7670
rect 13358 7600 13378 7640
rect 13418 7600 13438 7640
rect 13358 7540 13438 7600
rect 13358 7500 13378 7540
rect 13418 7500 13438 7540
rect 13358 7440 13438 7500
rect 13358 7400 13378 7440
rect 13418 7400 13438 7440
rect 13358 7340 13438 7400
rect 13358 7300 13378 7340
rect 13418 7300 13438 7340
rect 13358 7270 13438 7300
rect 13468 7640 13548 7670
rect 13468 7600 13488 7640
rect 13528 7600 13548 7640
rect 13468 7540 13548 7600
rect 13468 7500 13488 7540
rect 13528 7500 13548 7540
rect 13468 7440 13548 7500
rect 13468 7400 13488 7440
rect 13528 7400 13548 7440
rect 13468 7340 13548 7400
rect 13468 7300 13488 7340
rect 13528 7300 13548 7340
rect 13468 7270 13548 7300
rect 13768 7640 13848 7670
rect 13768 7600 13788 7640
rect 13828 7600 13848 7640
rect 13768 7540 13848 7600
rect 13768 7500 13788 7540
rect 13828 7500 13848 7540
rect 13768 7440 13848 7500
rect 13768 7400 13788 7440
rect 13828 7400 13848 7440
rect 13768 7340 13848 7400
rect 13768 7300 13788 7340
rect 13828 7300 13848 7340
rect 13768 7270 13848 7300
rect 13878 7640 13958 7670
rect 13878 7600 13898 7640
rect 13938 7600 13958 7640
rect 13878 7540 13958 7600
rect 13878 7500 13898 7540
rect 13938 7500 13958 7540
rect 13878 7440 13958 7500
rect 13878 7400 13898 7440
rect 13938 7400 13958 7440
rect 13878 7340 13958 7400
rect 13878 7300 13898 7340
rect 13938 7300 13958 7340
rect 13878 7270 13958 7300
rect 13988 7640 14068 7670
rect 14148 7640 14228 7670
rect 13988 7600 14008 7640
rect 14048 7600 14068 7640
rect 14148 7600 14168 7640
rect 14208 7600 14228 7640
rect 13988 7540 14068 7600
rect 14148 7540 14228 7600
rect 13988 7500 14008 7540
rect 14048 7500 14068 7540
rect 14148 7500 14168 7540
rect 14208 7500 14228 7540
rect 13988 7440 14068 7500
rect 14148 7440 14228 7500
rect 13988 7400 14008 7440
rect 14048 7400 14068 7440
rect 14148 7400 14168 7440
rect 14208 7400 14228 7440
rect 13988 7340 14068 7400
rect 14148 7340 14228 7400
rect 13988 7300 14008 7340
rect 14048 7300 14068 7340
rect 14148 7300 14168 7340
rect 14208 7300 14228 7340
rect 13988 7270 14068 7300
rect 14148 7270 14228 7300
rect 14258 7640 14338 7670
rect 14258 7600 14278 7640
rect 14318 7600 14338 7640
rect 14258 7540 14338 7600
rect 14258 7500 14278 7540
rect 14318 7500 14338 7540
rect 14258 7440 14338 7500
rect 14258 7400 14278 7440
rect 14318 7400 14338 7440
rect 14258 7340 14338 7400
rect 14258 7300 14278 7340
rect 14318 7300 14338 7340
rect 14258 7270 14338 7300
rect 14368 7640 14448 7670
rect 14368 7600 14388 7640
rect 14428 7600 14448 7640
rect 14368 7540 14448 7600
rect 14368 7500 14388 7540
rect 14428 7500 14448 7540
rect 14368 7440 14448 7500
rect 14368 7400 14388 7440
rect 14428 7400 14448 7440
rect 14368 7340 14448 7400
rect 14368 7300 14388 7340
rect 14428 7300 14448 7340
rect 14368 7270 14448 7300
rect 14668 7640 14748 7670
rect 14668 7600 14688 7640
rect 14728 7600 14748 7640
rect 14668 7540 14748 7600
rect 14668 7500 14688 7540
rect 14728 7500 14748 7540
rect 14668 7440 14748 7500
rect 14668 7400 14688 7440
rect 14728 7400 14748 7440
rect 14668 7340 14748 7400
rect 14668 7300 14688 7340
rect 14728 7300 14748 7340
rect 14668 7270 14748 7300
rect 14778 7640 14858 7670
rect 14778 7600 14798 7640
rect 14838 7600 14858 7640
rect 14778 7540 14858 7600
rect 14778 7500 14798 7540
rect 14838 7500 14858 7540
rect 14778 7440 14858 7500
rect 14778 7400 14798 7440
rect 14838 7400 14858 7440
rect 14778 7340 14858 7400
rect 14778 7300 14798 7340
rect 14838 7300 14858 7340
rect 14778 7270 14858 7300
rect 14888 7640 14968 7670
rect 14888 7600 14908 7640
rect 14948 7600 14968 7640
rect 14888 7540 14968 7600
rect 14888 7500 14908 7540
rect 14948 7500 14968 7540
rect 14888 7440 14968 7500
rect 14888 7400 14908 7440
rect 14948 7400 14968 7440
rect 14888 7340 14968 7400
rect 14888 7300 14908 7340
rect 14948 7300 14968 7340
rect 14888 7270 14968 7300
rect 15178 7640 15258 7670
rect 15178 7600 15198 7640
rect 15238 7600 15258 7640
rect 15178 7540 15258 7600
rect 15178 7500 15198 7540
rect 15238 7500 15258 7540
rect 15178 7440 15258 7500
rect 15178 7400 15198 7440
rect 15238 7400 15258 7440
rect 15178 7340 15258 7400
rect 15178 7300 15198 7340
rect 15238 7300 15258 7340
rect 15178 7270 15258 7300
rect 15288 7640 15368 7670
rect 15288 7600 15308 7640
rect 15348 7600 15368 7640
rect 15288 7540 15368 7600
rect 15288 7500 15308 7540
rect 15348 7500 15368 7540
rect 15288 7440 15368 7500
rect 15288 7400 15308 7440
rect 15348 7400 15368 7440
rect 15288 7340 15368 7400
rect 15288 7300 15308 7340
rect 15348 7300 15368 7340
rect 15288 7270 15368 7300
rect 15508 7640 15588 7670
rect 15508 7600 15528 7640
rect 15568 7600 15588 7640
rect 15508 7540 15588 7600
rect 15508 7500 15528 7540
rect 15568 7500 15588 7540
rect 15508 7440 15588 7500
rect 15508 7400 15528 7440
rect 15568 7400 15588 7440
rect 15508 7340 15588 7400
rect 15508 7300 15528 7340
rect 15568 7300 15588 7340
rect 15508 7270 15588 7300
rect 15618 7640 15698 7670
rect 15618 7600 15638 7640
rect 15678 7600 15698 7640
rect 15618 7540 15698 7600
rect 15618 7500 15638 7540
rect 15678 7500 15698 7540
rect 15618 7440 15698 7500
rect 15618 7400 15638 7440
rect 15678 7400 15698 7440
rect 15618 7340 15698 7400
rect 15618 7300 15638 7340
rect 15678 7300 15698 7340
rect 15618 7270 15698 7300
rect 15838 7640 15918 7670
rect 15838 7600 15858 7640
rect 15898 7600 15918 7640
rect 15838 7540 15918 7600
rect 15838 7500 15858 7540
rect 15898 7500 15918 7540
rect 15838 7440 15918 7500
rect 15838 7400 15858 7440
rect 15898 7400 15918 7440
rect 15838 7340 15918 7400
rect 15838 7300 15858 7340
rect 15898 7300 15918 7340
rect 15838 7270 15918 7300
rect 15948 7640 16028 7670
rect 15948 7600 15968 7640
rect 16008 7600 16028 7640
rect 15948 7540 16028 7600
rect 15948 7500 15968 7540
rect 16008 7500 16028 7540
rect 15948 7440 16028 7500
rect 15948 7400 15968 7440
rect 16008 7400 16028 7440
rect 15948 7340 16028 7400
rect 15948 7300 15968 7340
rect 16008 7300 16028 7340
rect 15948 7270 16028 7300
rect 16378 7640 16478 7670
rect 16378 7600 16408 7640
rect 16448 7600 16478 7640
rect 16378 7540 16478 7600
rect 16378 7500 16408 7540
rect 16448 7500 16478 7540
rect 16378 7440 16478 7500
rect 16378 7400 16408 7440
rect 16448 7400 16478 7440
rect 16378 7340 16478 7400
rect 16378 7300 16408 7340
rect 16448 7300 16478 7340
rect 16378 7270 16478 7300
rect 16508 7640 16608 7670
rect 16508 7600 16538 7640
rect 16578 7600 16608 7640
rect 16508 7540 16608 7600
rect 16508 7500 16538 7540
rect 16578 7500 16608 7540
rect 16508 7440 16608 7500
rect 16508 7400 16538 7440
rect 16578 7400 16608 7440
rect 16508 7340 16608 7400
rect 16508 7300 16538 7340
rect 16578 7300 16608 7340
rect 16508 7270 16608 7300
rect 16768 7640 16868 7670
rect 16768 7600 16798 7640
rect 16838 7600 16868 7640
rect 16768 7540 16868 7600
rect 16768 7500 16798 7540
rect 16838 7500 16868 7540
rect 16768 7440 16868 7500
rect 16768 7400 16798 7440
rect 16838 7400 16868 7440
rect 16768 7340 16868 7400
rect 16768 7300 16798 7340
rect 16838 7300 16868 7340
rect 16768 7270 16868 7300
rect 16898 7640 16998 7670
rect 16898 7600 16928 7640
rect 16968 7600 16998 7640
rect 16898 7540 16998 7600
rect 16898 7500 16928 7540
rect 16968 7500 16998 7540
rect 16898 7440 16998 7500
rect 16898 7400 16928 7440
rect 16968 7400 16998 7440
rect 16898 7340 16998 7400
rect 16898 7300 16928 7340
rect 16968 7300 16998 7340
rect 16898 7270 16998 7300
rect 17158 7640 17258 7670
rect 17158 7600 17188 7640
rect 17228 7600 17258 7640
rect 17158 7540 17258 7600
rect 17158 7500 17188 7540
rect 17228 7500 17258 7540
rect 17158 7440 17258 7500
rect 17158 7400 17188 7440
rect 17228 7400 17258 7440
rect 17158 7340 17258 7400
rect 17158 7300 17188 7340
rect 17228 7300 17258 7340
rect 17158 7270 17258 7300
rect 17288 7640 17388 7670
rect 17288 7600 17318 7640
rect 17358 7600 17388 7640
rect 17288 7540 17388 7600
rect 17288 7500 17318 7540
rect 17358 7500 17388 7540
rect 17288 7440 17388 7500
rect 17288 7400 17318 7440
rect 17358 7400 17388 7440
rect 17288 7340 17388 7400
rect 17288 7300 17318 7340
rect 17358 7300 17388 7340
rect 17288 7270 17388 7300
rect 17448 7640 17548 7670
rect 17448 7600 17478 7640
rect 17518 7600 17548 7640
rect 17448 7540 17548 7600
rect 17448 7500 17478 7540
rect 17518 7500 17548 7540
rect 17448 7440 17548 7500
rect 17448 7400 17478 7440
rect 17518 7400 17548 7440
rect 17448 7340 17548 7400
rect 17448 7300 17478 7340
rect 17518 7300 17548 7340
rect 17448 7270 17548 7300
rect 17578 7640 17678 7670
rect 17578 7600 17608 7640
rect 17648 7600 17678 7640
rect 17578 7540 17678 7600
rect 17578 7500 17608 7540
rect 17648 7500 17678 7540
rect 17578 7440 17678 7500
rect 17578 7400 17608 7440
rect 17648 7400 17678 7440
rect 17578 7340 17678 7400
rect 17578 7300 17608 7340
rect 17648 7300 17678 7340
rect 17578 7270 17678 7300
rect 19528 6910 19628 6940
rect 13248 6880 13328 6910
rect 13248 6840 13268 6880
rect 13308 6840 13328 6880
rect 13248 6780 13328 6840
rect 13248 6740 13268 6780
rect 13308 6740 13328 6780
rect 13248 6680 13328 6740
rect 13248 6640 13268 6680
rect 13308 6640 13328 6680
rect 13248 6580 13328 6640
rect 13248 6540 13268 6580
rect 13308 6540 13328 6580
rect 13248 6510 13328 6540
rect 13358 6880 13438 6910
rect 13358 6840 13378 6880
rect 13418 6840 13438 6880
rect 13358 6780 13438 6840
rect 13358 6740 13378 6780
rect 13418 6740 13438 6780
rect 13358 6680 13438 6740
rect 13358 6640 13378 6680
rect 13418 6640 13438 6680
rect 13358 6580 13438 6640
rect 13358 6540 13378 6580
rect 13418 6540 13438 6580
rect 13358 6510 13438 6540
rect 13468 6880 13548 6910
rect 13468 6840 13488 6880
rect 13528 6840 13548 6880
rect 13468 6780 13548 6840
rect 13468 6740 13488 6780
rect 13528 6740 13548 6780
rect 13468 6680 13548 6740
rect 13468 6640 13488 6680
rect 13528 6640 13548 6680
rect 13468 6580 13548 6640
rect 13468 6540 13488 6580
rect 13528 6540 13548 6580
rect 13468 6510 13548 6540
rect 13768 6880 13848 6910
rect 13768 6840 13788 6880
rect 13828 6840 13848 6880
rect 13768 6780 13848 6840
rect 13768 6740 13788 6780
rect 13828 6740 13848 6780
rect 13768 6680 13848 6740
rect 13768 6640 13788 6680
rect 13828 6640 13848 6680
rect 13768 6580 13848 6640
rect 13768 6540 13788 6580
rect 13828 6540 13848 6580
rect 13768 6510 13848 6540
rect 13878 6880 13958 6910
rect 13878 6840 13898 6880
rect 13938 6840 13958 6880
rect 13878 6780 13958 6840
rect 13878 6740 13898 6780
rect 13938 6740 13958 6780
rect 13878 6680 13958 6740
rect 13878 6640 13898 6680
rect 13938 6640 13958 6680
rect 13878 6580 13958 6640
rect 13878 6540 13898 6580
rect 13938 6540 13958 6580
rect 13878 6510 13958 6540
rect 13988 6880 14068 6910
rect 14148 6880 14228 6910
rect 13988 6840 14008 6880
rect 14048 6840 14068 6880
rect 14148 6840 14168 6880
rect 14208 6840 14228 6880
rect 13988 6780 14068 6840
rect 14148 6780 14228 6840
rect 13988 6740 14008 6780
rect 14048 6740 14068 6780
rect 14148 6740 14168 6780
rect 14208 6740 14228 6780
rect 13988 6680 14068 6740
rect 14148 6680 14228 6740
rect 13988 6640 14008 6680
rect 14048 6640 14068 6680
rect 14148 6640 14168 6680
rect 14208 6640 14228 6680
rect 13988 6580 14068 6640
rect 14148 6580 14228 6640
rect 13988 6540 14008 6580
rect 14048 6540 14068 6580
rect 14148 6540 14168 6580
rect 14208 6540 14228 6580
rect 13988 6510 14068 6540
rect 14148 6510 14228 6540
rect 14258 6880 14338 6910
rect 14258 6840 14278 6880
rect 14318 6840 14338 6880
rect 14258 6780 14338 6840
rect 14258 6740 14278 6780
rect 14318 6740 14338 6780
rect 14258 6680 14338 6740
rect 14258 6640 14278 6680
rect 14318 6640 14338 6680
rect 14258 6580 14338 6640
rect 14258 6540 14278 6580
rect 14318 6540 14338 6580
rect 14258 6510 14338 6540
rect 14368 6880 14448 6910
rect 14368 6840 14388 6880
rect 14428 6840 14448 6880
rect 14368 6780 14448 6840
rect 14368 6740 14388 6780
rect 14428 6740 14448 6780
rect 14368 6680 14448 6740
rect 14368 6640 14388 6680
rect 14428 6640 14448 6680
rect 14368 6580 14448 6640
rect 14368 6540 14388 6580
rect 14428 6540 14448 6580
rect 14368 6510 14448 6540
rect 14668 6880 14748 6910
rect 14668 6840 14688 6880
rect 14728 6840 14748 6880
rect 14668 6780 14748 6840
rect 14668 6740 14688 6780
rect 14728 6740 14748 6780
rect 14668 6680 14748 6740
rect 14668 6640 14688 6680
rect 14728 6640 14748 6680
rect 14668 6580 14748 6640
rect 14668 6540 14688 6580
rect 14728 6540 14748 6580
rect 14668 6510 14748 6540
rect 14778 6880 14858 6910
rect 14778 6840 14798 6880
rect 14838 6840 14858 6880
rect 14778 6780 14858 6840
rect 14778 6740 14798 6780
rect 14838 6740 14858 6780
rect 14778 6680 14858 6740
rect 14778 6640 14798 6680
rect 14838 6640 14858 6680
rect 14778 6580 14858 6640
rect 14778 6540 14798 6580
rect 14838 6540 14858 6580
rect 14778 6510 14858 6540
rect 14888 6880 14968 6910
rect 14888 6840 14908 6880
rect 14948 6840 14968 6880
rect 14888 6780 14968 6840
rect 14888 6740 14908 6780
rect 14948 6740 14968 6780
rect 14888 6680 14968 6740
rect 14888 6640 14908 6680
rect 14948 6640 14968 6680
rect 14888 6580 14968 6640
rect 14888 6540 14908 6580
rect 14948 6540 14968 6580
rect 14888 6510 14968 6540
rect 15168 6900 15268 6910
rect 15188 6880 15268 6900
rect 15188 6840 15208 6880
rect 15248 6840 15268 6880
rect 15188 6780 15268 6840
rect 15188 6740 15208 6780
rect 15248 6740 15268 6780
rect 15188 6680 15268 6740
rect 15188 6640 15208 6680
rect 15248 6640 15268 6680
rect 15188 6580 15268 6640
rect 15188 6540 15208 6580
rect 15248 6540 15268 6580
rect 15188 6510 15268 6540
rect 15298 6880 15378 6910
rect 15298 6840 15318 6880
rect 15358 6840 15378 6880
rect 15298 6780 15378 6840
rect 15298 6740 15318 6780
rect 15358 6740 15378 6780
rect 15298 6680 15378 6740
rect 15298 6640 15318 6680
rect 15358 6640 15378 6680
rect 15298 6580 15378 6640
rect 15298 6540 15318 6580
rect 15358 6540 15378 6580
rect 15298 6510 15378 6540
rect 15408 6880 15488 6910
rect 15408 6840 15428 6880
rect 15468 6840 15488 6880
rect 15408 6780 15488 6840
rect 15408 6740 15428 6780
rect 15468 6740 15488 6780
rect 15408 6680 15488 6740
rect 15408 6640 15428 6680
rect 15468 6640 15488 6680
rect 15408 6580 15488 6640
rect 15408 6540 15428 6580
rect 15468 6540 15488 6580
rect 15408 6510 15488 6540
rect 15628 6880 15708 6910
rect 15628 6840 15648 6880
rect 15688 6840 15708 6880
rect 15628 6780 15708 6840
rect 15628 6740 15648 6780
rect 15688 6740 15708 6780
rect 15628 6680 15708 6740
rect 15628 6640 15648 6680
rect 15688 6640 15708 6680
rect 15628 6580 15708 6640
rect 15628 6540 15648 6580
rect 15688 6540 15708 6580
rect 15628 6510 15708 6540
rect 15738 6880 15818 6910
rect 15738 6840 15758 6880
rect 15798 6840 15818 6880
rect 15738 6780 15818 6840
rect 15738 6740 15758 6780
rect 15798 6740 15818 6780
rect 15738 6680 15818 6740
rect 15738 6640 15758 6680
rect 15798 6640 15818 6680
rect 15738 6580 15818 6640
rect 15738 6540 15758 6580
rect 15798 6540 15818 6580
rect 15738 6510 15818 6540
rect 15958 6880 16038 6910
rect 15958 6840 15978 6880
rect 16018 6840 16038 6880
rect 15958 6780 16038 6840
rect 15958 6740 15978 6780
rect 16018 6740 16038 6780
rect 15958 6680 16038 6740
rect 15958 6640 15978 6680
rect 16018 6640 16038 6680
rect 15958 6580 16038 6640
rect 15958 6540 15978 6580
rect 16018 6540 16038 6580
rect 15958 6510 16038 6540
rect 16068 6880 16148 6910
rect 16068 6840 16088 6880
rect 16128 6840 16148 6880
rect 16068 6780 16148 6840
rect 16068 6740 16088 6780
rect 16128 6740 16148 6780
rect 16068 6680 16148 6740
rect 16068 6640 16088 6680
rect 16128 6640 16148 6680
rect 16068 6580 16148 6640
rect 16068 6540 16088 6580
rect 16128 6540 16148 6580
rect 16068 6510 16148 6540
rect 16378 6880 16478 6910
rect 16378 6840 16408 6880
rect 16448 6840 16478 6880
rect 16378 6780 16478 6840
rect 16378 6740 16408 6780
rect 16448 6740 16478 6780
rect 16378 6680 16478 6740
rect 16378 6640 16408 6680
rect 16448 6640 16478 6680
rect 16378 6580 16478 6640
rect 16378 6540 16408 6580
rect 16448 6540 16478 6580
rect 16378 6510 16478 6540
rect 16508 6880 16608 6910
rect 16508 6840 16538 6880
rect 16578 6840 16608 6880
rect 16508 6780 16608 6840
rect 16508 6740 16538 6780
rect 16578 6740 16608 6780
rect 16508 6680 16608 6740
rect 16508 6640 16538 6680
rect 16578 6640 16608 6680
rect 16508 6580 16608 6640
rect 16508 6540 16538 6580
rect 16578 6540 16608 6580
rect 16508 6510 16608 6540
rect 16768 6880 16868 6910
rect 16768 6840 16798 6880
rect 16838 6840 16868 6880
rect 16768 6780 16868 6840
rect 16768 6740 16798 6780
rect 16838 6740 16868 6780
rect 16768 6680 16868 6740
rect 16768 6640 16798 6680
rect 16838 6640 16868 6680
rect 16768 6580 16868 6640
rect 16768 6540 16798 6580
rect 16838 6540 16868 6580
rect 16768 6510 16868 6540
rect 16898 6880 16998 6910
rect 16898 6840 16928 6880
rect 16968 6840 16998 6880
rect 16898 6780 16998 6840
rect 16898 6740 16928 6780
rect 16968 6740 16998 6780
rect 16898 6680 16998 6740
rect 16898 6640 16928 6680
rect 16968 6640 16998 6680
rect 16898 6580 16998 6640
rect 16898 6540 16928 6580
rect 16968 6540 16998 6580
rect 16898 6510 16998 6540
rect 17158 6880 17258 6910
rect 17158 6840 17188 6880
rect 17228 6840 17258 6880
rect 17158 6780 17258 6840
rect 17158 6740 17188 6780
rect 17228 6740 17258 6780
rect 17158 6680 17258 6740
rect 17158 6640 17188 6680
rect 17228 6640 17258 6680
rect 17158 6580 17258 6640
rect 17158 6540 17188 6580
rect 17228 6540 17258 6580
rect 17158 6510 17258 6540
rect 17288 6880 17388 6910
rect 17288 6840 17318 6880
rect 17358 6840 17388 6880
rect 17288 6780 17388 6840
rect 17288 6740 17318 6780
rect 17358 6740 17388 6780
rect 17288 6680 17388 6740
rect 17288 6640 17318 6680
rect 17358 6640 17388 6680
rect 17288 6580 17388 6640
rect 17288 6540 17318 6580
rect 17358 6540 17388 6580
rect 17288 6510 17388 6540
rect 17448 6880 17548 6910
rect 17448 6840 17478 6880
rect 17518 6840 17548 6880
rect 17448 6780 17548 6840
rect 17448 6740 17478 6780
rect 17518 6740 17548 6780
rect 17448 6680 17548 6740
rect 17448 6640 17478 6680
rect 17518 6640 17548 6680
rect 17448 6580 17548 6640
rect 17448 6540 17478 6580
rect 17518 6540 17548 6580
rect 17448 6510 17548 6540
rect 17578 6880 17678 6910
rect 17578 6840 17608 6880
rect 17648 6840 17678 6880
rect 17578 6780 17678 6840
rect 17578 6740 17608 6780
rect 17648 6740 17678 6780
rect 17578 6680 17678 6740
rect 17578 6640 17608 6680
rect 17648 6640 17678 6680
rect 17578 6580 17678 6640
rect 17578 6540 17608 6580
rect 17648 6540 17678 6580
rect 17578 6510 17678 6540
rect 17838 6880 17938 6910
rect 17838 6840 17868 6880
rect 17908 6840 17938 6880
rect 17838 6780 17938 6840
rect 17838 6740 17868 6780
rect 17908 6740 17938 6780
rect 17838 6680 17938 6740
rect 17838 6640 17868 6680
rect 17908 6640 17938 6680
rect 17838 6580 17938 6640
rect 17838 6540 17868 6580
rect 17908 6540 17938 6580
rect 17838 6510 17938 6540
rect 17968 6880 18068 6910
rect 17968 6840 17998 6880
rect 18038 6840 18068 6880
rect 17968 6780 18068 6840
rect 17968 6740 17998 6780
rect 18038 6740 18068 6780
rect 17968 6680 18068 6740
rect 17968 6640 17998 6680
rect 18038 6640 18068 6680
rect 17968 6580 18068 6640
rect 17968 6540 17998 6580
rect 18038 6540 18068 6580
rect 19528 6870 19558 6910
rect 19598 6870 19628 6910
rect 19528 6810 19628 6870
rect 19528 6770 19558 6810
rect 19598 6770 19628 6810
rect 19528 6710 19628 6770
rect 19528 6670 19558 6710
rect 19598 6670 19628 6710
rect 19528 6610 19628 6670
rect 19528 6570 19558 6610
rect 19598 6570 19628 6610
rect 19528 6540 19628 6570
rect 19748 6910 19848 6940
rect 19748 6870 19778 6910
rect 19818 6870 19848 6910
rect 19748 6810 19848 6870
rect 19748 6770 19778 6810
rect 19818 6770 19848 6810
rect 19748 6710 19848 6770
rect 19748 6670 19778 6710
rect 19818 6670 19848 6710
rect 19748 6610 19848 6670
rect 19748 6570 19778 6610
rect 19818 6570 19848 6610
rect 19748 6540 19848 6570
rect 19968 6910 20068 6940
rect 19968 6870 19998 6910
rect 20038 6870 20068 6910
rect 19968 6810 20068 6870
rect 19968 6770 19998 6810
rect 20038 6770 20068 6810
rect 19968 6710 20068 6770
rect 19968 6670 19998 6710
rect 20038 6670 20068 6710
rect 19968 6610 20068 6670
rect 19968 6570 19998 6610
rect 20038 6570 20068 6610
rect 19968 6540 20068 6570
rect 20188 6910 20288 6940
rect 20188 6870 20218 6910
rect 20258 6870 20288 6910
rect 20188 6810 20288 6870
rect 20188 6770 20218 6810
rect 20258 6770 20288 6810
rect 20188 6710 20288 6770
rect 20188 6670 20218 6710
rect 20258 6670 20288 6710
rect 20188 6610 20288 6670
rect 20188 6570 20218 6610
rect 20258 6570 20288 6610
rect 20188 6540 20288 6570
rect 20408 6910 20508 6940
rect 20408 6870 20438 6910
rect 20478 6870 20508 6910
rect 20408 6810 20508 6870
rect 20408 6770 20438 6810
rect 20478 6770 20508 6810
rect 20408 6710 20508 6770
rect 20408 6670 20438 6710
rect 20478 6670 20508 6710
rect 20408 6610 20508 6670
rect 20408 6570 20438 6610
rect 20478 6570 20508 6610
rect 20408 6540 20508 6570
rect 20628 6910 20728 6940
rect 20628 6870 20658 6910
rect 20698 6870 20728 6910
rect 20628 6810 20728 6870
rect 20628 6770 20658 6810
rect 20698 6770 20728 6810
rect 20628 6710 20728 6770
rect 20628 6670 20658 6710
rect 20698 6670 20728 6710
rect 20628 6610 20728 6670
rect 20628 6570 20658 6610
rect 20698 6570 20728 6610
rect 20628 6540 20728 6570
rect 20848 6910 20948 6940
rect 21048 6910 21148 6940
rect 20848 6870 20878 6910
rect 20918 6870 20948 6910
rect 21048 6870 21078 6910
rect 21118 6870 21148 6910
rect 20848 6810 20948 6870
rect 21048 6810 21148 6870
rect 20848 6770 20878 6810
rect 20918 6770 20948 6810
rect 21048 6770 21078 6810
rect 21118 6770 21148 6810
rect 20848 6710 20948 6770
rect 21048 6710 21148 6770
rect 20848 6670 20878 6710
rect 20918 6670 20948 6710
rect 21048 6670 21078 6710
rect 21118 6670 21148 6710
rect 20848 6610 20948 6670
rect 21048 6610 21148 6670
rect 20848 6570 20878 6610
rect 20918 6570 20948 6610
rect 21048 6570 21078 6610
rect 21118 6570 21148 6610
rect 20848 6540 20948 6570
rect 21048 6540 21148 6570
rect 21268 6910 21368 6940
rect 21268 6870 21298 6910
rect 21338 6870 21368 6910
rect 21268 6810 21368 6870
rect 21268 6770 21298 6810
rect 21338 6770 21368 6810
rect 21268 6710 21368 6770
rect 21268 6670 21298 6710
rect 21338 6670 21368 6710
rect 21268 6610 21368 6670
rect 21268 6570 21298 6610
rect 21338 6570 21368 6610
rect 21268 6540 21368 6570
rect 21488 6910 21588 6940
rect 21488 6870 21518 6910
rect 21558 6870 21588 6910
rect 21488 6810 21588 6870
rect 21488 6770 21518 6810
rect 21558 6770 21588 6810
rect 21488 6710 21588 6770
rect 21488 6670 21518 6710
rect 21558 6670 21588 6710
rect 21488 6610 21588 6670
rect 21488 6570 21518 6610
rect 21558 6570 21588 6610
rect 21488 6540 21588 6570
rect 21708 6910 21808 6940
rect 21708 6870 21738 6910
rect 21778 6870 21808 6910
rect 21708 6810 21808 6870
rect 21708 6770 21738 6810
rect 21778 6770 21808 6810
rect 21708 6710 21808 6770
rect 21708 6670 21738 6710
rect 21778 6670 21808 6710
rect 21708 6610 21808 6670
rect 21708 6570 21738 6610
rect 21778 6570 21808 6610
rect 21708 6540 21808 6570
rect 21928 6910 22028 6940
rect 21928 6870 21958 6910
rect 21998 6870 22028 6910
rect 21928 6810 22028 6870
rect 21928 6770 21958 6810
rect 21998 6770 22028 6810
rect 21928 6710 22028 6770
rect 21928 6670 21958 6710
rect 21998 6670 22028 6710
rect 21928 6610 22028 6670
rect 21928 6570 21958 6610
rect 21998 6570 22028 6610
rect 21928 6540 22028 6570
rect 22148 6910 22248 6940
rect 22148 6870 22178 6910
rect 22218 6870 22248 6910
rect 22148 6810 22248 6870
rect 22148 6770 22178 6810
rect 22218 6770 22248 6810
rect 22148 6710 22248 6770
rect 22148 6670 22178 6710
rect 22218 6670 22248 6710
rect 22148 6610 22248 6670
rect 22148 6570 22178 6610
rect 22218 6570 22248 6610
rect 22148 6540 22248 6570
rect 22368 6910 22468 6940
rect 22368 6870 22398 6910
rect 22438 6870 22468 6910
rect 22368 6810 22468 6870
rect 22368 6770 22398 6810
rect 22438 6770 22468 6810
rect 22368 6710 22468 6770
rect 22368 6670 22398 6710
rect 22438 6670 22468 6710
rect 22368 6610 22468 6670
rect 22368 6570 22398 6610
rect 22438 6570 22468 6610
rect 22368 6540 22468 6570
rect 17968 6510 18068 6540
rect 23198 5400 23278 5430
rect 23198 5360 23218 5400
rect 23258 5360 23278 5400
rect 23198 5300 23278 5360
rect 23198 5260 23218 5300
rect 23258 5260 23278 5300
rect 23198 5200 23278 5260
rect 23198 5160 23218 5200
rect 23258 5160 23278 5200
rect 23198 5100 23278 5160
rect 23198 5060 23218 5100
rect 23258 5060 23278 5100
rect 23198 5030 23278 5060
rect 23578 5400 23658 5430
rect 23578 5360 23598 5400
rect 23638 5360 23658 5400
rect 23578 5300 23658 5360
rect 23578 5260 23598 5300
rect 23638 5260 23658 5300
rect 23578 5200 23658 5260
rect 23578 5160 23598 5200
rect 23638 5160 23658 5200
rect 23578 5100 23658 5160
rect 23578 5060 23598 5100
rect 23638 5060 23658 5100
rect 23578 5030 23658 5060
rect 23718 5400 23798 5430
rect 23718 5360 23738 5400
rect 23778 5360 23798 5400
rect 23718 5300 23798 5360
rect 23718 5260 23738 5300
rect 23778 5260 23798 5300
rect 23718 5200 23798 5260
rect 23718 5160 23738 5200
rect 23778 5160 23798 5200
rect 23718 5100 23798 5160
rect 23718 5060 23738 5100
rect 23778 5060 23798 5100
rect 23718 5030 23798 5060
rect 24098 5400 24178 5430
rect 24098 5360 24118 5400
rect 24158 5360 24178 5400
rect 24098 5300 24178 5360
rect 24098 5260 24118 5300
rect 24158 5260 24178 5300
rect 24098 5200 24178 5260
rect 24098 5160 24118 5200
rect 24158 5160 24178 5200
rect 24098 5100 24178 5160
rect 24098 5060 24118 5100
rect 24158 5060 24178 5100
rect 24098 5030 24178 5060
rect 24238 5400 24318 5430
rect 24238 5360 24258 5400
rect 24298 5360 24318 5400
rect 24238 5300 24318 5360
rect 24238 5260 24258 5300
rect 24298 5260 24318 5300
rect 24238 5200 24318 5260
rect 24238 5160 24258 5200
rect 24298 5160 24318 5200
rect 24238 5100 24318 5160
rect 24238 5060 24258 5100
rect 24298 5060 24318 5100
rect 24238 5030 24318 5060
rect 24618 5400 24698 5430
rect 24618 5360 24638 5400
rect 24678 5360 24698 5400
rect 24618 5300 24698 5360
rect 24618 5260 24638 5300
rect 24678 5260 24698 5300
rect 24618 5200 24698 5260
rect 24618 5160 24638 5200
rect 24678 5160 24698 5200
rect 24618 5100 24698 5160
rect 24618 5060 24638 5100
rect 24678 5060 24698 5100
rect 24618 5030 24698 5060
rect 24758 5400 24838 5430
rect 24758 5360 24778 5400
rect 24818 5360 24838 5400
rect 24758 5300 24838 5360
rect 24758 5260 24778 5300
rect 24818 5260 24838 5300
rect 24758 5200 24838 5260
rect 24758 5160 24778 5200
rect 24818 5160 24838 5200
rect 24758 5100 24838 5160
rect 24758 5060 24778 5100
rect 24818 5060 24838 5100
rect 24758 5030 24838 5060
rect 25138 5400 25218 5430
rect 25138 5360 25158 5400
rect 25198 5360 25218 5400
rect 25138 5300 25218 5360
rect 25138 5260 25158 5300
rect 25198 5260 25218 5300
rect 25138 5200 25218 5260
rect 25138 5160 25158 5200
rect 25198 5160 25218 5200
rect 25138 5100 25218 5160
rect 25138 5060 25158 5100
rect 25198 5060 25218 5100
rect 25138 5030 25218 5060
rect 12588 3500 12668 3530
rect 12588 3460 12608 3500
rect 12648 3460 12668 3500
rect 12588 3430 12668 3460
rect 12698 3500 12778 3530
rect 12698 3460 12718 3500
rect 12758 3460 12778 3500
rect 12698 3430 12778 3460
rect 13008 3500 13088 3530
rect 13008 3460 13028 3500
rect 13068 3460 13088 3500
rect 13008 3430 13088 3460
rect 13118 3500 13198 3530
rect 13118 3460 13138 3500
rect 13178 3460 13198 3500
rect 13118 3430 13198 3460
rect 13228 3500 13308 3530
rect 13228 3460 13248 3500
rect 13288 3460 13308 3500
rect 13228 3430 13308 3460
rect 13678 3500 13758 3530
rect 13678 3460 13698 3500
rect 13738 3460 13758 3500
rect 13678 3430 13758 3460
rect 13788 3500 13868 3530
rect 13788 3460 13808 3500
rect 13848 3460 13868 3500
rect 13788 3430 13868 3460
rect 13898 3500 13978 3530
rect 13898 3460 13918 3500
rect 13958 3460 13978 3500
rect 13898 3430 13978 3460
rect 14118 3500 14198 3530
rect 14118 3460 14138 3500
rect 14178 3460 14198 3500
rect 14118 3430 14198 3460
rect 14228 3500 14308 3530
rect 14228 3460 14248 3500
rect 14288 3460 14308 3500
rect 14228 3430 14308 3460
rect 14338 3500 14418 3530
rect 14338 3460 14358 3500
rect 14398 3460 14418 3500
rect 14338 3430 14418 3460
rect 14448 3500 14528 3530
rect 14448 3460 14468 3500
rect 14508 3460 14528 3500
rect 14448 3430 14528 3460
rect 14958 3500 15038 3530
rect 14958 3460 14978 3500
rect 15018 3460 15038 3500
rect 14958 3430 15038 3460
rect 15068 3500 15148 3530
rect 15068 3460 15088 3500
rect 15128 3460 15148 3500
rect 15068 3430 15148 3460
rect 15378 3500 15458 3530
rect 15378 3460 15398 3500
rect 15438 3460 15458 3500
rect 15378 3430 15458 3460
rect 15488 3500 15568 3530
rect 15488 3460 15508 3500
rect 15548 3460 15568 3500
rect 15488 3430 15568 3460
rect 15598 3500 15678 3530
rect 15598 3460 15618 3500
rect 15658 3460 15678 3500
rect 15598 3430 15678 3460
rect 15828 3500 15908 3530
rect 15828 3460 15848 3500
rect 15888 3460 15908 3500
rect 15828 3430 15908 3460
rect 15938 3500 16018 3530
rect 15938 3460 15958 3500
rect 15998 3460 16018 3500
rect 15938 3430 16018 3460
rect 16048 3500 16128 3530
rect 16048 3460 16068 3500
rect 16108 3460 16128 3500
rect 16048 3430 16128 3460
rect 16188 3500 16268 3530
rect 16188 3460 16208 3500
rect 16248 3460 16268 3500
rect 16188 3430 16268 3460
rect 16298 3500 16378 3530
rect 16298 3460 16318 3500
rect 16358 3460 16378 3500
rect 16298 3430 16378 3460
rect 16408 3500 16488 3530
rect 16408 3460 16428 3500
rect 16468 3460 16488 3500
rect 16408 3430 16488 3460
rect 16768 3500 16848 3530
rect 16768 3460 16788 3500
rect 16828 3460 16848 3500
rect 16768 3430 16848 3460
rect 16878 3500 16958 3530
rect 16878 3460 16898 3500
rect 16938 3460 16958 3500
rect 16878 3430 16958 3460
rect 16988 3500 17068 3530
rect 16988 3460 17008 3500
rect 17048 3460 17068 3500
rect 16988 3430 17068 3460
rect 17208 3500 17288 3530
rect 17208 3460 17228 3500
rect 17268 3460 17288 3500
rect 17208 3430 17288 3460
rect 17318 3500 17398 3530
rect 17318 3460 17338 3500
rect 17378 3460 17398 3500
rect 17318 3430 17398 3460
rect 17428 3500 17508 3530
rect 17428 3460 17448 3500
rect 17488 3460 17508 3500
rect 17428 3430 17508 3460
rect 17828 3500 17908 3530
rect 17828 3460 17848 3500
rect 17888 3460 17908 3500
rect 17828 3430 17908 3460
rect 17938 3500 18018 3530
rect 17938 3460 17958 3500
rect 17998 3460 18018 3500
rect 17938 3430 18018 3460
rect 18168 3500 18248 3530
rect 18168 3460 18188 3500
rect 18228 3460 18248 3500
rect 18168 3430 18248 3460
rect 18278 3500 18358 3530
rect 18278 3460 18298 3500
rect 18338 3460 18358 3500
rect 18278 3430 18358 3460
rect 18388 3500 18468 3530
rect 18388 3460 18408 3500
rect 18448 3460 18468 3500
rect 18388 3430 18468 3460
rect 18528 3500 18608 3530
rect 18528 3460 18548 3500
rect 18588 3460 18608 3500
rect 18528 3430 18608 3460
rect 18638 3500 18718 3530
rect 18638 3460 18658 3500
rect 18698 3460 18718 3500
rect 18638 3430 18718 3460
rect 18748 3500 18828 3530
rect 18748 3460 18768 3500
rect 18808 3460 18828 3500
rect 18748 3430 18828 3460
rect 19128 3500 19208 3530
rect 19128 3460 19148 3500
rect 19188 3460 19208 3500
rect 19128 3430 19208 3460
rect 19238 3500 19318 3530
rect 19238 3460 19258 3500
rect 19298 3460 19318 3500
rect 19238 3430 19318 3460
rect 19468 3500 19548 3530
rect 19468 3460 19488 3500
rect 19528 3460 19548 3500
rect 19468 3430 19548 3460
rect 19578 3500 19658 3530
rect 19578 3460 19598 3500
rect 19638 3460 19658 3500
rect 19578 3430 19658 3460
rect 19688 3500 19768 3530
rect 19688 3460 19708 3500
rect 19748 3460 19768 3500
rect 19688 3430 19768 3460
rect 19828 3500 19908 3530
rect 19828 3460 19848 3500
rect 19888 3460 19908 3500
rect 19828 3430 19908 3460
rect 19938 3500 20018 3530
rect 19938 3460 19958 3500
rect 19998 3460 20018 3500
rect 19938 3430 20018 3460
rect 20048 3500 20128 3530
rect 20048 3460 20068 3500
rect 20108 3460 20128 3500
rect 20048 3430 20128 3460
rect 20428 3500 20508 3530
rect 20428 3460 20448 3500
rect 20488 3460 20508 3500
rect 20428 3430 20508 3460
rect 20538 3500 20618 3530
rect 20538 3460 20558 3500
rect 20598 3460 20618 3500
rect 20538 3430 20618 3460
rect 20768 3500 20848 3530
rect 20768 3460 20788 3500
rect 20828 3460 20848 3500
rect 20768 3430 20848 3460
rect 20878 3500 20958 3530
rect 20878 3460 20898 3500
rect 20938 3460 20958 3500
rect 20878 3430 20958 3460
rect 20988 3500 21068 3530
rect 20988 3460 21008 3500
rect 21048 3460 21068 3500
rect 20988 3430 21068 3460
rect 21128 3500 21208 3530
rect 21128 3460 21148 3500
rect 21188 3460 21208 3500
rect 21128 3430 21208 3460
rect 21238 3500 21318 3530
rect 21238 3460 21258 3500
rect 21298 3460 21318 3500
rect 21238 3430 21318 3460
rect 21348 3500 21428 3530
rect 21348 3460 21368 3500
rect 21408 3460 21428 3500
rect 21348 3430 21428 3460
rect 21728 3500 21808 3530
rect 21728 3460 21748 3500
rect 21788 3460 21808 3500
rect 21728 3430 21808 3460
rect 21838 3500 21918 3530
rect 21838 3460 21858 3500
rect 21898 3460 21918 3500
rect 21838 3430 21918 3460
rect 22068 3500 22148 3530
rect 22068 3460 22088 3500
rect 22128 3460 22148 3500
rect 22068 3430 22148 3460
rect 22178 3500 22258 3530
rect 22178 3460 22198 3500
rect 22238 3460 22258 3500
rect 22178 3430 22258 3460
rect 22288 3500 22368 3530
rect 22288 3460 22308 3500
rect 22348 3460 22368 3500
rect 22288 3430 22368 3460
rect 22428 3500 22508 3530
rect 22428 3460 22448 3500
rect 22488 3460 22508 3500
rect 22428 3430 22508 3460
rect 22538 3500 22618 3530
rect 22538 3460 22558 3500
rect 22598 3460 22618 3500
rect 22538 3430 22618 3460
rect 22648 3500 22728 3530
rect 22648 3460 22668 3500
rect 22708 3460 22728 3500
rect 22648 3430 22728 3460
rect 23198 4710 23278 4740
rect 23198 4670 23218 4710
rect 23258 4670 23278 4710
rect 23198 4610 23278 4670
rect 23198 4570 23218 4610
rect 23258 4570 23278 4610
rect 23198 4510 23278 4570
rect 23198 4470 23218 4510
rect 23258 4470 23278 4510
rect 23198 4410 23278 4470
rect 23198 4370 23218 4410
rect 23258 4370 23278 4410
rect 23198 4310 23278 4370
rect 23198 4270 23218 4310
rect 23258 4270 23278 4310
rect 23198 4210 23278 4270
rect 23198 4170 23218 4210
rect 23258 4170 23278 4210
rect 23198 4140 23278 4170
rect 23308 4710 23388 4740
rect 23308 4670 23328 4710
rect 23368 4670 23388 4710
rect 23308 4610 23388 4670
rect 23308 4570 23328 4610
rect 23368 4570 23388 4610
rect 23308 4510 23388 4570
rect 23308 4470 23328 4510
rect 23368 4470 23388 4510
rect 23308 4410 23388 4470
rect 23308 4370 23328 4410
rect 23368 4370 23388 4410
rect 23308 4310 23388 4370
rect 23308 4270 23328 4310
rect 23368 4270 23388 4310
rect 23308 4210 23388 4270
rect 23308 4170 23328 4210
rect 23368 4170 23388 4210
rect 23308 4140 23388 4170
rect 23718 4710 23798 4740
rect 23718 4670 23738 4710
rect 23778 4670 23798 4710
rect 23718 4610 23798 4670
rect 23718 4570 23738 4610
rect 23778 4570 23798 4610
rect 23718 4510 23798 4570
rect 23718 4470 23738 4510
rect 23778 4470 23798 4510
rect 23718 4410 23798 4470
rect 23718 4370 23738 4410
rect 23778 4370 23798 4410
rect 23718 4310 23798 4370
rect 23718 4270 23738 4310
rect 23778 4270 23798 4310
rect 23718 4210 23798 4270
rect 23718 4170 23738 4210
rect 23778 4170 23798 4210
rect 23718 4140 23798 4170
rect 23828 4710 23908 4740
rect 23828 4670 23848 4710
rect 23888 4670 23908 4710
rect 23828 4610 23908 4670
rect 23828 4570 23848 4610
rect 23888 4570 23908 4610
rect 23828 4510 23908 4570
rect 23828 4470 23848 4510
rect 23888 4470 23908 4510
rect 23828 4410 23908 4470
rect 23828 4370 23848 4410
rect 23888 4370 23908 4410
rect 23828 4310 23908 4370
rect 23828 4270 23848 4310
rect 23888 4270 23908 4310
rect 23828 4210 23908 4270
rect 23828 4170 23848 4210
rect 23888 4170 23908 4210
rect 23828 4140 23908 4170
rect 24238 4710 24318 4740
rect 24238 4670 24258 4710
rect 24298 4670 24318 4710
rect 24238 4610 24318 4670
rect 24238 4570 24258 4610
rect 24298 4570 24318 4610
rect 24238 4510 24318 4570
rect 24238 4470 24258 4510
rect 24298 4470 24318 4510
rect 24238 4410 24318 4470
rect 24238 4370 24258 4410
rect 24298 4370 24318 4410
rect 24238 4310 24318 4370
rect 24238 4270 24258 4310
rect 24298 4270 24318 4310
rect 24238 4210 24318 4270
rect 24238 4170 24258 4210
rect 24298 4170 24318 4210
rect 24238 4140 24318 4170
rect 24348 4710 24428 4740
rect 24348 4670 24368 4710
rect 24408 4670 24428 4710
rect 24348 4610 24428 4670
rect 24348 4570 24368 4610
rect 24408 4570 24428 4610
rect 24348 4510 24428 4570
rect 24348 4470 24368 4510
rect 24408 4470 24428 4510
rect 24348 4410 24428 4470
rect 24348 4370 24368 4410
rect 24408 4370 24428 4410
rect 24348 4310 24428 4370
rect 24348 4270 24368 4310
rect 24408 4270 24428 4310
rect 24348 4210 24428 4270
rect 24348 4170 24368 4210
rect 24408 4170 24428 4210
rect 24348 4140 24428 4170
rect 23196 3930 23276 3960
rect 23196 3890 23216 3930
rect 23256 3890 23276 3930
rect 23196 3830 23276 3890
rect 23196 3790 23216 3830
rect 23256 3790 23276 3830
rect 23196 3730 23276 3790
rect 23196 3690 23216 3730
rect 23256 3690 23276 3730
rect 23196 3630 23276 3690
rect 23196 3590 23216 3630
rect 23256 3590 23276 3630
rect 23196 3560 23276 3590
rect 23308 3930 23388 3960
rect 23308 3890 23328 3930
rect 23368 3890 23388 3930
rect 23308 3830 23388 3890
rect 23308 3790 23328 3830
rect 23368 3790 23388 3830
rect 23308 3730 23388 3790
rect 23308 3690 23328 3730
rect 23368 3690 23388 3730
rect 23308 3630 23388 3690
rect 23308 3590 23328 3630
rect 23368 3590 23388 3630
rect 23308 3560 23388 3590
rect 23716 3930 23796 3960
rect 23716 3890 23736 3930
rect 23776 3890 23796 3930
rect 23716 3830 23796 3890
rect 23716 3790 23736 3830
rect 23776 3790 23796 3830
rect 23716 3730 23796 3790
rect 23716 3690 23736 3730
rect 23776 3690 23796 3730
rect 23716 3630 23796 3690
rect 23716 3590 23736 3630
rect 23776 3590 23796 3630
rect 23716 3560 23796 3590
rect 23828 3930 23908 3960
rect 23828 3890 23848 3930
rect 23888 3890 23908 3930
rect 23828 3830 23908 3890
rect 23828 3790 23848 3830
rect 23888 3790 23908 3830
rect 23828 3730 23908 3790
rect 23828 3690 23848 3730
rect 23888 3690 23908 3730
rect 23828 3630 23908 3690
rect 23828 3590 23848 3630
rect 23888 3590 23908 3630
rect 23828 3560 23908 3590
rect 24236 3930 24316 3960
rect 24236 3890 24256 3930
rect 24296 3890 24316 3930
rect 24236 3830 24316 3890
rect 24236 3790 24256 3830
rect 24296 3790 24316 3830
rect 24236 3730 24316 3790
rect 24236 3690 24256 3730
rect 24296 3690 24316 3730
rect 24236 3630 24316 3690
rect 24236 3590 24256 3630
rect 24296 3590 24316 3630
rect 24236 3560 24316 3590
rect 24348 3930 24428 3960
rect 24348 3890 24368 3930
rect 24408 3890 24428 3930
rect 24348 3830 24428 3890
rect 24348 3790 24368 3830
rect 24408 3790 24428 3830
rect 24348 3730 24428 3790
rect 24348 3690 24368 3730
rect 24408 3690 24428 3730
rect 24348 3630 24428 3690
rect 24348 3590 24368 3630
rect 24408 3590 24428 3630
rect 24348 3560 24428 3590
<< ndiffc >>
rect 11178 14210 11218 14250
rect 11178 14110 11218 14150
rect 13258 14210 13298 14250
rect 13258 14110 13298 14150
rect 15338 14210 15378 14250
rect 15338 14110 15378 14150
rect 10758 13600 10798 13640
rect 10758 13500 10798 13540
rect 10758 13400 10798 13440
rect 10758 13300 10798 13340
rect 10758 13200 10798 13240
rect 11838 13600 11878 13640
rect 11998 13600 12038 13640
rect 11838 13500 11878 13540
rect 11998 13500 12038 13540
rect 11838 13400 11878 13440
rect 11998 13400 12038 13440
rect 11838 13300 11878 13340
rect 11998 13300 12038 13340
rect 11838 13200 11878 13240
rect 11998 13200 12038 13240
rect 13078 13600 13118 13640
rect 13078 13500 13118 13540
rect 13078 13400 13118 13440
rect 13078 13300 13118 13340
rect 13078 13200 13118 13240
rect 13438 13600 13478 13640
rect 13438 13500 13478 13540
rect 13438 13400 13478 13440
rect 13438 13300 13478 13340
rect 13438 13200 13478 13240
rect 14518 13600 14558 13640
rect 14678 13600 14718 13640
rect 14518 13500 14558 13540
rect 14678 13500 14718 13540
rect 14518 13400 14558 13440
rect 14678 13400 14718 13440
rect 14518 13300 14558 13340
rect 14678 13300 14718 13340
rect 14518 13200 14558 13240
rect 14678 13200 14718 13240
rect 15758 13600 15798 13640
rect 15758 13500 15798 13540
rect 15758 13400 15798 13440
rect 15758 13300 15798 13340
rect 15758 13200 15798 13240
rect 11378 12590 11418 12630
rect 11498 12590 11538 12630
rect 11618 12590 11658 12630
rect 11738 12590 11778 12630
rect 11858 12590 11898 12630
rect 11978 12590 12018 12630
rect 12098 12590 12138 12630
rect 12218 12590 12258 12630
rect 12338 12590 12378 12630
rect 12458 12590 12498 12630
rect 12578 12590 12618 12630
rect 13938 12590 13978 12630
rect 14058 12590 14098 12630
rect 14178 12590 14218 12630
rect 14298 12590 14338 12630
rect 14418 12590 14458 12630
rect 14538 12590 14578 12630
rect 14658 12590 14698 12630
rect 14778 12590 14818 12630
rect 14898 12590 14938 12630
rect 15018 12590 15058 12630
rect 15138 12590 15178 12630
rect 19468 10990 19508 11030
rect 19598 10990 19638 11030
rect 19728 10990 19768 11030
rect 19858 10990 19898 11030
rect 19988 10990 20028 11030
rect 20118 10990 20158 11030
rect 20248 10990 20288 11030
rect 20608 10990 20648 11030
rect 20738 10990 20778 11030
rect 20868 10990 20908 11030
rect 20998 10990 21038 11030
rect 21128 10990 21168 11030
rect 21258 10990 21298 11030
rect 21388 10990 21428 11030
rect 21748 10990 21788 11030
rect 21878 10990 21918 11030
rect 22008 10990 22048 11030
rect 22138 10990 22178 11030
rect 22268 10990 22308 11030
rect 22398 10990 22438 11030
rect 22528 10990 22568 11030
rect 19418 10440 19458 10490
rect 19418 10300 19458 10350
rect 19618 10440 19658 10490
rect 19618 10300 19658 10350
rect 19818 10440 19858 10490
rect 19818 10300 19858 10350
rect 20018 10440 20058 10490
rect 20018 10300 20058 10350
rect 20218 10440 20258 10490
rect 20218 10300 20258 10350
rect 20418 10440 20458 10490
rect 20418 10300 20458 10350
rect 20618 10440 20658 10490
rect 20618 10300 20658 10350
rect 20818 10440 20858 10490
rect 20818 10300 20858 10350
rect 21018 10440 21058 10490
rect 21018 10300 21058 10350
rect 21218 10440 21258 10490
rect 21218 10300 21258 10350
rect 21418 10440 21458 10490
rect 21418 10300 21458 10350
rect 13268 8020 13308 8060
rect 13268 7920 13308 7960
rect 13378 8020 13418 8060
rect 13378 7920 13418 7960
rect 13488 8020 13528 8060
rect 13488 7920 13528 7960
rect 13788 8020 13828 8060
rect 13788 7920 13828 7960
rect 13898 8020 13938 8060
rect 13898 7920 13938 7960
rect 14008 8020 14048 8060
rect 14168 8020 14208 8060
rect 14008 7920 14048 7960
rect 14168 7920 14208 7960
rect 14278 8020 14318 8060
rect 14278 7920 14318 7960
rect 14388 8020 14428 8060
rect 14388 7920 14428 7960
rect 14688 8020 14728 8060
rect 14688 7920 14728 7960
rect 14798 8020 14838 8060
rect 14798 7920 14838 7960
rect 14908 8020 14948 8060
rect 14908 7920 14948 7960
rect 15198 8020 15238 8060
rect 15198 7920 15238 7960
rect 15308 8020 15348 8060
rect 15308 7920 15348 7960
rect 15528 8020 15568 8060
rect 15528 7920 15568 7960
rect 15638 8020 15678 8060
rect 15638 7920 15678 7960
rect 15858 8020 15898 8060
rect 15858 7920 15898 7960
rect 15968 8020 16008 8060
rect 15968 7920 16008 7960
rect 16408 8020 16448 8060
rect 16408 7920 16448 7960
rect 16538 8020 16578 8060
rect 16538 7920 16578 7960
rect 16798 8020 16838 8060
rect 16798 7920 16838 7960
rect 16928 8020 16968 8060
rect 16928 7920 16968 7960
rect 17188 8020 17228 8060
rect 17188 7920 17228 7960
rect 17318 8020 17358 8060
rect 17318 7920 17358 7960
rect 17478 8020 17518 8060
rect 17478 7920 17518 7960
rect 17608 8020 17648 8060
rect 17608 7920 17648 7960
rect 17868 8020 17908 8060
rect 17868 7920 17908 7960
rect 17998 8020 18038 8060
rect 17998 7920 18038 7960
rect 19358 7970 19398 8010
rect 19358 7870 19398 7910
rect 19358 7770 19398 7810
rect 19358 7670 19398 7710
rect 19578 7970 19618 8010
rect 19578 7870 19618 7910
rect 19578 7770 19618 7810
rect 19578 7670 19618 7710
rect 19798 7970 19838 8010
rect 19798 7870 19838 7910
rect 19798 7770 19838 7810
rect 19798 7670 19838 7710
rect 20018 7970 20058 8010
rect 20018 7870 20058 7910
rect 20018 7770 20058 7810
rect 20018 7670 20058 7710
rect 20238 7970 20278 8010
rect 20438 7970 20478 8010
rect 20238 7870 20278 7910
rect 20438 7870 20478 7910
rect 20238 7770 20278 7810
rect 20438 7770 20478 7810
rect 20238 7670 20278 7710
rect 20438 7670 20478 7710
rect 20658 7970 20698 8010
rect 20658 7870 20698 7910
rect 20658 7770 20698 7810
rect 20658 7670 20698 7710
rect 20878 7970 20918 8010
rect 20878 7870 20918 7910
rect 20878 7770 20918 7810
rect 20878 7670 20918 7710
rect 21098 7970 21138 8010
rect 21098 7870 21138 7910
rect 21098 7770 21138 7810
rect 21098 7670 21138 7710
rect 21318 7970 21358 8010
rect 21518 7970 21558 8010
rect 21318 7870 21358 7910
rect 21518 7870 21558 7910
rect 21318 7770 21358 7810
rect 21518 7770 21558 7810
rect 21318 7670 21358 7710
rect 21518 7670 21558 7710
rect 21738 7970 21778 8010
rect 21738 7870 21778 7910
rect 21738 7770 21778 7810
rect 21738 7670 21778 7710
rect 21958 7970 21998 8010
rect 21958 7870 21998 7910
rect 21958 7770 21998 7810
rect 21958 7670 21998 7710
rect 22178 7970 22218 8010
rect 22178 7870 22218 7910
rect 22178 7770 22218 7810
rect 22178 7670 22218 7710
rect 22398 7970 22438 8010
rect 22398 7870 22438 7910
rect 22398 7770 22438 7810
rect 22398 7670 22438 7710
rect 13268 6220 13308 6260
rect 13268 6120 13308 6160
rect 13378 6220 13418 6260
rect 13378 6120 13418 6160
rect 13488 6220 13528 6260
rect 13488 6120 13528 6160
rect 13788 6220 13828 6260
rect 13788 6120 13828 6160
rect 13898 6220 13938 6260
rect 13898 6120 13938 6160
rect 14008 6220 14048 6260
rect 14168 6220 14208 6260
rect 14008 6120 14048 6160
rect 14168 6120 14208 6160
rect 14278 6220 14318 6260
rect 14278 6120 14318 6160
rect 14388 6220 14428 6260
rect 14388 6120 14428 6160
rect 14688 6220 14728 6260
rect 14688 6120 14728 6160
rect 14798 6220 14838 6260
rect 14798 6120 14838 6160
rect 14908 6220 14948 6260
rect 14908 6120 14948 6160
rect 15208 6220 15248 6260
rect 15208 6120 15248 6160
rect 15318 6220 15358 6260
rect 15318 6120 15358 6160
rect 15428 6220 15468 6260
rect 15428 6120 15468 6160
rect 15648 6220 15688 6260
rect 15648 6120 15688 6160
rect 15758 6220 15798 6260
rect 15758 6120 15798 6160
rect 15978 6220 16018 6260
rect 15978 6120 16018 6160
rect 16088 6220 16128 6260
rect 16088 6120 16128 6160
rect 16408 6220 16448 6260
rect 16408 6120 16448 6160
rect 16538 6220 16578 6260
rect 16538 6120 16578 6160
rect 16798 6220 16838 6260
rect 16798 6120 16838 6160
rect 16928 6220 16968 6260
rect 16928 6120 16968 6160
rect 17188 6220 17228 6260
rect 17188 6120 17228 6160
rect 17318 6220 17358 6260
rect 17318 6120 17358 6160
rect 17478 6220 17518 6260
rect 17478 6120 17518 6160
rect 17608 6220 17648 6260
rect 17608 6120 17648 6160
rect 12448 3140 12488 3180
rect 12558 3140 12598 3180
rect 12668 3140 12708 3180
rect 12778 3140 12818 3180
rect 12888 3140 12928 3180
rect 13028 3140 13068 3180
rect 13138 3140 13178 3180
rect 13248 3140 13288 3180
rect 13478 3140 13518 3180
rect 13588 3140 13628 3180
rect 13698 3140 13738 3180
rect 13808 3140 13848 3180
rect 13918 3140 13958 3180
rect 14138 3140 14178 3180
rect 14248 3140 14288 3180
rect 14358 3140 14398 3180
rect 14468 3140 14508 3180
rect 14578 3140 14618 3180
rect 14818 3140 14858 3180
rect 14928 3140 14968 3180
rect 15038 3140 15078 3180
rect 15148 3140 15188 3180
rect 15258 3140 15298 3180
rect 15398 3140 15438 3180
rect 15508 3140 15548 3180
rect 15618 3140 15658 3180
rect 15958 3140 15998 3180
rect 16068 3140 16108 3180
rect 16318 3140 16358 3180
rect 16428 3140 16468 3180
rect 16568 3140 16608 3180
rect 16678 3140 16718 3180
rect 16788 3140 16828 3180
rect 16898 3140 16938 3180
rect 17008 3140 17048 3180
rect 17228 3140 17268 3180
rect 17338 3140 17378 3180
rect 17448 3140 17488 3180
rect 17558 3140 17598 3180
rect 17778 3140 17818 3180
rect 17888 3140 17928 3180
rect 17998 3140 18038 3180
rect 18108 3140 18148 3180
rect 18218 3140 18258 3180
rect 18438 3140 18478 3180
rect 18548 3140 18588 3180
rect 18658 3140 18698 3180
rect 18768 3140 18808 3180
rect 19078 3050 19118 3090
rect 19188 3050 19228 3090
rect 19298 3050 19338 3090
rect 19408 3050 19448 3090
rect 19518 3050 19558 3090
rect 19738 3050 19778 3090
rect 19848 3050 19888 3090
rect 19958 3050 19998 3090
rect 20068 3050 20108 3090
rect 20378 3050 20418 3090
rect 20488 3050 20528 3090
rect 20598 3050 20638 3090
rect 20708 3050 20748 3090
rect 20818 3050 20858 3090
rect 21038 3050 21078 3090
rect 21148 3050 21188 3090
rect 21258 3050 21298 3090
rect 21368 3050 21408 3090
rect 21678 3050 21718 3090
rect 21788 3050 21828 3090
rect 21898 3050 21938 3090
rect 22008 3050 22048 3090
rect 22118 3050 22158 3090
rect 22338 3050 22378 3090
rect 22448 3050 22488 3090
rect 22558 3050 22598 3090
rect 22668 3050 22708 3090
rect 23216 2970 23256 3010
rect 23216 2870 23256 2910
rect 23328 2970 23368 3010
rect 23328 2870 23368 2910
rect 23736 2970 23776 3010
rect 23736 2870 23776 2910
rect 23848 2970 23888 3010
rect 23848 2870 23888 2910
rect 24256 2970 24296 3010
rect 24256 2870 24296 2910
rect 24368 2970 24408 3010
rect 24368 2870 24408 2910
rect 23218 2590 23258 2630
rect 23218 2490 23258 2530
rect 23218 2390 23258 2430
rect 23328 2590 23368 2630
rect 23328 2490 23368 2530
rect 23328 2390 23368 2430
rect 23738 2590 23778 2630
rect 23738 2490 23778 2530
rect 23738 2390 23778 2430
rect 23848 2590 23888 2630
rect 23848 2490 23888 2530
rect 23848 2390 23888 2430
rect 24258 2590 24298 2630
rect 24258 2490 24298 2530
rect 24258 2390 24298 2430
rect 24368 2590 24408 2630
rect 24368 2490 24408 2530
rect 24368 2390 24408 2430
rect 23218 2110 23258 2150
rect 23218 2010 23258 2050
rect 23328 2110 23368 2150
rect 23328 2010 23368 2050
rect 23738 2110 23778 2150
rect 23738 2010 23778 2050
rect 23848 2110 23888 2150
rect 23848 2010 23888 2050
rect 24258 2110 24298 2150
rect 24258 2010 24298 2050
rect 24368 2110 24408 2150
rect 24368 2010 24408 2050
rect 24858 2110 24898 2150
rect 24858 2010 24898 2050
rect 24968 2110 25008 2150
rect 24968 2010 25008 2050
<< pdiffc >>
rect 11630 18392 11664 18426
rect 11720 18392 11754 18426
rect 11810 18392 11844 18426
rect 11900 18392 11934 18426
rect 11990 18392 12024 18426
rect 12080 18392 12114 18426
rect 12170 18392 12204 18426
rect 11630 18302 11664 18336
rect 11720 18302 11754 18336
rect 11810 18302 11844 18336
rect 11900 18302 11934 18336
rect 11990 18302 12024 18336
rect 12080 18302 12114 18336
rect 12170 18302 12204 18336
rect 11630 18212 11664 18246
rect 11720 18212 11754 18246
rect 11810 18212 11844 18246
rect 11900 18212 11934 18246
rect 11990 18212 12024 18246
rect 12080 18212 12114 18246
rect 12170 18212 12204 18246
rect 11630 18122 11664 18156
rect 11720 18122 11754 18156
rect 11810 18122 11844 18156
rect 11900 18122 11934 18156
rect 11990 18122 12024 18156
rect 12080 18122 12114 18156
rect 12170 18122 12204 18156
rect 11630 18032 11664 18066
rect 11720 18032 11754 18066
rect 11810 18032 11844 18066
rect 11900 18032 11934 18066
rect 11990 18032 12024 18066
rect 12080 18032 12114 18066
rect 12170 18032 12204 18066
rect 11630 17942 11664 17976
rect 11720 17942 11754 17976
rect 11810 17942 11844 17976
rect 11900 17942 11934 17976
rect 11990 17942 12024 17976
rect 12080 17942 12114 17976
rect 12170 17942 12204 17976
rect 11630 17852 11664 17886
rect 11720 17852 11754 17886
rect 11810 17852 11844 17886
rect 11900 17852 11934 17886
rect 11990 17852 12024 17886
rect 12080 17852 12114 17886
rect 12170 17852 12204 17886
rect 12990 18392 13024 18426
rect 13080 18392 13114 18426
rect 13170 18392 13204 18426
rect 13260 18392 13294 18426
rect 13350 18392 13384 18426
rect 13440 18392 13474 18426
rect 13530 18392 13564 18426
rect 12990 18302 13024 18336
rect 13080 18302 13114 18336
rect 13170 18302 13204 18336
rect 13260 18302 13294 18336
rect 13350 18302 13384 18336
rect 13440 18302 13474 18336
rect 13530 18302 13564 18336
rect 12990 18212 13024 18246
rect 13080 18212 13114 18246
rect 13170 18212 13204 18246
rect 13260 18212 13294 18246
rect 13350 18212 13384 18246
rect 13440 18212 13474 18246
rect 13530 18212 13564 18246
rect 12990 18122 13024 18156
rect 13080 18122 13114 18156
rect 13170 18122 13204 18156
rect 13260 18122 13294 18156
rect 13350 18122 13384 18156
rect 13440 18122 13474 18156
rect 13530 18122 13564 18156
rect 12990 18032 13024 18066
rect 13080 18032 13114 18066
rect 13170 18032 13204 18066
rect 13260 18032 13294 18066
rect 13350 18032 13384 18066
rect 13440 18032 13474 18066
rect 13530 18032 13564 18066
rect 12990 17942 13024 17976
rect 13080 17942 13114 17976
rect 13170 17942 13204 17976
rect 13260 17942 13294 17976
rect 13350 17942 13384 17976
rect 13440 17942 13474 17976
rect 13530 17942 13564 17976
rect 12990 17852 13024 17886
rect 13080 17852 13114 17886
rect 13170 17852 13204 17886
rect 13260 17852 13294 17886
rect 13350 17852 13384 17886
rect 13440 17852 13474 17886
rect 13530 17852 13564 17886
rect 14350 18392 14384 18426
rect 14440 18392 14474 18426
rect 14530 18392 14564 18426
rect 14620 18392 14654 18426
rect 14710 18392 14744 18426
rect 14800 18392 14834 18426
rect 14890 18392 14924 18426
rect 14350 18302 14384 18336
rect 14440 18302 14474 18336
rect 14530 18302 14564 18336
rect 14620 18302 14654 18336
rect 14710 18302 14744 18336
rect 14800 18302 14834 18336
rect 14890 18302 14924 18336
rect 14350 18212 14384 18246
rect 14440 18212 14474 18246
rect 14530 18212 14564 18246
rect 14620 18212 14654 18246
rect 14710 18212 14744 18246
rect 14800 18212 14834 18246
rect 14890 18212 14924 18246
rect 14350 18122 14384 18156
rect 14440 18122 14474 18156
rect 14530 18122 14564 18156
rect 14620 18122 14654 18156
rect 14710 18122 14744 18156
rect 14800 18122 14834 18156
rect 14890 18122 14924 18156
rect 14350 18032 14384 18066
rect 14440 18032 14474 18066
rect 14530 18032 14564 18066
rect 14620 18032 14654 18066
rect 14710 18032 14744 18066
rect 14800 18032 14834 18066
rect 14890 18032 14924 18066
rect 14350 17942 14384 17976
rect 14440 17942 14474 17976
rect 14530 17942 14564 17976
rect 14620 17942 14654 17976
rect 14710 17942 14744 17976
rect 14800 17942 14834 17976
rect 14890 17942 14924 17976
rect 14350 17852 14384 17886
rect 14440 17852 14474 17886
rect 14530 17852 14564 17886
rect 14620 17852 14654 17886
rect 14710 17852 14744 17886
rect 14800 17852 14834 17886
rect 14890 17852 14924 17886
rect 11630 17032 11664 17066
rect 11720 17032 11754 17066
rect 11810 17032 11844 17066
rect 11900 17032 11934 17066
rect 11990 17032 12024 17066
rect 12080 17032 12114 17066
rect 12170 17032 12204 17066
rect 11630 16942 11664 16976
rect 11720 16942 11754 16976
rect 11810 16942 11844 16976
rect 11900 16942 11934 16976
rect 11990 16942 12024 16976
rect 12080 16942 12114 16976
rect 12170 16942 12204 16976
rect 11630 16852 11664 16886
rect 11720 16852 11754 16886
rect 11810 16852 11844 16886
rect 11900 16852 11934 16886
rect 11990 16852 12024 16886
rect 12080 16852 12114 16886
rect 12170 16852 12204 16886
rect 11630 16762 11664 16796
rect 11720 16762 11754 16796
rect 11810 16762 11844 16796
rect 11900 16762 11934 16796
rect 11990 16762 12024 16796
rect 12080 16762 12114 16796
rect 12170 16762 12204 16796
rect 11630 16672 11664 16706
rect 11720 16672 11754 16706
rect 11810 16672 11844 16706
rect 11900 16672 11934 16706
rect 11990 16672 12024 16706
rect 12080 16672 12114 16706
rect 12170 16672 12204 16706
rect 11630 16582 11664 16616
rect 11720 16582 11754 16616
rect 11810 16582 11844 16616
rect 11900 16582 11934 16616
rect 11990 16582 12024 16616
rect 12080 16582 12114 16616
rect 12170 16582 12204 16616
rect 11630 16492 11664 16526
rect 11720 16492 11754 16526
rect 11810 16492 11844 16526
rect 11900 16492 11934 16526
rect 11990 16492 12024 16526
rect 12080 16492 12114 16526
rect 12170 16492 12204 16526
rect 12990 17032 13024 17066
rect 13080 17032 13114 17066
rect 13170 17032 13204 17066
rect 13260 17032 13294 17066
rect 13350 17032 13384 17066
rect 13440 17032 13474 17066
rect 13530 17032 13564 17066
rect 12990 16942 13024 16976
rect 13080 16942 13114 16976
rect 13170 16942 13204 16976
rect 13260 16942 13294 16976
rect 13350 16942 13384 16976
rect 13440 16942 13474 16976
rect 13530 16942 13564 16976
rect 12990 16852 13024 16886
rect 13080 16852 13114 16886
rect 13170 16852 13204 16886
rect 13260 16852 13294 16886
rect 13350 16852 13384 16886
rect 13440 16852 13474 16886
rect 13530 16852 13564 16886
rect 12990 16762 13024 16796
rect 13080 16762 13114 16796
rect 13170 16762 13204 16796
rect 13260 16762 13294 16796
rect 13350 16762 13384 16796
rect 13440 16762 13474 16796
rect 13530 16762 13564 16796
rect 12990 16672 13024 16706
rect 13080 16672 13114 16706
rect 13170 16672 13204 16706
rect 13260 16672 13294 16706
rect 13350 16672 13384 16706
rect 13440 16672 13474 16706
rect 13530 16672 13564 16706
rect 12990 16582 13024 16616
rect 13080 16582 13114 16616
rect 13170 16582 13204 16616
rect 13260 16582 13294 16616
rect 13350 16582 13384 16616
rect 13440 16582 13474 16616
rect 13530 16582 13564 16616
rect 12990 16492 13024 16526
rect 13080 16492 13114 16526
rect 13170 16492 13204 16526
rect 13260 16492 13294 16526
rect 13350 16492 13384 16526
rect 13440 16492 13474 16526
rect 13530 16492 13564 16526
rect 14350 17032 14384 17066
rect 14440 17032 14474 17066
rect 14530 17032 14564 17066
rect 14620 17032 14654 17066
rect 14710 17032 14744 17066
rect 14800 17032 14834 17066
rect 14890 17032 14924 17066
rect 14350 16942 14384 16976
rect 14440 16942 14474 16976
rect 14530 16942 14564 16976
rect 14620 16942 14654 16976
rect 14710 16942 14744 16976
rect 14800 16942 14834 16976
rect 14890 16942 14924 16976
rect 14350 16852 14384 16886
rect 14440 16852 14474 16886
rect 14530 16852 14564 16886
rect 14620 16852 14654 16886
rect 14710 16852 14744 16886
rect 14800 16852 14834 16886
rect 14890 16852 14924 16886
rect 14350 16762 14384 16796
rect 14440 16762 14474 16796
rect 14530 16762 14564 16796
rect 14620 16762 14654 16796
rect 14710 16762 14744 16796
rect 14800 16762 14834 16796
rect 14890 16762 14924 16796
rect 14350 16672 14384 16706
rect 14440 16672 14474 16706
rect 14530 16672 14564 16706
rect 14620 16672 14654 16706
rect 14710 16672 14744 16706
rect 14800 16672 14834 16706
rect 14890 16672 14924 16706
rect 14350 16582 14384 16616
rect 14440 16582 14474 16616
rect 14530 16582 14564 16616
rect 14620 16582 14654 16616
rect 14710 16582 14744 16616
rect 14800 16582 14834 16616
rect 14890 16582 14924 16616
rect 14350 16492 14384 16526
rect 14440 16492 14474 16526
rect 14530 16492 14564 16526
rect 14620 16492 14654 16526
rect 14710 16492 14744 16526
rect 14800 16492 14834 16526
rect 14890 16492 14924 16526
rect 11630 15672 11664 15706
rect 11720 15672 11754 15706
rect 11810 15672 11844 15706
rect 11900 15672 11934 15706
rect 11990 15672 12024 15706
rect 12080 15672 12114 15706
rect 12170 15672 12204 15706
rect 11630 15582 11664 15616
rect 11720 15582 11754 15616
rect 11810 15582 11844 15616
rect 11900 15582 11934 15616
rect 11990 15582 12024 15616
rect 12080 15582 12114 15616
rect 12170 15582 12204 15616
rect 11630 15492 11664 15526
rect 11720 15492 11754 15526
rect 11810 15492 11844 15526
rect 11900 15492 11934 15526
rect 11990 15492 12024 15526
rect 12080 15492 12114 15526
rect 12170 15492 12204 15526
rect 11630 15402 11664 15436
rect 11720 15402 11754 15436
rect 11810 15402 11844 15436
rect 11900 15402 11934 15436
rect 11990 15402 12024 15436
rect 12080 15402 12114 15436
rect 12170 15402 12204 15436
rect 11630 15312 11664 15346
rect 11720 15312 11754 15346
rect 11810 15312 11844 15346
rect 11900 15312 11934 15346
rect 11990 15312 12024 15346
rect 12080 15312 12114 15346
rect 12170 15312 12204 15346
rect 11630 15222 11664 15256
rect 11720 15222 11754 15256
rect 11810 15222 11844 15256
rect 11900 15222 11934 15256
rect 11990 15222 12024 15256
rect 12080 15222 12114 15256
rect 12170 15222 12204 15256
rect 11630 15132 11664 15166
rect 11720 15132 11754 15166
rect 11810 15132 11844 15166
rect 11900 15132 11934 15166
rect 11990 15132 12024 15166
rect 12080 15132 12114 15166
rect 12170 15132 12204 15166
rect 12990 15672 13024 15706
rect 13080 15672 13114 15706
rect 13170 15672 13204 15706
rect 13260 15672 13294 15706
rect 13350 15672 13384 15706
rect 13440 15672 13474 15706
rect 13530 15672 13564 15706
rect 12990 15582 13024 15616
rect 13080 15582 13114 15616
rect 13170 15582 13204 15616
rect 13260 15582 13294 15616
rect 13350 15582 13384 15616
rect 13440 15582 13474 15616
rect 13530 15582 13564 15616
rect 12990 15492 13024 15526
rect 13080 15492 13114 15526
rect 13170 15492 13204 15526
rect 13260 15492 13294 15526
rect 13350 15492 13384 15526
rect 13440 15492 13474 15526
rect 13530 15492 13564 15526
rect 12990 15402 13024 15436
rect 13080 15402 13114 15436
rect 13170 15402 13204 15436
rect 13260 15402 13294 15436
rect 13350 15402 13384 15436
rect 13440 15402 13474 15436
rect 13530 15402 13564 15436
rect 12990 15312 13024 15346
rect 13080 15312 13114 15346
rect 13170 15312 13204 15346
rect 13260 15312 13294 15346
rect 13350 15312 13384 15346
rect 13440 15312 13474 15346
rect 13530 15312 13564 15346
rect 12990 15222 13024 15256
rect 13080 15222 13114 15256
rect 13170 15222 13204 15256
rect 13260 15222 13294 15256
rect 13350 15222 13384 15256
rect 13440 15222 13474 15256
rect 13530 15222 13564 15256
rect 12990 15132 13024 15166
rect 13080 15132 13114 15166
rect 13170 15132 13204 15166
rect 13260 15132 13294 15166
rect 13350 15132 13384 15166
rect 13440 15132 13474 15166
rect 13530 15132 13564 15166
rect 14350 15672 14384 15706
rect 14440 15672 14474 15706
rect 14530 15672 14564 15706
rect 14620 15672 14654 15706
rect 14710 15672 14744 15706
rect 14800 15672 14834 15706
rect 14890 15672 14924 15706
rect 14350 15582 14384 15616
rect 14440 15582 14474 15616
rect 14530 15582 14564 15616
rect 14620 15582 14654 15616
rect 14710 15582 14744 15616
rect 14800 15582 14834 15616
rect 14890 15582 14924 15616
rect 14350 15492 14384 15526
rect 14440 15492 14474 15526
rect 14530 15492 14564 15526
rect 14620 15492 14654 15526
rect 14710 15492 14744 15526
rect 14800 15492 14834 15526
rect 14890 15492 14924 15526
rect 14350 15402 14384 15436
rect 14440 15402 14474 15436
rect 14530 15402 14564 15436
rect 14620 15402 14654 15436
rect 14710 15402 14744 15436
rect 14800 15402 14834 15436
rect 14890 15402 14924 15436
rect 14350 15312 14384 15346
rect 14440 15312 14474 15346
rect 14530 15312 14564 15346
rect 14620 15312 14654 15346
rect 14710 15312 14744 15346
rect 14800 15312 14834 15346
rect 14890 15312 14924 15346
rect 14350 15222 14384 15256
rect 14440 15222 14474 15256
rect 14530 15222 14564 15256
rect 14620 15222 14654 15256
rect 14710 15222 14744 15256
rect 14800 15222 14834 15256
rect 14890 15222 14924 15256
rect 14350 15132 14384 15166
rect 14440 15132 14474 15166
rect 14530 15132 14564 15166
rect 14620 15132 14654 15166
rect 14710 15132 14744 15166
rect 14800 15132 14834 15166
rect 14890 15132 14924 15166
rect 19538 12620 19578 12660
rect 19538 12520 19578 12560
rect 19538 12420 19578 12460
rect 19538 12320 19578 12360
rect 19538 12220 19578 12260
rect 19738 12620 19778 12660
rect 19738 12520 19778 12560
rect 19738 12420 19778 12460
rect 19738 12320 19778 12360
rect 19738 12220 19778 12260
rect 19938 12620 19978 12660
rect 19938 12520 19978 12560
rect 19938 12420 19978 12460
rect 19938 12320 19978 12360
rect 19938 12220 19978 12260
rect 20138 12620 20178 12660
rect 20138 12520 20178 12560
rect 20138 12420 20178 12460
rect 20138 12320 20178 12360
rect 20138 12220 20178 12260
rect 20338 12620 20378 12660
rect 20338 12520 20378 12560
rect 20338 12420 20378 12460
rect 20338 12320 20378 12360
rect 20338 12220 20378 12260
rect 20538 12620 20578 12660
rect 20538 12520 20578 12560
rect 20538 12420 20578 12460
rect 20538 12320 20578 12360
rect 20538 12220 20578 12260
rect 20738 12620 20778 12660
rect 20738 12520 20778 12560
rect 20738 12420 20778 12460
rect 20738 12320 20778 12360
rect 20738 12220 20778 12260
rect 20938 12620 20978 12660
rect 20938 12520 20978 12560
rect 20938 12420 20978 12460
rect 20938 12320 20978 12360
rect 20938 12220 20978 12260
rect 21138 12620 21178 12660
rect 21138 12520 21178 12560
rect 21138 12420 21178 12460
rect 21138 12320 21178 12360
rect 21138 12220 21178 12260
rect 21338 12620 21378 12660
rect 21338 12520 21378 12560
rect 21338 12420 21378 12460
rect 21338 12320 21378 12360
rect 21338 12220 21378 12260
rect 21538 12620 21578 12660
rect 21538 12520 21578 12560
rect 21538 12420 21578 12460
rect 21538 12320 21578 12360
rect 21538 12220 21578 12260
rect 10538 11750 10578 11790
rect 10538 11650 10578 11690
rect 10658 11750 10698 11790
rect 10658 11650 10698 11690
rect 10778 11750 10818 11790
rect 10778 11650 10818 11690
rect 10898 11750 10938 11790
rect 10898 11650 10938 11690
rect 11018 11750 11058 11790
rect 11018 11650 11058 11690
rect 11138 11750 11178 11790
rect 11138 11650 11178 11690
rect 11258 11750 11298 11790
rect 11258 11650 11298 11690
rect 11378 11750 11418 11790
rect 11378 11650 11418 11690
rect 11498 11750 11538 11790
rect 11498 11650 11538 11690
rect 11618 11750 11658 11790
rect 11618 11650 11658 11690
rect 11738 11750 11778 11790
rect 11738 11650 11778 11690
rect 11858 11750 11898 11790
rect 11858 11650 11898 11690
rect 11978 11750 12018 11790
rect 11978 11650 12018 11690
rect 12098 11750 12138 11790
rect 12098 11650 12138 11690
rect 12218 11750 12258 11790
rect 12218 11650 12258 11690
rect 12338 11750 12378 11790
rect 12338 11650 12378 11690
rect 12458 11750 12498 11790
rect 12458 11650 12498 11690
rect 12578 11750 12618 11790
rect 12578 11650 12618 11690
rect 12698 11750 12738 11790
rect 12698 11650 12738 11690
rect 12818 11750 12858 11790
rect 12818 11650 12858 11690
rect 12938 11750 12978 11790
rect 12938 11650 12978 11690
rect 13578 11750 13618 11790
rect 13578 11650 13618 11690
rect 13698 11750 13738 11790
rect 13698 11650 13738 11690
rect 13818 11750 13858 11790
rect 13818 11650 13858 11690
rect 13938 11750 13978 11790
rect 13938 11650 13978 11690
rect 14058 11750 14098 11790
rect 14058 11650 14098 11690
rect 14178 11750 14218 11790
rect 14178 11650 14218 11690
rect 14298 11750 14338 11790
rect 14298 11650 14338 11690
rect 14418 11750 14458 11790
rect 14418 11650 14458 11690
rect 14538 11750 14578 11790
rect 14538 11650 14578 11690
rect 14658 11750 14698 11790
rect 14658 11650 14698 11690
rect 14778 11750 14818 11790
rect 14778 11650 14818 11690
rect 14898 11750 14938 11790
rect 14898 11650 14938 11690
rect 15018 11750 15058 11790
rect 15018 11650 15058 11690
rect 15138 11750 15178 11790
rect 15138 11650 15178 11690
rect 15258 11750 15298 11790
rect 15258 11650 15298 11690
rect 15378 11750 15418 11790
rect 15378 11650 15418 11690
rect 15498 11750 15538 11790
rect 15498 11650 15538 11690
rect 15618 11750 15658 11790
rect 15618 11650 15658 11690
rect 15738 11750 15778 11790
rect 15738 11650 15778 11690
rect 15858 11750 15898 11790
rect 15858 11650 15898 11690
rect 15978 11750 16018 11790
rect 15978 11650 16018 11690
rect 19468 11670 19508 11710
rect 19468 11570 19508 11610
rect 19598 11670 19638 11710
rect 19598 11570 19638 11610
rect 19728 11670 19768 11710
rect 19728 11570 19768 11610
rect 19858 11670 19898 11710
rect 19858 11570 19898 11610
rect 19988 11670 20028 11710
rect 19988 11570 20028 11610
rect 20118 11670 20158 11710
rect 20118 11570 20158 11610
rect 20248 11670 20288 11710
rect 20248 11570 20288 11610
rect 20608 11670 20648 11710
rect 20608 11570 20648 11610
rect 20738 11670 20778 11710
rect 20738 11570 20778 11610
rect 20868 11670 20908 11710
rect 20868 11570 20908 11610
rect 20998 11670 21038 11710
rect 20998 11570 21038 11610
rect 21128 11670 21168 11710
rect 21128 11570 21168 11610
rect 21258 11670 21298 11710
rect 21258 11570 21298 11610
rect 21388 11670 21428 11710
rect 21388 11570 21428 11610
rect 21748 11670 21788 11710
rect 21748 11570 21788 11610
rect 21878 11670 21918 11710
rect 21878 11570 21918 11610
rect 22008 11670 22048 11710
rect 22008 11570 22048 11610
rect 22138 11670 22178 11710
rect 22138 11570 22178 11610
rect 22268 11670 22308 11710
rect 22268 11570 22308 11610
rect 22398 11670 22438 11710
rect 22398 11570 22438 11610
rect 22528 11670 22568 11710
rect 22528 11570 22568 11610
rect 11638 10590 11678 10630
rect 11638 10490 11678 10530
rect 11638 10390 11678 10430
rect 11638 10290 11678 10330
rect 11638 10190 11678 10230
rect 11638 10090 11678 10130
rect 11818 10590 11858 10630
rect 11818 10490 11858 10530
rect 11818 10390 11858 10430
rect 11818 10290 11858 10330
rect 11818 10190 11858 10230
rect 11818 10090 11858 10130
rect 11998 10590 12038 10630
rect 11998 10490 12038 10530
rect 11998 10390 12038 10430
rect 11998 10290 12038 10330
rect 11998 10190 12038 10230
rect 11998 10090 12038 10130
rect 12178 10590 12218 10630
rect 12178 10490 12218 10530
rect 12178 10390 12218 10430
rect 12178 10290 12218 10330
rect 12178 10190 12218 10230
rect 12178 10090 12218 10130
rect 12358 10590 12398 10630
rect 12358 10490 12398 10530
rect 12358 10390 12398 10430
rect 12358 10290 12398 10330
rect 12358 10190 12398 10230
rect 12358 10090 12398 10130
rect 12538 10590 12578 10630
rect 12538 10490 12578 10530
rect 12538 10390 12578 10430
rect 12538 10290 12578 10330
rect 12538 10190 12578 10230
rect 12538 10090 12578 10130
rect 12718 10590 12758 10630
rect 12718 10490 12758 10530
rect 12718 10390 12758 10430
rect 12718 10290 12758 10330
rect 12718 10190 12758 10230
rect 12718 10090 12758 10130
rect 12898 10590 12938 10630
rect 12898 10490 12938 10530
rect 12898 10390 12938 10430
rect 12898 10290 12938 10330
rect 12898 10190 12938 10230
rect 12898 10090 12938 10130
rect 13078 10590 13118 10630
rect 13078 10490 13118 10530
rect 13078 10390 13118 10430
rect 13078 10290 13118 10330
rect 13078 10190 13118 10230
rect 13078 10090 13118 10130
rect 13258 10590 13298 10630
rect 13258 10490 13298 10530
rect 13258 10390 13298 10430
rect 13258 10290 13298 10330
rect 13258 10190 13298 10230
rect 13258 10090 13298 10130
rect 13438 10590 13478 10630
rect 13438 10490 13478 10530
rect 13438 10390 13478 10430
rect 13438 10290 13478 10330
rect 13438 10190 13478 10230
rect 13438 10090 13478 10130
rect 13618 10590 13658 10630
rect 13618 10490 13658 10530
rect 13618 10390 13658 10430
rect 13618 10290 13658 10330
rect 13618 10190 13658 10230
rect 13618 10090 13658 10130
rect 13798 10590 13838 10630
rect 13798 10490 13838 10530
rect 13798 10390 13838 10430
rect 13798 10290 13838 10330
rect 13798 10190 13838 10230
rect 13798 10090 13838 10130
rect 13978 10590 14018 10630
rect 13978 10490 14018 10530
rect 13978 10390 14018 10430
rect 13978 10290 14018 10330
rect 13978 10190 14018 10230
rect 13978 10090 14018 10130
rect 14158 10590 14198 10630
rect 14158 10490 14198 10530
rect 14158 10390 14198 10430
rect 14158 10290 14198 10330
rect 14158 10190 14198 10230
rect 14158 10090 14198 10130
rect 14338 10590 14378 10630
rect 14338 10490 14378 10530
rect 14338 10390 14378 10430
rect 14338 10290 14378 10330
rect 14338 10190 14378 10230
rect 14338 10090 14378 10130
rect 14518 10590 14558 10630
rect 14518 10490 14558 10530
rect 14518 10390 14558 10430
rect 14518 10290 14558 10330
rect 14518 10190 14558 10230
rect 14518 10090 14558 10130
rect 14698 10590 14738 10630
rect 14698 10490 14738 10530
rect 14698 10390 14738 10430
rect 14698 10290 14738 10330
rect 14698 10190 14738 10230
rect 14698 10090 14738 10130
rect 14878 10590 14918 10630
rect 14878 10490 14918 10530
rect 14878 10390 14918 10430
rect 14878 10290 14918 10330
rect 15508 10390 15548 10430
rect 15508 10290 15548 10330
rect 15618 10390 15658 10430
rect 15618 10290 15658 10330
rect 15728 10390 15768 10430
rect 15728 10290 15768 10330
rect 15838 10390 15878 10430
rect 15838 10290 15878 10330
rect 15948 10390 15988 10430
rect 15948 10290 15988 10330
rect 14878 10190 14918 10230
rect 14878 10090 14918 10130
rect 11648 9590 11688 9630
rect 11648 9490 11688 9530
rect 11758 9590 11798 9630
rect 11758 9490 11798 9530
rect 11868 9590 11908 9630
rect 11868 9490 11908 9530
rect 11978 9590 12018 9630
rect 11978 9490 12018 9530
rect 12088 9590 12128 9630
rect 12088 9490 12128 9530
rect 12198 9590 12238 9630
rect 12198 9490 12238 9530
rect 12308 9590 12348 9630
rect 12308 9490 12348 9530
rect 12418 9590 12458 9630
rect 12418 9490 12458 9530
rect 12528 9590 12568 9630
rect 12528 9490 12568 9530
rect 12638 9590 12678 9630
rect 12638 9490 12678 9530
rect 12748 9590 12788 9630
rect 12748 9490 12788 9530
rect 12858 9590 12898 9630
rect 12858 9490 12898 9530
rect 12968 9590 13008 9630
rect 12968 9490 13008 9530
rect 13548 9590 13588 9630
rect 13548 9490 13588 9530
rect 13658 9590 13698 9630
rect 13658 9490 13698 9530
rect 13768 9590 13808 9630
rect 13768 9490 13808 9530
rect 13878 9590 13918 9630
rect 13878 9490 13918 9530
rect 13988 9590 14028 9630
rect 13988 9490 14028 9530
rect 14098 9590 14138 9630
rect 14098 9490 14138 9530
rect 14208 9590 14248 9630
rect 14208 9490 14248 9530
rect 14318 9590 14358 9630
rect 14318 9490 14358 9530
rect 14428 9590 14468 9630
rect 14428 9490 14468 9530
rect 14538 9590 14578 9630
rect 14538 9490 14578 9530
rect 14648 9590 14688 9630
rect 14648 9490 14688 9530
rect 14758 9590 14798 9630
rect 14758 9490 14798 9530
rect 14868 9590 14908 9630
rect 14868 9490 14908 9530
rect 13268 7600 13308 7640
rect 13268 7500 13308 7540
rect 13268 7400 13308 7440
rect 13268 7300 13308 7340
rect 13378 7600 13418 7640
rect 13378 7500 13418 7540
rect 13378 7400 13418 7440
rect 13378 7300 13418 7340
rect 13488 7600 13528 7640
rect 13488 7500 13528 7540
rect 13488 7400 13528 7440
rect 13488 7300 13528 7340
rect 13788 7600 13828 7640
rect 13788 7500 13828 7540
rect 13788 7400 13828 7440
rect 13788 7300 13828 7340
rect 13898 7600 13938 7640
rect 13898 7500 13938 7540
rect 13898 7400 13938 7440
rect 13898 7300 13938 7340
rect 14008 7600 14048 7640
rect 14168 7600 14208 7640
rect 14008 7500 14048 7540
rect 14168 7500 14208 7540
rect 14008 7400 14048 7440
rect 14168 7400 14208 7440
rect 14008 7300 14048 7340
rect 14168 7300 14208 7340
rect 14278 7600 14318 7640
rect 14278 7500 14318 7540
rect 14278 7400 14318 7440
rect 14278 7300 14318 7340
rect 14388 7600 14428 7640
rect 14388 7500 14428 7540
rect 14388 7400 14428 7440
rect 14388 7300 14428 7340
rect 14688 7600 14728 7640
rect 14688 7500 14728 7540
rect 14688 7400 14728 7440
rect 14688 7300 14728 7340
rect 14798 7600 14838 7640
rect 14798 7500 14838 7540
rect 14798 7400 14838 7440
rect 14798 7300 14838 7340
rect 14908 7600 14948 7640
rect 14908 7500 14948 7540
rect 14908 7400 14948 7440
rect 14908 7300 14948 7340
rect 15198 7600 15238 7640
rect 15198 7500 15238 7540
rect 15198 7400 15238 7440
rect 15198 7300 15238 7340
rect 15308 7600 15348 7640
rect 15308 7500 15348 7540
rect 15308 7400 15348 7440
rect 15308 7300 15348 7340
rect 15528 7600 15568 7640
rect 15528 7500 15568 7540
rect 15528 7400 15568 7440
rect 15528 7300 15568 7340
rect 15638 7600 15678 7640
rect 15638 7500 15678 7540
rect 15638 7400 15678 7440
rect 15638 7300 15678 7340
rect 15858 7600 15898 7640
rect 15858 7500 15898 7540
rect 15858 7400 15898 7440
rect 15858 7300 15898 7340
rect 15968 7600 16008 7640
rect 15968 7500 16008 7540
rect 15968 7400 16008 7440
rect 15968 7300 16008 7340
rect 16408 7600 16448 7640
rect 16408 7500 16448 7540
rect 16408 7400 16448 7440
rect 16408 7300 16448 7340
rect 16538 7600 16578 7640
rect 16538 7500 16578 7540
rect 16538 7400 16578 7440
rect 16538 7300 16578 7340
rect 16798 7600 16838 7640
rect 16798 7500 16838 7540
rect 16798 7400 16838 7440
rect 16798 7300 16838 7340
rect 16928 7600 16968 7640
rect 16928 7500 16968 7540
rect 16928 7400 16968 7440
rect 16928 7300 16968 7340
rect 17188 7600 17228 7640
rect 17188 7500 17228 7540
rect 17188 7400 17228 7440
rect 17188 7300 17228 7340
rect 17318 7600 17358 7640
rect 17318 7500 17358 7540
rect 17318 7400 17358 7440
rect 17318 7300 17358 7340
rect 17478 7600 17518 7640
rect 17478 7500 17518 7540
rect 17478 7400 17518 7440
rect 17478 7300 17518 7340
rect 17608 7600 17648 7640
rect 17608 7500 17648 7540
rect 17608 7400 17648 7440
rect 17608 7300 17648 7340
rect 13268 6840 13308 6880
rect 13268 6740 13308 6780
rect 13268 6640 13308 6680
rect 13268 6540 13308 6580
rect 13378 6840 13418 6880
rect 13378 6740 13418 6780
rect 13378 6640 13418 6680
rect 13378 6540 13418 6580
rect 13488 6840 13528 6880
rect 13488 6740 13528 6780
rect 13488 6640 13528 6680
rect 13488 6540 13528 6580
rect 13788 6840 13828 6880
rect 13788 6740 13828 6780
rect 13788 6640 13828 6680
rect 13788 6540 13828 6580
rect 13898 6840 13938 6880
rect 13898 6740 13938 6780
rect 13898 6640 13938 6680
rect 13898 6540 13938 6580
rect 14008 6840 14048 6880
rect 14168 6840 14208 6880
rect 14008 6740 14048 6780
rect 14168 6740 14208 6780
rect 14008 6640 14048 6680
rect 14168 6640 14208 6680
rect 14008 6540 14048 6580
rect 14168 6540 14208 6580
rect 14278 6840 14318 6880
rect 14278 6740 14318 6780
rect 14278 6640 14318 6680
rect 14278 6540 14318 6580
rect 14388 6840 14428 6880
rect 14388 6740 14428 6780
rect 14388 6640 14428 6680
rect 14388 6540 14428 6580
rect 14688 6840 14728 6880
rect 14688 6740 14728 6780
rect 14688 6640 14728 6680
rect 14688 6540 14728 6580
rect 14798 6840 14838 6880
rect 14798 6740 14838 6780
rect 14798 6640 14838 6680
rect 14798 6540 14838 6580
rect 14908 6840 14948 6880
rect 14908 6740 14948 6780
rect 14908 6640 14948 6680
rect 14908 6540 14948 6580
rect 15208 6840 15248 6880
rect 15208 6740 15248 6780
rect 15208 6640 15248 6680
rect 15208 6540 15248 6580
rect 15318 6840 15358 6880
rect 15318 6740 15358 6780
rect 15318 6640 15358 6680
rect 15318 6540 15358 6580
rect 15428 6840 15468 6880
rect 15428 6740 15468 6780
rect 15428 6640 15468 6680
rect 15428 6540 15468 6580
rect 15648 6840 15688 6880
rect 15648 6740 15688 6780
rect 15648 6640 15688 6680
rect 15648 6540 15688 6580
rect 15758 6840 15798 6880
rect 15758 6740 15798 6780
rect 15758 6640 15798 6680
rect 15758 6540 15798 6580
rect 15978 6840 16018 6880
rect 15978 6740 16018 6780
rect 15978 6640 16018 6680
rect 15978 6540 16018 6580
rect 16088 6840 16128 6880
rect 16088 6740 16128 6780
rect 16088 6640 16128 6680
rect 16088 6540 16128 6580
rect 16408 6840 16448 6880
rect 16408 6740 16448 6780
rect 16408 6640 16448 6680
rect 16408 6540 16448 6580
rect 16538 6840 16578 6880
rect 16538 6740 16578 6780
rect 16538 6640 16578 6680
rect 16538 6540 16578 6580
rect 16798 6840 16838 6880
rect 16798 6740 16838 6780
rect 16798 6640 16838 6680
rect 16798 6540 16838 6580
rect 16928 6840 16968 6880
rect 16928 6740 16968 6780
rect 16928 6640 16968 6680
rect 16928 6540 16968 6580
rect 17188 6840 17228 6880
rect 17188 6740 17228 6780
rect 17188 6640 17228 6680
rect 17188 6540 17228 6580
rect 17318 6840 17358 6880
rect 17318 6740 17358 6780
rect 17318 6640 17358 6680
rect 17318 6540 17358 6580
rect 17478 6840 17518 6880
rect 17478 6740 17518 6780
rect 17478 6640 17518 6680
rect 17478 6540 17518 6580
rect 17608 6840 17648 6880
rect 17608 6740 17648 6780
rect 17608 6640 17648 6680
rect 17608 6540 17648 6580
rect 17868 6840 17908 6880
rect 17868 6740 17908 6780
rect 17868 6640 17908 6680
rect 17868 6540 17908 6580
rect 17998 6840 18038 6880
rect 17998 6740 18038 6780
rect 17998 6640 18038 6680
rect 17998 6540 18038 6580
rect 19558 6870 19598 6910
rect 19558 6770 19598 6810
rect 19558 6670 19598 6710
rect 19558 6570 19598 6610
rect 19778 6870 19818 6910
rect 19778 6770 19818 6810
rect 19778 6670 19818 6710
rect 19778 6570 19818 6610
rect 19998 6870 20038 6910
rect 19998 6770 20038 6810
rect 19998 6670 20038 6710
rect 19998 6570 20038 6610
rect 20218 6870 20258 6910
rect 20218 6770 20258 6810
rect 20218 6670 20258 6710
rect 20218 6570 20258 6610
rect 20438 6870 20478 6910
rect 20438 6770 20478 6810
rect 20438 6670 20478 6710
rect 20438 6570 20478 6610
rect 20658 6870 20698 6910
rect 20658 6770 20698 6810
rect 20658 6670 20698 6710
rect 20658 6570 20698 6610
rect 20878 6870 20918 6910
rect 21078 6870 21118 6910
rect 20878 6770 20918 6810
rect 21078 6770 21118 6810
rect 20878 6670 20918 6710
rect 21078 6670 21118 6710
rect 20878 6570 20918 6610
rect 21078 6570 21118 6610
rect 21298 6870 21338 6910
rect 21298 6770 21338 6810
rect 21298 6670 21338 6710
rect 21298 6570 21338 6610
rect 21518 6870 21558 6910
rect 21518 6770 21558 6810
rect 21518 6670 21558 6710
rect 21518 6570 21558 6610
rect 21738 6870 21778 6910
rect 21738 6770 21778 6810
rect 21738 6670 21778 6710
rect 21738 6570 21778 6610
rect 21958 6870 21998 6910
rect 21958 6770 21998 6810
rect 21958 6670 21998 6710
rect 21958 6570 21998 6610
rect 22178 6870 22218 6910
rect 22178 6770 22218 6810
rect 22178 6670 22218 6710
rect 22178 6570 22218 6610
rect 22398 6870 22438 6910
rect 22398 6770 22438 6810
rect 22398 6670 22438 6710
rect 22398 6570 22438 6610
rect 23218 5360 23258 5400
rect 23218 5260 23258 5300
rect 23218 5160 23258 5200
rect 23218 5060 23258 5100
rect 23598 5360 23638 5400
rect 23598 5260 23638 5300
rect 23598 5160 23638 5200
rect 23598 5060 23638 5100
rect 23738 5360 23778 5400
rect 23738 5260 23778 5300
rect 23738 5160 23778 5200
rect 23738 5060 23778 5100
rect 24118 5360 24158 5400
rect 24118 5260 24158 5300
rect 24118 5160 24158 5200
rect 24118 5060 24158 5100
rect 24258 5360 24298 5400
rect 24258 5260 24298 5300
rect 24258 5160 24298 5200
rect 24258 5060 24298 5100
rect 24638 5360 24678 5400
rect 24638 5260 24678 5300
rect 24638 5160 24678 5200
rect 24638 5060 24678 5100
rect 24778 5360 24818 5400
rect 24778 5260 24818 5300
rect 24778 5160 24818 5200
rect 24778 5060 24818 5100
rect 25158 5360 25198 5400
rect 25158 5260 25198 5300
rect 25158 5160 25198 5200
rect 25158 5060 25198 5100
rect 12608 3460 12648 3500
rect 12718 3460 12758 3500
rect 13028 3460 13068 3500
rect 13138 3460 13178 3500
rect 13248 3460 13288 3500
rect 13698 3460 13738 3500
rect 13808 3460 13848 3500
rect 13918 3460 13958 3500
rect 14138 3460 14178 3500
rect 14248 3460 14288 3500
rect 14358 3460 14398 3500
rect 14468 3460 14508 3500
rect 14978 3460 15018 3500
rect 15088 3460 15128 3500
rect 15398 3460 15438 3500
rect 15508 3460 15548 3500
rect 15618 3460 15658 3500
rect 15848 3460 15888 3500
rect 15958 3460 15998 3500
rect 16068 3460 16108 3500
rect 16208 3460 16248 3500
rect 16318 3460 16358 3500
rect 16428 3460 16468 3500
rect 16788 3460 16828 3500
rect 16898 3460 16938 3500
rect 17008 3460 17048 3500
rect 17228 3460 17268 3500
rect 17338 3460 17378 3500
rect 17448 3460 17488 3500
rect 17848 3460 17888 3500
rect 17958 3460 17998 3500
rect 18188 3460 18228 3500
rect 18298 3460 18338 3500
rect 18408 3460 18448 3500
rect 18548 3460 18588 3500
rect 18658 3460 18698 3500
rect 18768 3460 18808 3500
rect 19148 3460 19188 3500
rect 19258 3460 19298 3500
rect 19488 3460 19528 3500
rect 19598 3460 19638 3500
rect 19708 3460 19748 3500
rect 19848 3460 19888 3500
rect 19958 3460 19998 3500
rect 20068 3460 20108 3500
rect 20448 3460 20488 3500
rect 20558 3460 20598 3500
rect 20788 3460 20828 3500
rect 20898 3460 20938 3500
rect 21008 3460 21048 3500
rect 21148 3460 21188 3500
rect 21258 3460 21298 3500
rect 21368 3460 21408 3500
rect 21748 3460 21788 3500
rect 21858 3460 21898 3500
rect 22088 3460 22128 3500
rect 22198 3460 22238 3500
rect 22308 3460 22348 3500
rect 22448 3460 22488 3500
rect 22558 3460 22598 3500
rect 22668 3460 22708 3500
rect 23218 4670 23258 4710
rect 23218 4570 23258 4610
rect 23218 4470 23258 4510
rect 23218 4370 23258 4410
rect 23218 4270 23258 4310
rect 23218 4170 23258 4210
rect 23328 4670 23368 4710
rect 23328 4570 23368 4610
rect 23328 4470 23368 4510
rect 23328 4370 23368 4410
rect 23328 4270 23368 4310
rect 23328 4170 23368 4210
rect 23738 4670 23778 4710
rect 23738 4570 23778 4610
rect 23738 4470 23778 4510
rect 23738 4370 23778 4410
rect 23738 4270 23778 4310
rect 23738 4170 23778 4210
rect 23848 4670 23888 4710
rect 23848 4570 23888 4610
rect 23848 4470 23888 4510
rect 23848 4370 23888 4410
rect 23848 4270 23888 4310
rect 23848 4170 23888 4210
rect 24258 4670 24298 4710
rect 24258 4570 24298 4610
rect 24258 4470 24298 4510
rect 24258 4370 24298 4410
rect 24258 4270 24298 4310
rect 24258 4170 24298 4210
rect 24368 4670 24408 4710
rect 24368 4570 24408 4610
rect 24368 4470 24408 4510
rect 24368 4370 24408 4410
rect 24368 4270 24408 4310
rect 24368 4170 24408 4210
rect 23216 3890 23256 3930
rect 23216 3790 23256 3830
rect 23216 3690 23256 3730
rect 23216 3590 23256 3630
rect 23328 3890 23368 3930
rect 23328 3790 23368 3830
rect 23328 3690 23368 3730
rect 23328 3590 23368 3630
rect 23736 3890 23776 3930
rect 23736 3790 23776 3830
rect 23736 3690 23776 3730
rect 23736 3590 23776 3630
rect 23848 3890 23888 3930
rect 23848 3790 23888 3830
rect 23848 3690 23888 3730
rect 23848 3590 23888 3630
rect 24256 3890 24296 3930
rect 24256 3790 24296 3830
rect 24256 3690 24296 3730
rect 24256 3590 24296 3630
rect 24368 3890 24408 3930
rect 24368 3790 24408 3830
rect 24368 3690 24408 3730
rect 24368 3590 24408 3630
<< psubdiff >>
rect 13228 19070 13328 19100
rect 13228 19030 13258 19070
rect 13298 19030 13328 19070
rect 13228 18990 13328 19030
rect 13228 18950 13258 18990
rect 13298 18950 13328 18990
rect 13228 18910 13328 18950
rect 13228 18870 13258 18910
rect 13298 18870 13328 18910
rect 13228 18840 13328 18870
rect 11274 18752 12562 18784
rect 11274 18718 11408 18752
rect 11442 18718 11498 18752
rect 11532 18718 11588 18752
rect 11622 18718 11678 18752
rect 11712 18718 11768 18752
rect 11802 18718 11858 18752
rect 11892 18718 11948 18752
rect 11982 18718 12038 18752
rect 12072 18718 12128 18752
rect 12162 18718 12218 18752
rect 12252 18718 12308 18752
rect 12342 18718 12398 18752
rect 12432 18718 12562 18752
rect 11274 18683 12562 18718
rect 11274 18668 11375 18683
rect 11274 18634 11307 18668
rect 11341 18634 11375 18668
rect 11274 18578 11375 18634
rect 12461 18668 12562 18683
rect 12461 18634 12494 18668
rect 12528 18634 12562 18668
rect 11274 18544 11307 18578
rect 11341 18544 11375 18578
rect 11274 18488 11375 18544
rect 11274 18454 11307 18488
rect 11341 18454 11375 18488
rect 11274 18398 11375 18454
rect 11274 18364 11307 18398
rect 11341 18364 11375 18398
rect 11274 18308 11375 18364
rect 11274 18274 11307 18308
rect 11341 18274 11375 18308
rect 11274 18218 11375 18274
rect 11274 18184 11307 18218
rect 11341 18184 11375 18218
rect 11274 18128 11375 18184
rect 11274 18094 11307 18128
rect 11341 18094 11375 18128
rect 11274 18038 11375 18094
rect 11274 18004 11307 18038
rect 11341 18004 11375 18038
rect 11274 17948 11375 18004
rect 11274 17914 11307 17948
rect 11341 17914 11375 17948
rect 11274 17858 11375 17914
rect 11274 17824 11307 17858
rect 11341 17824 11375 17858
rect 11274 17768 11375 17824
rect 11274 17734 11307 17768
rect 11341 17734 11375 17768
rect 11274 17678 11375 17734
rect 11274 17644 11307 17678
rect 11341 17644 11375 17678
rect 12461 18578 12562 18634
rect 12461 18544 12494 18578
rect 12528 18544 12562 18578
rect 12461 18488 12562 18544
rect 12461 18454 12494 18488
rect 12528 18454 12562 18488
rect 12461 18398 12562 18454
rect 12461 18364 12494 18398
rect 12528 18364 12562 18398
rect 12461 18308 12562 18364
rect 12461 18274 12494 18308
rect 12528 18274 12562 18308
rect 12461 18218 12562 18274
rect 12461 18184 12494 18218
rect 12528 18184 12562 18218
rect 12461 18128 12562 18184
rect 12461 18094 12494 18128
rect 12528 18094 12562 18128
rect 12461 18038 12562 18094
rect 12461 18004 12494 18038
rect 12528 18004 12562 18038
rect 12461 17948 12562 18004
rect 12461 17914 12494 17948
rect 12528 17914 12562 17948
rect 12461 17858 12562 17914
rect 12461 17824 12494 17858
rect 12528 17824 12562 17858
rect 12461 17768 12562 17824
rect 12461 17734 12494 17768
rect 12528 17734 12562 17768
rect 12461 17678 12562 17734
rect 11274 17597 11375 17644
rect 12461 17644 12494 17678
rect 12528 17644 12562 17678
rect 12461 17597 12562 17644
rect 11274 17588 12562 17597
rect 11274 17554 11307 17588
rect 11341 17565 12494 17588
rect 11341 17554 11408 17565
rect 11274 17531 11408 17554
rect 11442 17531 11498 17565
rect 11532 17531 11588 17565
rect 11622 17531 11678 17565
rect 11712 17531 11768 17565
rect 11802 17531 11858 17565
rect 11892 17531 11948 17565
rect 11982 17531 12038 17565
rect 12072 17531 12128 17565
rect 12162 17531 12218 17565
rect 12252 17531 12308 17565
rect 12342 17531 12398 17565
rect 12432 17554 12494 17565
rect 12528 17554 12562 17588
rect 12432 17531 12562 17554
rect 11274 17496 12562 17531
rect 12634 18752 13922 18784
rect 12634 18718 12768 18752
rect 12802 18718 12858 18752
rect 12892 18718 12948 18752
rect 12982 18718 13038 18752
rect 13072 18718 13128 18752
rect 13162 18718 13218 18752
rect 13252 18718 13308 18752
rect 13342 18718 13398 18752
rect 13432 18718 13488 18752
rect 13522 18718 13578 18752
rect 13612 18718 13668 18752
rect 13702 18718 13758 18752
rect 13792 18718 13922 18752
rect 12634 18683 13922 18718
rect 12634 18668 12735 18683
rect 12634 18634 12667 18668
rect 12701 18634 12735 18668
rect 12634 18578 12735 18634
rect 13821 18668 13922 18683
rect 13821 18634 13854 18668
rect 13888 18634 13922 18668
rect 12634 18544 12667 18578
rect 12701 18544 12735 18578
rect 12634 18488 12735 18544
rect 12634 18454 12667 18488
rect 12701 18454 12735 18488
rect 12634 18398 12735 18454
rect 12634 18364 12667 18398
rect 12701 18364 12735 18398
rect 12634 18308 12735 18364
rect 12634 18274 12667 18308
rect 12701 18274 12735 18308
rect 12634 18218 12735 18274
rect 12634 18184 12667 18218
rect 12701 18184 12735 18218
rect 12634 18128 12735 18184
rect 12634 18094 12667 18128
rect 12701 18094 12735 18128
rect 12634 18038 12735 18094
rect 12634 18004 12667 18038
rect 12701 18004 12735 18038
rect 12634 17948 12735 18004
rect 12634 17914 12667 17948
rect 12701 17914 12735 17948
rect 12634 17858 12735 17914
rect 12634 17824 12667 17858
rect 12701 17824 12735 17858
rect 12634 17768 12735 17824
rect 12634 17734 12667 17768
rect 12701 17734 12735 17768
rect 12634 17678 12735 17734
rect 12634 17644 12667 17678
rect 12701 17644 12735 17678
rect 13821 18578 13922 18634
rect 13821 18544 13854 18578
rect 13888 18544 13922 18578
rect 13821 18488 13922 18544
rect 13821 18454 13854 18488
rect 13888 18454 13922 18488
rect 13821 18398 13922 18454
rect 13821 18364 13854 18398
rect 13888 18364 13922 18398
rect 13821 18308 13922 18364
rect 13821 18274 13854 18308
rect 13888 18274 13922 18308
rect 13821 18218 13922 18274
rect 13821 18184 13854 18218
rect 13888 18184 13922 18218
rect 13821 18128 13922 18184
rect 13821 18094 13854 18128
rect 13888 18094 13922 18128
rect 13821 18038 13922 18094
rect 13821 18004 13854 18038
rect 13888 18004 13922 18038
rect 13821 17948 13922 18004
rect 13821 17914 13854 17948
rect 13888 17914 13922 17948
rect 13821 17858 13922 17914
rect 13821 17824 13854 17858
rect 13888 17824 13922 17858
rect 13821 17768 13922 17824
rect 13821 17734 13854 17768
rect 13888 17734 13922 17768
rect 13821 17678 13922 17734
rect 12634 17597 12735 17644
rect 13821 17644 13854 17678
rect 13888 17644 13922 17678
rect 13821 17597 13922 17644
rect 12634 17588 13922 17597
rect 12634 17554 12667 17588
rect 12701 17565 13854 17588
rect 12701 17554 12768 17565
rect 12634 17531 12768 17554
rect 12802 17531 12858 17565
rect 12892 17531 12948 17565
rect 12982 17531 13038 17565
rect 13072 17531 13128 17565
rect 13162 17531 13218 17565
rect 13252 17531 13308 17565
rect 13342 17531 13398 17565
rect 13432 17531 13488 17565
rect 13522 17531 13578 17565
rect 13612 17531 13668 17565
rect 13702 17531 13758 17565
rect 13792 17554 13854 17565
rect 13888 17554 13922 17588
rect 13792 17531 13922 17554
rect 12634 17496 13922 17531
rect 13994 18752 15282 18784
rect 13994 18718 14128 18752
rect 14162 18718 14218 18752
rect 14252 18718 14308 18752
rect 14342 18718 14398 18752
rect 14432 18718 14488 18752
rect 14522 18718 14578 18752
rect 14612 18718 14668 18752
rect 14702 18718 14758 18752
rect 14792 18718 14848 18752
rect 14882 18718 14938 18752
rect 14972 18718 15028 18752
rect 15062 18718 15118 18752
rect 15152 18718 15282 18752
rect 13994 18683 15282 18718
rect 13994 18668 14095 18683
rect 13994 18634 14027 18668
rect 14061 18634 14095 18668
rect 13994 18578 14095 18634
rect 15181 18668 15282 18683
rect 15181 18634 15214 18668
rect 15248 18634 15282 18668
rect 13994 18544 14027 18578
rect 14061 18544 14095 18578
rect 13994 18488 14095 18544
rect 13994 18454 14027 18488
rect 14061 18454 14095 18488
rect 13994 18398 14095 18454
rect 13994 18364 14027 18398
rect 14061 18364 14095 18398
rect 13994 18308 14095 18364
rect 13994 18274 14027 18308
rect 14061 18274 14095 18308
rect 13994 18218 14095 18274
rect 13994 18184 14027 18218
rect 14061 18184 14095 18218
rect 13994 18128 14095 18184
rect 13994 18094 14027 18128
rect 14061 18094 14095 18128
rect 13994 18038 14095 18094
rect 13994 18004 14027 18038
rect 14061 18004 14095 18038
rect 13994 17948 14095 18004
rect 13994 17914 14027 17948
rect 14061 17914 14095 17948
rect 13994 17858 14095 17914
rect 13994 17824 14027 17858
rect 14061 17824 14095 17858
rect 13994 17768 14095 17824
rect 13994 17734 14027 17768
rect 14061 17734 14095 17768
rect 13994 17678 14095 17734
rect 13994 17644 14027 17678
rect 14061 17644 14095 17678
rect 15181 18578 15282 18634
rect 15181 18544 15214 18578
rect 15248 18544 15282 18578
rect 15181 18488 15282 18544
rect 15181 18454 15214 18488
rect 15248 18454 15282 18488
rect 15181 18398 15282 18454
rect 15181 18364 15214 18398
rect 15248 18364 15282 18398
rect 15181 18308 15282 18364
rect 15181 18274 15214 18308
rect 15248 18274 15282 18308
rect 15181 18218 15282 18274
rect 15181 18184 15214 18218
rect 15248 18184 15282 18218
rect 15181 18128 15282 18184
rect 15181 18094 15214 18128
rect 15248 18094 15282 18128
rect 15181 18038 15282 18094
rect 15181 18004 15214 18038
rect 15248 18004 15282 18038
rect 15181 17948 15282 18004
rect 15181 17914 15214 17948
rect 15248 17914 15282 17948
rect 15181 17858 15282 17914
rect 15181 17824 15214 17858
rect 15248 17824 15282 17858
rect 15181 17768 15282 17824
rect 15181 17734 15214 17768
rect 15248 17734 15282 17768
rect 15181 17678 15282 17734
rect 13994 17597 14095 17644
rect 15181 17644 15214 17678
rect 15248 17644 15282 17678
rect 15181 17597 15282 17644
rect 13994 17588 15282 17597
rect 13994 17554 14027 17588
rect 14061 17565 15214 17588
rect 14061 17554 14128 17565
rect 13994 17531 14128 17554
rect 14162 17531 14218 17565
rect 14252 17531 14308 17565
rect 14342 17531 14398 17565
rect 14432 17531 14488 17565
rect 14522 17531 14578 17565
rect 14612 17531 14668 17565
rect 14702 17531 14758 17565
rect 14792 17531 14848 17565
rect 14882 17531 14938 17565
rect 14972 17531 15028 17565
rect 15062 17531 15118 17565
rect 15152 17554 15214 17565
rect 15248 17554 15282 17588
rect 15152 17531 15282 17554
rect 13994 17496 15282 17531
rect 11274 17392 12562 17424
rect 11274 17358 11408 17392
rect 11442 17358 11498 17392
rect 11532 17358 11588 17392
rect 11622 17358 11678 17392
rect 11712 17358 11768 17392
rect 11802 17358 11858 17392
rect 11892 17358 11948 17392
rect 11982 17358 12038 17392
rect 12072 17358 12128 17392
rect 12162 17358 12218 17392
rect 12252 17358 12308 17392
rect 12342 17358 12398 17392
rect 12432 17358 12562 17392
rect 11274 17323 12562 17358
rect 11274 17308 11375 17323
rect 11274 17274 11307 17308
rect 11341 17274 11375 17308
rect 11274 17218 11375 17274
rect 12461 17308 12562 17323
rect 12461 17274 12494 17308
rect 12528 17274 12562 17308
rect 11274 17184 11307 17218
rect 11341 17184 11375 17218
rect 11274 17128 11375 17184
rect 11274 17094 11307 17128
rect 11341 17094 11375 17128
rect 11274 17038 11375 17094
rect 11274 17004 11307 17038
rect 11341 17004 11375 17038
rect 11274 16948 11375 17004
rect 11274 16914 11307 16948
rect 11341 16914 11375 16948
rect 11274 16858 11375 16914
rect 11274 16824 11307 16858
rect 11341 16824 11375 16858
rect 11274 16768 11375 16824
rect 11274 16734 11307 16768
rect 11341 16734 11375 16768
rect 11274 16678 11375 16734
rect 11274 16644 11307 16678
rect 11341 16644 11375 16678
rect 11274 16588 11375 16644
rect 11274 16554 11307 16588
rect 11341 16554 11375 16588
rect 11274 16498 11375 16554
rect 11274 16464 11307 16498
rect 11341 16464 11375 16498
rect 11274 16408 11375 16464
rect 11274 16374 11307 16408
rect 11341 16374 11375 16408
rect 11274 16318 11375 16374
rect 11274 16284 11307 16318
rect 11341 16284 11375 16318
rect 12461 17218 12562 17274
rect 12461 17184 12494 17218
rect 12528 17184 12562 17218
rect 12461 17128 12562 17184
rect 12461 17094 12494 17128
rect 12528 17094 12562 17128
rect 12461 17038 12562 17094
rect 12461 17004 12494 17038
rect 12528 17004 12562 17038
rect 12461 16948 12562 17004
rect 12461 16914 12494 16948
rect 12528 16914 12562 16948
rect 12461 16858 12562 16914
rect 12461 16824 12494 16858
rect 12528 16824 12562 16858
rect 12461 16768 12562 16824
rect 12461 16734 12494 16768
rect 12528 16734 12562 16768
rect 12461 16678 12562 16734
rect 12461 16644 12494 16678
rect 12528 16644 12562 16678
rect 12461 16588 12562 16644
rect 12461 16554 12494 16588
rect 12528 16554 12562 16588
rect 12461 16498 12562 16554
rect 12461 16464 12494 16498
rect 12528 16464 12562 16498
rect 12461 16408 12562 16464
rect 12461 16374 12494 16408
rect 12528 16374 12562 16408
rect 12461 16318 12562 16374
rect 11274 16237 11375 16284
rect 12461 16284 12494 16318
rect 12528 16284 12562 16318
rect 12461 16237 12562 16284
rect 11274 16228 12562 16237
rect 11274 16194 11307 16228
rect 11341 16205 12494 16228
rect 11341 16194 11408 16205
rect 11274 16171 11408 16194
rect 11442 16171 11498 16205
rect 11532 16171 11588 16205
rect 11622 16171 11678 16205
rect 11712 16171 11768 16205
rect 11802 16171 11858 16205
rect 11892 16171 11948 16205
rect 11982 16171 12038 16205
rect 12072 16171 12128 16205
rect 12162 16171 12218 16205
rect 12252 16171 12308 16205
rect 12342 16171 12398 16205
rect 12432 16194 12494 16205
rect 12528 16194 12562 16228
rect 12432 16171 12562 16194
rect 11274 16136 12562 16171
rect 12634 17392 13922 17424
rect 12634 17358 12768 17392
rect 12802 17358 12858 17392
rect 12892 17358 12948 17392
rect 12982 17358 13038 17392
rect 13072 17358 13128 17392
rect 13162 17358 13218 17392
rect 13252 17358 13308 17392
rect 13342 17358 13398 17392
rect 13432 17358 13488 17392
rect 13522 17358 13578 17392
rect 13612 17358 13668 17392
rect 13702 17358 13758 17392
rect 13792 17358 13922 17392
rect 12634 17323 13922 17358
rect 12634 17308 12735 17323
rect 12634 17274 12667 17308
rect 12701 17274 12735 17308
rect 12634 17218 12735 17274
rect 13821 17308 13922 17323
rect 13821 17274 13854 17308
rect 13888 17274 13922 17308
rect 12634 17184 12667 17218
rect 12701 17184 12735 17218
rect 12634 17128 12735 17184
rect 12634 17094 12667 17128
rect 12701 17094 12735 17128
rect 12634 17038 12735 17094
rect 12634 17004 12667 17038
rect 12701 17004 12735 17038
rect 12634 16948 12735 17004
rect 12634 16914 12667 16948
rect 12701 16914 12735 16948
rect 12634 16858 12735 16914
rect 12634 16824 12667 16858
rect 12701 16824 12735 16858
rect 12634 16768 12735 16824
rect 12634 16734 12667 16768
rect 12701 16734 12735 16768
rect 12634 16678 12735 16734
rect 12634 16644 12667 16678
rect 12701 16644 12735 16678
rect 12634 16588 12735 16644
rect 12634 16554 12667 16588
rect 12701 16554 12735 16588
rect 12634 16498 12735 16554
rect 12634 16464 12667 16498
rect 12701 16464 12735 16498
rect 12634 16408 12735 16464
rect 12634 16374 12667 16408
rect 12701 16374 12735 16408
rect 12634 16318 12735 16374
rect 12634 16284 12667 16318
rect 12701 16284 12735 16318
rect 13821 17218 13922 17274
rect 13821 17184 13854 17218
rect 13888 17184 13922 17218
rect 13821 17128 13922 17184
rect 13821 17094 13854 17128
rect 13888 17094 13922 17128
rect 13821 17038 13922 17094
rect 13821 17004 13854 17038
rect 13888 17004 13922 17038
rect 13821 16948 13922 17004
rect 13821 16914 13854 16948
rect 13888 16914 13922 16948
rect 13821 16858 13922 16914
rect 13821 16824 13854 16858
rect 13888 16824 13922 16858
rect 13821 16768 13922 16824
rect 13821 16734 13854 16768
rect 13888 16734 13922 16768
rect 13821 16678 13922 16734
rect 13821 16644 13854 16678
rect 13888 16644 13922 16678
rect 13821 16588 13922 16644
rect 13821 16554 13854 16588
rect 13888 16554 13922 16588
rect 13821 16498 13922 16554
rect 13821 16464 13854 16498
rect 13888 16464 13922 16498
rect 13821 16408 13922 16464
rect 13821 16374 13854 16408
rect 13888 16374 13922 16408
rect 13821 16318 13922 16374
rect 12634 16237 12735 16284
rect 13821 16284 13854 16318
rect 13888 16284 13922 16318
rect 13821 16237 13922 16284
rect 12634 16228 13922 16237
rect 12634 16194 12667 16228
rect 12701 16205 13854 16228
rect 12701 16194 12768 16205
rect 12634 16171 12768 16194
rect 12802 16171 12858 16205
rect 12892 16171 12948 16205
rect 12982 16171 13038 16205
rect 13072 16171 13128 16205
rect 13162 16171 13218 16205
rect 13252 16171 13308 16205
rect 13342 16171 13398 16205
rect 13432 16171 13488 16205
rect 13522 16171 13578 16205
rect 13612 16171 13668 16205
rect 13702 16171 13758 16205
rect 13792 16194 13854 16205
rect 13888 16194 13922 16228
rect 13792 16171 13922 16194
rect 12634 16136 13922 16171
rect 13994 17392 15282 17424
rect 13994 17358 14128 17392
rect 14162 17358 14218 17392
rect 14252 17358 14308 17392
rect 14342 17358 14398 17392
rect 14432 17358 14488 17392
rect 14522 17358 14578 17392
rect 14612 17358 14668 17392
rect 14702 17358 14758 17392
rect 14792 17358 14848 17392
rect 14882 17358 14938 17392
rect 14972 17358 15028 17392
rect 15062 17358 15118 17392
rect 15152 17358 15282 17392
rect 13994 17323 15282 17358
rect 13994 17308 14095 17323
rect 13994 17274 14027 17308
rect 14061 17274 14095 17308
rect 13994 17218 14095 17274
rect 15181 17308 15282 17323
rect 15181 17274 15214 17308
rect 15248 17274 15282 17308
rect 13994 17184 14027 17218
rect 14061 17184 14095 17218
rect 13994 17128 14095 17184
rect 13994 17094 14027 17128
rect 14061 17094 14095 17128
rect 13994 17038 14095 17094
rect 13994 17004 14027 17038
rect 14061 17004 14095 17038
rect 13994 16948 14095 17004
rect 13994 16914 14027 16948
rect 14061 16914 14095 16948
rect 13994 16858 14095 16914
rect 13994 16824 14027 16858
rect 14061 16824 14095 16858
rect 13994 16768 14095 16824
rect 13994 16734 14027 16768
rect 14061 16734 14095 16768
rect 13994 16678 14095 16734
rect 13994 16644 14027 16678
rect 14061 16644 14095 16678
rect 13994 16588 14095 16644
rect 13994 16554 14027 16588
rect 14061 16554 14095 16588
rect 13994 16498 14095 16554
rect 13994 16464 14027 16498
rect 14061 16464 14095 16498
rect 13994 16408 14095 16464
rect 13994 16374 14027 16408
rect 14061 16374 14095 16408
rect 13994 16318 14095 16374
rect 13994 16284 14027 16318
rect 14061 16284 14095 16318
rect 15181 17218 15282 17274
rect 15181 17184 15214 17218
rect 15248 17184 15282 17218
rect 15181 17128 15282 17184
rect 15181 17094 15214 17128
rect 15248 17094 15282 17128
rect 15181 17038 15282 17094
rect 15181 17004 15214 17038
rect 15248 17004 15282 17038
rect 15181 16948 15282 17004
rect 15181 16914 15214 16948
rect 15248 16914 15282 16948
rect 15181 16858 15282 16914
rect 15181 16824 15214 16858
rect 15248 16824 15282 16858
rect 15181 16768 15282 16824
rect 15181 16734 15214 16768
rect 15248 16734 15282 16768
rect 15181 16678 15282 16734
rect 15181 16644 15214 16678
rect 15248 16644 15282 16678
rect 15181 16588 15282 16644
rect 15181 16554 15214 16588
rect 15248 16554 15282 16588
rect 15181 16498 15282 16554
rect 15181 16464 15214 16498
rect 15248 16464 15282 16498
rect 15181 16408 15282 16464
rect 15181 16374 15214 16408
rect 15248 16374 15282 16408
rect 15181 16318 15282 16374
rect 13994 16237 14095 16284
rect 15181 16284 15214 16318
rect 15248 16284 15282 16318
rect 15181 16237 15282 16284
rect 13994 16228 15282 16237
rect 13994 16194 14027 16228
rect 14061 16205 15214 16228
rect 14061 16194 14128 16205
rect 13994 16171 14128 16194
rect 14162 16171 14218 16205
rect 14252 16171 14308 16205
rect 14342 16171 14398 16205
rect 14432 16171 14488 16205
rect 14522 16171 14578 16205
rect 14612 16171 14668 16205
rect 14702 16171 14758 16205
rect 14792 16171 14848 16205
rect 14882 16171 14938 16205
rect 14972 16171 15028 16205
rect 15062 16171 15118 16205
rect 15152 16194 15214 16205
rect 15248 16194 15282 16228
rect 15152 16171 15282 16194
rect 13994 16136 15282 16171
rect 11274 16032 12562 16064
rect 11274 15998 11408 16032
rect 11442 15998 11498 16032
rect 11532 15998 11588 16032
rect 11622 15998 11678 16032
rect 11712 15998 11768 16032
rect 11802 15998 11858 16032
rect 11892 15998 11948 16032
rect 11982 15998 12038 16032
rect 12072 15998 12128 16032
rect 12162 15998 12218 16032
rect 12252 15998 12308 16032
rect 12342 15998 12398 16032
rect 12432 15998 12562 16032
rect 11274 15963 12562 15998
rect 11274 15948 11375 15963
rect 11274 15914 11307 15948
rect 11341 15914 11375 15948
rect 11274 15858 11375 15914
rect 12461 15948 12562 15963
rect 12461 15914 12494 15948
rect 12528 15914 12562 15948
rect 11274 15824 11307 15858
rect 11341 15824 11375 15858
rect 11274 15768 11375 15824
rect 11274 15734 11307 15768
rect 11341 15734 11375 15768
rect 11274 15678 11375 15734
rect 11274 15644 11307 15678
rect 11341 15644 11375 15678
rect 11274 15588 11375 15644
rect 11274 15554 11307 15588
rect 11341 15554 11375 15588
rect 11274 15498 11375 15554
rect 11274 15464 11307 15498
rect 11341 15464 11375 15498
rect 11274 15408 11375 15464
rect 11274 15374 11307 15408
rect 11341 15374 11375 15408
rect 11274 15318 11375 15374
rect 11274 15284 11307 15318
rect 11341 15284 11375 15318
rect 11274 15228 11375 15284
rect 11274 15194 11307 15228
rect 11341 15194 11375 15228
rect 11274 15138 11375 15194
rect 11274 15104 11307 15138
rect 11341 15104 11375 15138
rect 11274 15048 11375 15104
rect 11274 15014 11307 15048
rect 11341 15014 11375 15048
rect 11274 14958 11375 15014
rect 11274 14924 11307 14958
rect 11341 14924 11375 14958
rect 12461 15858 12562 15914
rect 12461 15824 12494 15858
rect 12528 15824 12562 15858
rect 12461 15768 12562 15824
rect 12461 15734 12494 15768
rect 12528 15734 12562 15768
rect 12461 15678 12562 15734
rect 12461 15644 12494 15678
rect 12528 15644 12562 15678
rect 12461 15588 12562 15644
rect 12461 15554 12494 15588
rect 12528 15554 12562 15588
rect 12461 15498 12562 15554
rect 12461 15464 12494 15498
rect 12528 15464 12562 15498
rect 12461 15408 12562 15464
rect 12461 15374 12494 15408
rect 12528 15374 12562 15408
rect 12461 15318 12562 15374
rect 12461 15284 12494 15318
rect 12528 15284 12562 15318
rect 12461 15228 12562 15284
rect 12461 15194 12494 15228
rect 12528 15194 12562 15228
rect 12461 15138 12562 15194
rect 12461 15104 12494 15138
rect 12528 15104 12562 15138
rect 12461 15048 12562 15104
rect 12461 15014 12494 15048
rect 12528 15014 12562 15048
rect 12461 14958 12562 15014
rect 11274 14877 11375 14924
rect 12461 14924 12494 14958
rect 12528 14924 12562 14958
rect 12461 14877 12562 14924
rect 11274 14868 12562 14877
rect 11274 14834 11307 14868
rect 11341 14845 12494 14868
rect 11341 14834 11408 14845
rect 11274 14811 11408 14834
rect 11442 14811 11498 14845
rect 11532 14811 11588 14845
rect 11622 14811 11678 14845
rect 11712 14811 11768 14845
rect 11802 14811 11858 14845
rect 11892 14811 11948 14845
rect 11982 14811 12038 14845
rect 12072 14811 12128 14845
rect 12162 14811 12218 14845
rect 12252 14811 12308 14845
rect 12342 14811 12398 14845
rect 12432 14834 12494 14845
rect 12528 14834 12562 14868
rect 12432 14811 12562 14834
rect 11274 14776 12562 14811
rect 12634 16032 13922 16064
rect 12634 15998 12768 16032
rect 12802 15998 12858 16032
rect 12892 15998 12948 16032
rect 12982 15998 13038 16032
rect 13072 15998 13128 16032
rect 13162 15998 13218 16032
rect 13252 15998 13308 16032
rect 13342 15998 13398 16032
rect 13432 15998 13488 16032
rect 13522 15998 13578 16032
rect 13612 15998 13668 16032
rect 13702 15998 13758 16032
rect 13792 15998 13922 16032
rect 12634 15963 13922 15998
rect 12634 15948 12735 15963
rect 12634 15914 12667 15948
rect 12701 15914 12735 15948
rect 12634 15858 12735 15914
rect 13821 15948 13922 15963
rect 13821 15914 13854 15948
rect 13888 15914 13922 15948
rect 12634 15824 12667 15858
rect 12701 15824 12735 15858
rect 12634 15768 12735 15824
rect 12634 15734 12667 15768
rect 12701 15734 12735 15768
rect 12634 15678 12735 15734
rect 12634 15644 12667 15678
rect 12701 15644 12735 15678
rect 12634 15588 12735 15644
rect 12634 15554 12667 15588
rect 12701 15554 12735 15588
rect 12634 15498 12735 15554
rect 12634 15464 12667 15498
rect 12701 15464 12735 15498
rect 12634 15408 12735 15464
rect 12634 15374 12667 15408
rect 12701 15374 12735 15408
rect 12634 15318 12735 15374
rect 12634 15284 12667 15318
rect 12701 15284 12735 15318
rect 12634 15228 12735 15284
rect 12634 15194 12667 15228
rect 12701 15194 12735 15228
rect 12634 15138 12735 15194
rect 12634 15104 12667 15138
rect 12701 15104 12735 15138
rect 12634 15048 12735 15104
rect 12634 15014 12667 15048
rect 12701 15014 12735 15048
rect 12634 14958 12735 15014
rect 12634 14924 12667 14958
rect 12701 14924 12735 14958
rect 13821 15858 13922 15914
rect 13821 15824 13854 15858
rect 13888 15824 13922 15858
rect 13821 15768 13922 15824
rect 13821 15734 13854 15768
rect 13888 15734 13922 15768
rect 13821 15678 13922 15734
rect 13821 15644 13854 15678
rect 13888 15644 13922 15678
rect 13821 15588 13922 15644
rect 13821 15554 13854 15588
rect 13888 15554 13922 15588
rect 13821 15498 13922 15554
rect 13821 15464 13854 15498
rect 13888 15464 13922 15498
rect 13821 15408 13922 15464
rect 13821 15374 13854 15408
rect 13888 15374 13922 15408
rect 13821 15318 13922 15374
rect 13821 15284 13854 15318
rect 13888 15284 13922 15318
rect 13821 15228 13922 15284
rect 13821 15194 13854 15228
rect 13888 15194 13922 15228
rect 13821 15138 13922 15194
rect 13821 15104 13854 15138
rect 13888 15104 13922 15138
rect 13821 15048 13922 15104
rect 13821 15014 13854 15048
rect 13888 15014 13922 15048
rect 13821 14958 13922 15014
rect 12634 14877 12735 14924
rect 13821 14924 13854 14958
rect 13888 14924 13922 14958
rect 13821 14877 13922 14924
rect 12634 14868 13922 14877
rect 12634 14834 12667 14868
rect 12701 14845 13854 14868
rect 12701 14834 12768 14845
rect 12634 14811 12768 14834
rect 12802 14811 12858 14845
rect 12892 14811 12948 14845
rect 12982 14811 13038 14845
rect 13072 14811 13128 14845
rect 13162 14811 13218 14845
rect 13252 14811 13308 14845
rect 13342 14811 13398 14845
rect 13432 14811 13488 14845
rect 13522 14811 13578 14845
rect 13612 14811 13668 14845
rect 13702 14811 13758 14845
rect 13792 14834 13854 14845
rect 13888 14834 13922 14868
rect 13792 14811 13922 14834
rect 12634 14776 13922 14811
rect 13994 16032 15282 16064
rect 13994 15998 14128 16032
rect 14162 15998 14218 16032
rect 14252 15998 14308 16032
rect 14342 15998 14398 16032
rect 14432 15998 14488 16032
rect 14522 15998 14578 16032
rect 14612 15998 14668 16032
rect 14702 15998 14758 16032
rect 14792 15998 14848 16032
rect 14882 15998 14938 16032
rect 14972 15998 15028 16032
rect 15062 15998 15118 16032
rect 15152 15998 15282 16032
rect 13994 15963 15282 15998
rect 13994 15948 14095 15963
rect 13994 15914 14027 15948
rect 14061 15914 14095 15948
rect 13994 15858 14095 15914
rect 15181 15948 15282 15963
rect 15181 15914 15214 15948
rect 15248 15914 15282 15948
rect 13994 15824 14027 15858
rect 14061 15824 14095 15858
rect 13994 15768 14095 15824
rect 13994 15734 14027 15768
rect 14061 15734 14095 15768
rect 13994 15678 14095 15734
rect 13994 15644 14027 15678
rect 14061 15644 14095 15678
rect 13994 15588 14095 15644
rect 13994 15554 14027 15588
rect 14061 15554 14095 15588
rect 13994 15498 14095 15554
rect 13994 15464 14027 15498
rect 14061 15464 14095 15498
rect 13994 15408 14095 15464
rect 13994 15374 14027 15408
rect 14061 15374 14095 15408
rect 13994 15318 14095 15374
rect 13994 15284 14027 15318
rect 14061 15284 14095 15318
rect 13994 15228 14095 15284
rect 13994 15194 14027 15228
rect 14061 15194 14095 15228
rect 13994 15138 14095 15194
rect 13994 15104 14027 15138
rect 14061 15104 14095 15138
rect 13994 15048 14095 15104
rect 13994 15014 14027 15048
rect 14061 15014 14095 15048
rect 13994 14958 14095 15014
rect 13994 14924 14027 14958
rect 14061 14924 14095 14958
rect 15181 15858 15282 15914
rect 15181 15824 15214 15858
rect 15248 15824 15282 15858
rect 15181 15768 15282 15824
rect 15181 15734 15214 15768
rect 15248 15734 15282 15768
rect 15181 15678 15282 15734
rect 15181 15644 15214 15678
rect 15248 15644 15282 15678
rect 15181 15588 15282 15644
rect 15181 15554 15214 15588
rect 15248 15554 15282 15588
rect 15181 15498 15282 15554
rect 15181 15464 15214 15498
rect 15248 15464 15282 15498
rect 15181 15408 15282 15464
rect 15181 15374 15214 15408
rect 15248 15374 15282 15408
rect 15181 15318 15282 15374
rect 15181 15284 15214 15318
rect 15248 15284 15282 15318
rect 15181 15228 15282 15284
rect 15181 15194 15214 15228
rect 15248 15194 15282 15228
rect 15181 15138 15282 15194
rect 15181 15104 15214 15138
rect 15248 15104 15282 15138
rect 15181 15048 15282 15104
rect 15181 15014 15214 15048
rect 15248 15014 15282 15048
rect 15181 14958 15282 15014
rect 13994 14877 14095 14924
rect 15181 14924 15214 14958
rect 15248 14924 15282 14958
rect 15181 14877 15282 14924
rect 13994 14868 15282 14877
rect 13994 14834 14027 14868
rect 14061 14845 15214 14868
rect 14061 14834 14128 14845
rect 13994 14811 14128 14834
rect 14162 14811 14218 14845
rect 14252 14811 14308 14845
rect 14342 14811 14398 14845
rect 14432 14811 14488 14845
rect 14522 14811 14578 14845
rect 14612 14811 14668 14845
rect 14702 14811 14758 14845
rect 14792 14811 14848 14845
rect 14882 14811 14938 14845
rect 14972 14811 15028 14845
rect 15062 14811 15118 14845
rect 15152 14834 15214 14845
rect 15248 14834 15282 14868
rect 15152 14811 15282 14834
rect 13994 14776 15282 14811
rect 15398 14250 15478 14280
rect 15398 14210 15418 14250
rect 15458 14210 15478 14250
rect 15398 14150 15478 14210
rect 15398 14110 15418 14150
rect 15458 14110 15478 14150
rect 15398 14080 15478 14110
rect 11898 13640 11978 13670
rect 11898 13600 11918 13640
rect 11958 13600 11978 13640
rect 11898 13540 11978 13600
rect 11898 13500 11918 13540
rect 11958 13500 11978 13540
rect 11898 13440 11978 13500
rect 11898 13400 11918 13440
rect 11958 13400 11978 13440
rect 11898 13340 11978 13400
rect 11898 13300 11918 13340
rect 11958 13300 11978 13340
rect 11898 13240 11978 13300
rect 11898 13200 11918 13240
rect 11958 13200 11978 13240
rect 11898 13170 11978 13200
rect 14578 13640 14658 13660
rect 14578 13600 14598 13640
rect 14638 13600 14658 13640
rect 14578 13540 14658 13600
rect 14578 13500 14598 13540
rect 14638 13500 14658 13540
rect 14578 13440 14658 13500
rect 14578 13400 14598 13440
rect 14638 13400 14658 13440
rect 14578 13340 14658 13400
rect 14578 13300 14598 13340
rect 14638 13300 14658 13340
rect 14578 13240 14658 13300
rect 14578 13200 14598 13240
rect 14638 13200 14658 13240
rect 14578 13170 14658 13200
rect 12798 12720 12878 12750
rect 12798 12680 12818 12720
rect 12858 12680 12878 12720
rect 12798 12640 12878 12680
rect 12798 12600 12818 12640
rect 12858 12600 12878 12640
rect 12798 12560 12878 12600
rect 12798 12520 12818 12560
rect 12858 12520 12878 12560
rect 12798 12490 12878 12520
rect 13678 12720 13758 12750
rect 13678 12680 13698 12720
rect 13738 12680 13758 12720
rect 13678 12640 13758 12680
rect 13678 12600 13698 12640
rect 13738 12600 13758 12640
rect 13678 12560 13758 12600
rect 13678 12520 13698 12560
rect 13738 12520 13758 12560
rect 13678 12490 13758 12520
rect 19338 11030 19438 11060
rect 19338 10990 19368 11030
rect 19408 10990 19438 11030
rect 19338 10960 19438 10990
rect 20318 11030 20418 11060
rect 20318 10990 20348 11030
rect 20388 10990 20418 11030
rect 20318 10960 20418 10990
rect 21618 11030 21718 11060
rect 21618 10990 21648 11030
rect 21688 10990 21718 11030
rect 21618 10960 21718 10990
rect 22598 11030 22698 11060
rect 22598 10990 22628 11030
rect 22668 10990 22698 11030
rect 22598 10960 22698 10990
rect 19288 10490 19388 10520
rect 19288 10440 19318 10490
rect 19358 10440 19388 10490
rect 19288 10350 19388 10440
rect 19288 10300 19318 10350
rect 19358 10300 19388 10350
rect 19288 10270 19388 10300
rect 21488 10490 21588 10520
rect 21488 10440 21518 10490
rect 21558 10440 21588 10490
rect 21488 10350 21588 10440
rect 21488 10300 21518 10350
rect 21558 10300 21588 10350
rect 21488 10270 21588 10300
rect 13168 8060 13248 8090
rect 13168 8020 13188 8060
rect 13228 8020 13248 8060
rect 13168 7960 13248 8020
rect 13168 7920 13188 7960
rect 13228 7920 13248 7960
rect 13168 7890 13248 7920
rect 14068 8060 14148 8090
rect 14068 8020 14088 8060
rect 14128 8020 14148 8060
rect 14068 7960 14148 8020
rect 14068 7920 14088 7960
rect 14128 7920 14148 7960
rect 14068 7890 14148 7920
rect 14968 8060 15048 8090
rect 14968 8020 14988 8060
rect 15028 8020 15048 8060
rect 14968 7960 15048 8020
rect 14968 7920 14988 7960
rect 15028 7920 15048 7960
rect 14968 7890 15048 7920
rect 15368 8060 15448 8090
rect 15368 8020 15388 8060
rect 15428 8020 15448 8060
rect 15368 7960 15448 8020
rect 15368 7920 15388 7960
rect 15428 7920 15448 7960
rect 15368 7890 15448 7920
rect 15698 8060 15778 8090
rect 15698 8020 15718 8060
rect 15758 8020 15778 8060
rect 15698 7960 15778 8020
rect 15698 7920 15718 7960
rect 15758 7920 15778 7960
rect 15698 7890 15778 7920
rect 16028 8060 16108 8090
rect 16028 8020 16048 8060
rect 16088 8020 16108 8060
rect 16028 7960 16108 8020
rect 16028 7920 16048 7960
rect 16088 7920 16108 7960
rect 16028 7890 16108 7920
rect 16278 8060 16378 8090
rect 16278 8020 16308 8060
rect 16348 8020 16378 8060
rect 16278 7960 16378 8020
rect 16278 7920 16308 7960
rect 16348 7920 16378 7960
rect 16278 7890 16378 7920
rect 17058 8060 17158 8090
rect 17058 8020 17088 8060
rect 17128 8020 17158 8060
rect 17058 7960 17158 8020
rect 17058 7920 17088 7960
rect 17128 7920 17158 7960
rect 17058 7890 17158 7920
rect 17738 8060 17838 8090
rect 17738 8020 17768 8060
rect 17808 8020 17838 8060
rect 17738 7960 17838 8020
rect 17738 7920 17768 7960
rect 17808 7920 17838 7960
rect 17738 7890 17838 7920
rect 19228 8010 19328 8040
rect 19228 7970 19258 8010
rect 19298 7970 19328 8010
rect 19228 7910 19328 7970
rect 19228 7870 19258 7910
rect 19298 7870 19328 7910
rect 19228 7810 19328 7870
rect 19228 7770 19258 7810
rect 19298 7770 19328 7810
rect 19228 7710 19328 7770
rect 19228 7670 19258 7710
rect 19298 7670 19328 7710
rect 19228 7640 19328 7670
rect 20308 8010 20408 8040
rect 20308 7970 20338 8010
rect 20378 7970 20408 8010
rect 20308 7910 20408 7970
rect 20308 7870 20338 7910
rect 20378 7870 20408 7910
rect 20308 7810 20408 7870
rect 20308 7770 20338 7810
rect 20378 7770 20408 7810
rect 20308 7710 20408 7770
rect 20308 7670 20338 7710
rect 20378 7670 20408 7710
rect 20308 7640 20408 7670
rect 21388 8010 21488 8040
rect 21388 7970 21418 8010
rect 21458 7970 21488 8010
rect 21388 7910 21488 7970
rect 21388 7870 21418 7910
rect 21458 7870 21488 7910
rect 21388 7810 21488 7870
rect 21388 7770 21418 7810
rect 21458 7770 21488 7810
rect 21388 7710 21488 7770
rect 21388 7670 21418 7710
rect 21458 7670 21488 7710
rect 21388 7640 21488 7670
rect 22468 8010 22568 8040
rect 22468 7970 22498 8010
rect 22538 7970 22568 8010
rect 22468 7910 22568 7970
rect 22468 7870 22498 7910
rect 22538 7870 22568 7910
rect 22468 7810 22568 7870
rect 22468 7770 22498 7810
rect 22538 7770 22568 7810
rect 22468 7710 22568 7770
rect 22468 7670 22498 7710
rect 22538 7670 22568 7710
rect 22468 7640 22568 7670
rect 13168 6260 13248 6290
rect 13168 6220 13188 6260
rect 13228 6220 13248 6260
rect 13168 6160 13248 6220
rect 13168 6120 13188 6160
rect 13228 6120 13248 6160
rect 13168 6090 13248 6120
rect 14068 6260 14148 6290
rect 14068 6220 14088 6260
rect 14128 6220 14148 6260
rect 14068 6160 14148 6220
rect 14068 6120 14088 6160
rect 14128 6120 14148 6160
rect 14068 6090 14148 6120
rect 14968 6260 15048 6290
rect 14968 6220 14988 6260
rect 15028 6220 15048 6260
rect 14968 6160 15048 6220
rect 14968 6120 14988 6160
rect 15028 6120 15048 6160
rect 14968 6090 15048 6120
rect 15108 6260 15188 6290
rect 15108 6220 15128 6260
rect 15168 6220 15188 6260
rect 15108 6160 15188 6220
rect 15108 6120 15128 6160
rect 15168 6120 15188 6160
rect 15108 6090 15188 6120
rect 15548 6260 15628 6290
rect 15548 6220 15568 6260
rect 15608 6220 15628 6260
rect 15548 6160 15628 6220
rect 15548 6120 15568 6160
rect 15608 6120 15628 6160
rect 15548 6090 15628 6120
rect 15878 6260 15958 6290
rect 15878 6220 15898 6260
rect 15938 6220 15958 6260
rect 15878 6160 15958 6220
rect 15878 6120 15898 6160
rect 15938 6120 15958 6160
rect 15878 6090 15958 6120
rect 16298 6260 16378 6290
rect 16298 6220 16318 6260
rect 16358 6220 16378 6260
rect 16298 6160 16378 6220
rect 16298 6120 16318 6160
rect 16358 6120 16378 6160
rect 16298 6090 16378 6120
rect 16688 6260 16768 6290
rect 16688 6220 16708 6260
rect 16748 6220 16768 6260
rect 16688 6160 16768 6220
rect 16688 6120 16708 6160
rect 16748 6120 16768 6160
rect 16688 6090 16768 6120
rect 17078 6260 17158 6290
rect 17078 6220 17098 6260
rect 17138 6220 17158 6260
rect 17078 6160 17158 6220
rect 17078 6120 17098 6160
rect 17138 6120 17158 6160
rect 17078 6090 17158 6120
rect 15678 3180 15758 3210
rect 15678 3140 15698 3180
rect 15738 3140 15758 3180
rect 15678 3110 15758 3140
rect 17128 3180 17208 3210
rect 17128 3140 17148 3180
rect 17188 3140 17208 3180
rect 17128 3110 17208 3140
rect 23088 3180 24228 3220
rect 24368 3180 25128 3220
rect 18918 3090 18998 3120
rect 18918 3050 18938 3090
rect 18978 3050 18998 3090
rect 18918 3020 18998 3050
rect 20218 3090 20298 3120
rect 20218 3050 20238 3090
rect 20278 3050 20298 3090
rect 20218 3020 20298 3050
rect 21518 3090 21598 3120
rect 21518 3050 21538 3090
rect 21578 3050 21598 3090
rect 21518 3020 21598 3050
rect 23088 2660 23128 3180
rect 25088 2660 25128 3180
rect 23088 1920 23128 2450
rect 25088 1920 25128 2450
rect 23088 1880 24228 1920
rect 24368 1880 25128 1920
<< nsubdiff >>
rect 14851 19663 14947 19697
rect 17369 19663 17465 19697
rect 14851 19601 14885 19663
rect 17431 19601 17465 19663
rect 14851 19279 14885 19341
rect 17431 19279 17465 19341
rect 14851 19245 14947 19279
rect 17369 19245 17465 19279
rect 8261 18563 8357 18597
rect 8617 18563 8713 18597
rect 8261 18501 8295 18563
rect 8679 18501 8713 18563
rect 8261 17111 8295 17173
rect 8679 17111 8713 17173
rect 8261 17077 8357 17111
rect 8617 17077 8713 17111
rect 9048 18566 9144 18600
rect 9736 18566 9832 18600
rect 9048 18504 9082 18566
rect 9798 18504 9832 18566
rect 9048 16712 9082 16774
rect 9798 16712 9832 16774
rect 9048 16678 9144 16712
rect 9736 16678 9832 16712
rect 10161 18563 10257 18597
rect 10849 18563 10945 18597
rect 10161 18501 10195 18563
rect 10911 18501 10945 18563
rect 10161 16181 10195 16243
rect 11437 18602 12399 18621
rect 11437 18568 11548 18602
rect 11582 18568 11638 18602
rect 11672 18568 11728 18602
rect 11762 18568 11818 18602
rect 11852 18568 11908 18602
rect 11942 18568 11998 18602
rect 12032 18568 12088 18602
rect 12122 18568 12178 18602
rect 12212 18568 12268 18602
rect 12302 18568 12399 18602
rect 11437 18549 12399 18568
rect 11437 18508 11509 18549
rect 11437 18474 11456 18508
rect 11490 18474 11509 18508
rect 12327 18489 12399 18549
rect 11437 18418 11509 18474
rect 11437 18384 11456 18418
rect 11490 18384 11509 18418
rect 11437 18328 11509 18384
rect 11437 18294 11456 18328
rect 11490 18294 11509 18328
rect 11437 18238 11509 18294
rect 11437 18204 11456 18238
rect 11490 18204 11509 18238
rect 11437 18148 11509 18204
rect 11437 18114 11456 18148
rect 11490 18114 11509 18148
rect 11437 18058 11509 18114
rect 11437 18024 11456 18058
rect 11490 18024 11509 18058
rect 11437 17968 11509 18024
rect 11437 17934 11456 17968
rect 11490 17934 11509 17968
rect 11437 17878 11509 17934
rect 11437 17844 11456 17878
rect 11490 17844 11509 17878
rect 11437 17788 11509 17844
rect 12327 18455 12346 18489
rect 12380 18455 12399 18489
rect 12327 18399 12399 18455
rect 12327 18365 12346 18399
rect 12380 18365 12399 18399
rect 12327 18309 12399 18365
rect 12327 18275 12346 18309
rect 12380 18275 12399 18309
rect 12327 18219 12399 18275
rect 12327 18185 12346 18219
rect 12380 18185 12399 18219
rect 12327 18129 12399 18185
rect 12327 18095 12346 18129
rect 12380 18095 12399 18129
rect 12327 18039 12399 18095
rect 12327 18005 12346 18039
rect 12380 18005 12399 18039
rect 12327 17949 12399 18005
rect 12327 17915 12346 17949
rect 12380 17915 12399 17949
rect 12327 17859 12399 17915
rect 12327 17825 12346 17859
rect 12380 17825 12399 17859
rect 11437 17754 11456 17788
rect 11490 17754 11509 17788
rect 11437 17731 11509 17754
rect 12327 17769 12399 17825
rect 12327 17735 12346 17769
rect 12380 17735 12399 17769
rect 12327 17731 12399 17735
rect 11437 17712 12399 17731
rect 11437 17678 11514 17712
rect 11548 17678 11604 17712
rect 11638 17678 11694 17712
rect 11728 17678 11784 17712
rect 11818 17678 11874 17712
rect 11908 17678 11964 17712
rect 11998 17678 12054 17712
rect 12088 17678 12144 17712
rect 12178 17678 12234 17712
rect 12268 17678 12399 17712
rect 11437 17659 12399 17678
rect 12797 18602 13759 18621
rect 12797 18568 12908 18602
rect 12942 18568 12998 18602
rect 13032 18568 13088 18602
rect 13122 18568 13178 18602
rect 13212 18568 13268 18602
rect 13302 18568 13358 18602
rect 13392 18568 13448 18602
rect 13482 18568 13538 18602
rect 13572 18568 13628 18602
rect 13662 18568 13759 18602
rect 12797 18549 13759 18568
rect 12797 18508 12869 18549
rect 12797 18474 12816 18508
rect 12850 18474 12869 18508
rect 13687 18489 13759 18549
rect 12797 18418 12869 18474
rect 12797 18384 12816 18418
rect 12850 18384 12869 18418
rect 12797 18328 12869 18384
rect 12797 18294 12816 18328
rect 12850 18294 12869 18328
rect 12797 18238 12869 18294
rect 12797 18204 12816 18238
rect 12850 18204 12869 18238
rect 12797 18148 12869 18204
rect 12797 18114 12816 18148
rect 12850 18114 12869 18148
rect 12797 18058 12869 18114
rect 12797 18024 12816 18058
rect 12850 18024 12869 18058
rect 12797 17968 12869 18024
rect 12797 17934 12816 17968
rect 12850 17934 12869 17968
rect 12797 17878 12869 17934
rect 12797 17844 12816 17878
rect 12850 17844 12869 17878
rect 12797 17788 12869 17844
rect 13687 18455 13706 18489
rect 13740 18455 13759 18489
rect 13687 18399 13759 18455
rect 13687 18365 13706 18399
rect 13740 18365 13759 18399
rect 13687 18309 13759 18365
rect 13687 18275 13706 18309
rect 13740 18275 13759 18309
rect 13687 18219 13759 18275
rect 13687 18185 13706 18219
rect 13740 18185 13759 18219
rect 13687 18129 13759 18185
rect 13687 18095 13706 18129
rect 13740 18095 13759 18129
rect 13687 18039 13759 18095
rect 13687 18005 13706 18039
rect 13740 18005 13759 18039
rect 13687 17949 13759 18005
rect 13687 17915 13706 17949
rect 13740 17915 13759 17949
rect 13687 17859 13759 17915
rect 13687 17825 13706 17859
rect 13740 17825 13759 17859
rect 12797 17754 12816 17788
rect 12850 17754 12869 17788
rect 12797 17731 12869 17754
rect 13687 17769 13759 17825
rect 13687 17735 13706 17769
rect 13740 17735 13759 17769
rect 13687 17731 13759 17735
rect 12797 17712 13759 17731
rect 12797 17678 12874 17712
rect 12908 17678 12964 17712
rect 12998 17678 13054 17712
rect 13088 17678 13144 17712
rect 13178 17678 13234 17712
rect 13268 17678 13324 17712
rect 13358 17678 13414 17712
rect 13448 17678 13504 17712
rect 13538 17678 13594 17712
rect 13628 17678 13759 17712
rect 12797 17659 13759 17678
rect 14157 18602 15119 18621
rect 14157 18568 14268 18602
rect 14302 18568 14358 18602
rect 14392 18568 14448 18602
rect 14482 18568 14538 18602
rect 14572 18568 14628 18602
rect 14662 18568 14718 18602
rect 14752 18568 14808 18602
rect 14842 18568 14898 18602
rect 14932 18568 14988 18602
rect 15022 18568 15119 18602
rect 14157 18549 15119 18568
rect 14157 18508 14229 18549
rect 14157 18474 14176 18508
rect 14210 18474 14229 18508
rect 15047 18489 15119 18549
rect 14157 18418 14229 18474
rect 14157 18384 14176 18418
rect 14210 18384 14229 18418
rect 14157 18328 14229 18384
rect 14157 18294 14176 18328
rect 14210 18294 14229 18328
rect 14157 18238 14229 18294
rect 14157 18204 14176 18238
rect 14210 18204 14229 18238
rect 14157 18148 14229 18204
rect 14157 18114 14176 18148
rect 14210 18114 14229 18148
rect 14157 18058 14229 18114
rect 14157 18024 14176 18058
rect 14210 18024 14229 18058
rect 14157 17968 14229 18024
rect 14157 17934 14176 17968
rect 14210 17934 14229 17968
rect 14157 17878 14229 17934
rect 14157 17844 14176 17878
rect 14210 17844 14229 17878
rect 14157 17788 14229 17844
rect 15047 18455 15066 18489
rect 15100 18455 15119 18489
rect 15047 18399 15119 18455
rect 15047 18365 15066 18399
rect 15100 18365 15119 18399
rect 15047 18309 15119 18365
rect 15047 18275 15066 18309
rect 15100 18275 15119 18309
rect 15047 18219 15119 18275
rect 15047 18185 15066 18219
rect 15100 18185 15119 18219
rect 15047 18129 15119 18185
rect 15047 18095 15066 18129
rect 15100 18095 15119 18129
rect 15047 18039 15119 18095
rect 15047 18005 15066 18039
rect 15100 18005 15119 18039
rect 15047 17949 15119 18005
rect 15047 17915 15066 17949
rect 15100 17915 15119 17949
rect 15047 17859 15119 17915
rect 15047 17825 15066 17859
rect 15100 17825 15119 17859
rect 14157 17754 14176 17788
rect 14210 17754 14229 17788
rect 14157 17731 14229 17754
rect 15047 17769 15119 17825
rect 15047 17735 15066 17769
rect 15100 17735 15119 17769
rect 15047 17731 15119 17735
rect 14157 17712 15119 17731
rect 14157 17678 14234 17712
rect 14268 17678 14324 17712
rect 14358 17678 14414 17712
rect 14448 17678 14504 17712
rect 14538 17678 14594 17712
rect 14628 17678 14684 17712
rect 14718 17678 14774 17712
rect 14808 17678 14864 17712
rect 14898 17678 14954 17712
rect 14988 17678 15119 17712
rect 14157 17659 15119 17678
rect 15481 18563 15577 18597
rect 16169 18563 16265 18597
rect 15481 18501 15515 18563
rect 10911 16181 10945 16243
rect 10161 16147 10257 16181
rect 10849 16147 10945 16181
rect 11437 17242 12399 17261
rect 11437 17208 11548 17242
rect 11582 17208 11638 17242
rect 11672 17208 11728 17242
rect 11762 17208 11818 17242
rect 11852 17208 11908 17242
rect 11942 17208 11998 17242
rect 12032 17208 12088 17242
rect 12122 17208 12178 17242
rect 12212 17208 12268 17242
rect 12302 17208 12399 17242
rect 11437 17189 12399 17208
rect 11437 17148 11509 17189
rect 11437 17114 11456 17148
rect 11490 17114 11509 17148
rect 12327 17129 12399 17189
rect 11437 17058 11509 17114
rect 11437 17024 11456 17058
rect 11490 17024 11509 17058
rect 11437 16968 11509 17024
rect 11437 16934 11456 16968
rect 11490 16934 11509 16968
rect 11437 16878 11509 16934
rect 11437 16844 11456 16878
rect 11490 16844 11509 16878
rect 11437 16788 11509 16844
rect 11437 16754 11456 16788
rect 11490 16754 11509 16788
rect 11437 16698 11509 16754
rect 11437 16664 11456 16698
rect 11490 16664 11509 16698
rect 11437 16608 11509 16664
rect 11437 16574 11456 16608
rect 11490 16574 11509 16608
rect 11437 16518 11509 16574
rect 11437 16484 11456 16518
rect 11490 16484 11509 16518
rect 11437 16428 11509 16484
rect 12327 17095 12346 17129
rect 12380 17095 12399 17129
rect 12327 17039 12399 17095
rect 12327 17005 12346 17039
rect 12380 17005 12399 17039
rect 12327 16949 12399 17005
rect 12327 16915 12346 16949
rect 12380 16915 12399 16949
rect 12327 16859 12399 16915
rect 12327 16825 12346 16859
rect 12380 16825 12399 16859
rect 12327 16769 12399 16825
rect 12327 16735 12346 16769
rect 12380 16735 12399 16769
rect 12327 16679 12399 16735
rect 12327 16645 12346 16679
rect 12380 16645 12399 16679
rect 12327 16589 12399 16645
rect 12327 16555 12346 16589
rect 12380 16555 12399 16589
rect 12327 16499 12399 16555
rect 12327 16465 12346 16499
rect 12380 16465 12399 16499
rect 11437 16394 11456 16428
rect 11490 16394 11509 16428
rect 11437 16371 11509 16394
rect 12327 16409 12399 16465
rect 12327 16375 12346 16409
rect 12380 16375 12399 16409
rect 12327 16371 12399 16375
rect 11437 16352 12399 16371
rect 11437 16318 11514 16352
rect 11548 16318 11604 16352
rect 11638 16318 11694 16352
rect 11728 16318 11784 16352
rect 11818 16318 11874 16352
rect 11908 16318 11964 16352
rect 11998 16318 12054 16352
rect 12088 16318 12144 16352
rect 12178 16318 12234 16352
rect 12268 16318 12399 16352
rect 11437 16299 12399 16318
rect 12797 17242 13759 17261
rect 12797 17208 12908 17242
rect 12942 17208 12998 17242
rect 13032 17208 13088 17242
rect 13122 17208 13178 17242
rect 13212 17208 13268 17242
rect 13302 17208 13358 17242
rect 13392 17208 13448 17242
rect 13482 17208 13538 17242
rect 13572 17208 13628 17242
rect 13662 17208 13759 17242
rect 12797 17189 13759 17208
rect 12797 17148 12869 17189
rect 12797 17114 12816 17148
rect 12850 17114 12869 17148
rect 13687 17129 13759 17189
rect 12797 17058 12869 17114
rect 12797 17024 12816 17058
rect 12850 17024 12869 17058
rect 12797 16968 12869 17024
rect 12797 16934 12816 16968
rect 12850 16934 12869 16968
rect 12797 16878 12869 16934
rect 12797 16844 12816 16878
rect 12850 16844 12869 16878
rect 12797 16788 12869 16844
rect 12797 16754 12816 16788
rect 12850 16754 12869 16788
rect 12797 16698 12869 16754
rect 12797 16664 12816 16698
rect 12850 16664 12869 16698
rect 12797 16608 12869 16664
rect 12797 16574 12816 16608
rect 12850 16574 12869 16608
rect 12797 16518 12869 16574
rect 12797 16484 12816 16518
rect 12850 16484 12869 16518
rect 12797 16428 12869 16484
rect 13687 17095 13706 17129
rect 13740 17095 13759 17129
rect 13687 17039 13759 17095
rect 13687 17005 13706 17039
rect 13740 17005 13759 17039
rect 13687 16949 13759 17005
rect 13687 16915 13706 16949
rect 13740 16915 13759 16949
rect 13687 16859 13759 16915
rect 13687 16825 13706 16859
rect 13740 16825 13759 16859
rect 13687 16769 13759 16825
rect 13687 16735 13706 16769
rect 13740 16735 13759 16769
rect 13687 16679 13759 16735
rect 13687 16645 13706 16679
rect 13740 16645 13759 16679
rect 13687 16589 13759 16645
rect 13687 16555 13706 16589
rect 13740 16555 13759 16589
rect 13687 16499 13759 16555
rect 13687 16465 13706 16499
rect 13740 16465 13759 16499
rect 12797 16394 12816 16428
rect 12850 16394 12869 16428
rect 12797 16371 12869 16394
rect 13687 16409 13759 16465
rect 13687 16375 13706 16409
rect 13740 16375 13759 16409
rect 13687 16371 13759 16375
rect 12797 16352 13759 16371
rect 12797 16318 12874 16352
rect 12908 16318 12964 16352
rect 12998 16318 13054 16352
rect 13088 16318 13144 16352
rect 13178 16318 13234 16352
rect 13268 16318 13324 16352
rect 13358 16318 13414 16352
rect 13448 16318 13504 16352
rect 13538 16318 13594 16352
rect 13628 16318 13759 16352
rect 12797 16299 13759 16318
rect 14157 17242 15119 17261
rect 14157 17208 14268 17242
rect 14302 17208 14358 17242
rect 14392 17208 14448 17242
rect 14482 17208 14538 17242
rect 14572 17208 14628 17242
rect 14662 17208 14718 17242
rect 14752 17208 14808 17242
rect 14842 17208 14898 17242
rect 14932 17208 14988 17242
rect 15022 17208 15119 17242
rect 14157 17189 15119 17208
rect 14157 17148 14229 17189
rect 14157 17114 14176 17148
rect 14210 17114 14229 17148
rect 15047 17129 15119 17189
rect 14157 17058 14229 17114
rect 14157 17024 14176 17058
rect 14210 17024 14229 17058
rect 14157 16968 14229 17024
rect 14157 16934 14176 16968
rect 14210 16934 14229 16968
rect 14157 16878 14229 16934
rect 14157 16844 14176 16878
rect 14210 16844 14229 16878
rect 14157 16788 14229 16844
rect 14157 16754 14176 16788
rect 14210 16754 14229 16788
rect 14157 16698 14229 16754
rect 14157 16664 14176 16698
rect 14210 16664 14229 16698
rect 14157 16608 14229 16664
rect 14157 16574 14176 16608
rect 14210 16574 14229 16608
rect 14157 16518 14229 16574
rect 14157 16484 14176 16518
rect 14210 16484 14229 16518
rect 14157 16428 14229 16484
rect 15047 17095 15066 17129
rect 15100 17095 15119 17129
rect 15047 17039 15119 17095
rect 15047 17005 15066 17039
rect 15100 17005 15119 17039
rect 15047 16949 15119 17005
rect 15047 16915 15066 16949
rect 15100 16915 15119 16949
rect 15047 16859 15119 16915
rect 15047 16825 15066 16859
rect 15100 16825 15119 16859
rect 15047 16769 15119 16825
rect 15047 16735 15066 16769
rect 15100 16735 15119 16769
rect 15047 16679 15119 16735
rect 15047 16645 15066 16679
rect 15100 16645 15119 16679
rect 15047 16589 15119 16645
rect 15047 16555 15066 16589
rect 15100 16555 15119 16589
rect 15047 16499 15119 16555
rect 15047 16465 15066 16499
rect 15100 16465 15119 16499
rect 14157 16394 14176 16428
rect 14210 16394 14229 16428
rect 14157 16371 14229 16394
rect 15047 16409 15119 16465
rect 15047 16375 15066 16409
rect 15100 16375 15119 16409
rect 15047 16371 15119 16375
rect 14157 16352 15119 16371
rect 14157 16318 14234 16352
rect 14268 16318 14324 16352
rect 14358 16318 14414 16352
rect 14448 16318 14504 16352
rect 14538 16318 14594 16352
rect 14628 16318 14684 16352
rect 14718 16318 14774 16352
rect 14808 16318 14864 16352
rect 14898 16318 14954 16352
rect 14988 16318 15119 16352
rect 14157 16299 15119 16318
rect 16231 18501 16265 18563
rect 15481 16181 15515 16243
rect 16594 18560 16690 18594
rect 16950 18560 17046 18594
rect 16594 18498 16628 18560
rect 17012 18498 17046 18560
rect 16594 17318 16628 17380
rect 17012 17318 17046 17380
rect 16594 17284 16690 17318
rect 16950 17284 17046 17318
rect 17381 18563 17477 18597
rect 17737 18563 17833 18597
rect 17381 18501 17415 18563
rect 17799 18501 17833 18563
rect 17381 17111 17415 17173
rect 17799 17111 17833 17173
rect 17381 17077 17477 17111
rect 17737 17077 17833 17111
rect 16231 16181 16265 16243
rect 15481 16147 15577 16181
rect 16169 16147 16265 16181
rect 11437 15882 12399 15901
rect 11437 15848 11548 15882
rect 11582 15848 11638 15882
rect 11672 15848 11728 15882
rect 11762 15848 11818 15882
rect 11852 15848 11908 15882
rect 11942 15848 11998 15882
rect 12032 15848 12088 15882
rect 12122 15848 12178 15882
rect 12212 15848 12268 15882
rect 12302 15848 12399 15882
rect 11437 15829 12399 15848
rect 11437 15788 11509 15829
rect 11437 15754 11456 15788
rect 11490 15754 11509 15788
rect 12327 15769 12399 15829
rect 11437 15698 11509 15754
rect 11437 15664 11456 15698
rect 11490 15664 11509 15698
rect 11437 15608 11509 15664
rect 11437 15574 11456 15608
rect 11490 15574 11509 15608
rect 11437 15518 11509 15574
rect 11437 15484 11456 15518
rect 11490 15484 11509 15518
rect 11437 15428 11509 15484
rect 11437 15394 11456 15428
rect 11490 15394 11509 15428
rect 11437 15338 11509 15394
rect 11437 15304 11456 15338
rect 11490 15304 11509 15338
rect 11437 15248 11509 15304
rect 11437 15214 11456 15248
rect 11490 15214 11509 15248
rect 11437 15158 11509 15214
rect 11437 15124 11456 15158
rect 11490 15124 11509 15158
rect 11437 15068 11509 15124
rect 12327 15735 12346 15769
rect 12380 15735 12399 15769
rect 12327 15679 12399 15735
rect 12327 15645 12346 15679
rect 12380 15645 12399 15679
rect 12327 15589 12399 15645
rect 12327 15555 12346 15589
rect 12380 15555 12399 15589
rect 12327 15499 12399 15555
rect 12327 15465 12346 15499
rect 12380 15465 12399 15499
rect 12327 15409 12399 15465
rect 12327 15375 12346 15409
rect 12380 15375 12399 15409
rect 12327 15319 12399 15375
rect 12327 15285 12346 15319
rect 12380 15285 12399 15319
rect 12327 15229 12399 15285
rect 12327 15195 12346 15229
rect 12380 15195 12399 15229
rect 12327 15139 12399 15195
rect 12327 15105 12346 15139
rect 12380 15105 12399 15139
rect 11437 15034 11456 15068
rect 11490 15034 11509 15068
rect 11437 15011 11509 15034
rect 12327 15049 12399 15105
rect 12327 15015 12346 15049
rect 12380 15015 12399 15049
rect 12327 15011 12399 15015
rect 11437 14992 12399 15011
rect 11437 14958 11514 14992
rect 11548 14958 11604 14992
rect 11638 14958 11694 14992
rect 11728 14958 11784 14992
rect 11818 14958 11874 14992
rect 11908 14958 11964 14992
rect 11998 14958 12054 14992
rect 12088 14958 12144 14992
rect 12178 14958 12234 14992
rect 12268 14958 12399 14992
rect 11437 14939 12399 14958
rect 12797 15882 13759 15901
rect 12797 15848 12908 15882
rect 12942 15848 12998 15882
rect 13032 15848 13088 15882
rect 13122 15848 13178 15882
rect 13212 15848 13268 15882
rect 13302 15848 13358 15882
rect 13392 15848 13448 15882
rect 13482 15848 13538 15882
rect 13572 15848 13628 15882
rect 13662 15848 13759 15882
rect 12797 15829 13759 15848
rect 12797 15788 12869 15829
rect 12797 15754 12816 15788
rect 12850 15754 12869 15788
rect 13687 15769 13759 15829
rect 12797 15698 12869 15754
rect 12797 15664 12816 15698
rect 12850 15664 12869 15698
rect 12797 15608 12869 15664
rect 12797 15574 12816 15608
rect 12850 15574 12869 15608
rect 12797 15518 12869 15574
rect 12797 15484 12816 15518
rect 12850 15484 12869 15518
rect 12797 15428 12869 15484
rect 12797 15394 12816 15428
rect 12850 15394 12869 15428
rect 12797 15338 12869 15394
rect 12797 15304 12816 15338
rect 12850 15304 12869 15338
rect 12797 15248 12869 15304
rect 12797 15214 12816 15248
rect 12850 15214 12869 15248
rect 12797 15158 12869 15214
rect 12797 15124 12816 15158
rect 12850 15124 12869 15158
rect 12797 15068 12869 15124
rect 13687 15735 13706 15769
rect 13740 15735 13759 15769
rect 13687 15679 13759 15735
rect 13687 15645 13706 15679
rect 13740 15645 13759 15679
rect 13687 15589 13759 15645
rect 13687 15555 13706 15589
rect 13740 15555 13759 15589
rect 13687 15499 13759 15555
rect 13687 15465 13706 15499
rect 13740 15465 13759 15499
rect 13687 15409 13759 15465
rect 13687 15375 13706 15409
rect 13740 15375 13759 15409
rect 13687 15319 13759 15375
rect 13687 15285 13706 15319
rect 13740 15285 13759 15319
rect 13687 15229 13759 15285
rect 13687 15195 13706 15229
rect 13740 15195 13759 15229
rect 13687 15139 13759 15195
rect 13687 15105 13706 15139
rect 13740 15105 13759 15139
rect 12797 15034 12816 15068
rect 12850 15034 12869 15068
rect 12797 15011 12869 15034
rect 13687 15049 13759 15105
rect 13687 15015 13706 15049
rect 13740 15015 13759 15049
rect 13687 15011 13759 15015
rect 12797 14992 13759 15011
rect 12797 14958 12874 14992
rect 12908 14958 12964 14992
rect 12998 14958 13054 14992
rect 13088 14958 13144 14992
rect 13178 14958 13234 14992
rect 13268 14958 13324 14992
rect 13358 14958 13414 14992
rect 13448 14958 13504 14992
rect 13538 14958 13594 14992
rect 13628 14958 13759 14992
rect 12797 14939 13759 14958
rect 14157 15882 15119 15901
rect 14157 15848 14268 15882
rect 14302 15848 14358 15882
rect 14392 15848 14448 15882
rect 14482 15848 14538 15882
rect 14572 15848 14628 15882
rect 14662 15848 14718 15882
rect 14752 15848 14808 15882
rect 14842 15848 14898 15882
rect 14932 15848 14988 15882
rect 15022 15848 15119 15882
rect 14157 15829 15119 15848
rect 14157 15788 14229 15829
rect 14157 15754 14176 15788
rect 14210 15754 14229 15788
rect 15047 15769 15119 15829
rect 14157 15698 14229 15754
rect 14157 15664 14176 15698
rect 14210 15664 14229 15698
rect 14157 15608 14229 15664
rect 14157 15574 14176 15608
rect 14210 15574 14229 15608
rect 14157 15518 14229 15574
rect 14157 15484 14176 15518
rect 14210 15484 14229 15518
rect 14157 15428 14229 15484
rect 14157 15394 14176 15428
rect 14210 15394 14229 15428
rect 14157 15338 14229 15394
rect 14157 15304 14176 15338
rect 14210 15304 14229 15338
rect 14157 15248 14229 15304
rect 14157 15214 14176 15248
rect 14210 15214 14229 15248
rect 14157 15158 14229 15214
rect 14157 15124 14176 15158
rect 14210 15124 14229 15158
rect 14157 15068 14229 15124
rect 15047 15735 15066 15769
rect 15100 15735 15119 15769
rect 15047 15679 15119 15735
rect 15047 15645 15066 15679
rect 15100 15645 15119 15679
rect 15047 15589 15119 15645
rect 15047 15555 15066 15589
rect 15100 15555 15119 15589
rect 15047 15499 15119 15555
rect 15047 15465 15066 15499
rect 15100 15465 15119 15499
rect 15047 15409 15119 15465
rect 15047 15375 15066 15409
rect 15100 15375 15119 15409
rect 15047 15319 15119 15375
rect 15047 15285 15066 15319
rect 15100 15285 15119 15319
rect 15047 15229 15119 15285
rect 15047 15195 15066 15229
rect 15100 15195 15119 15229
rect 15047 15139 15119 15195
rect 15047 15105 15066 15139
rect 15100 15105 15119 15139
rect 14157 15034 14176 15068
rect 14210 15034 14229 15068
rect 14157 15011 14229 15034
rect 15047 15049 15119 15105
rect 15047 15015 15066 15049
rect 15100 15015 15119 15049
rect 15047 15011 15119 15015
rect 14157 14992 15119 15011
rect 14157 14958 14234 14992
rect 14268 14958 14324 14992
rect 14358 14958 14414 14992
rect 14448 14958 14504 14992
rect 14538 14958 14594 14992
rect 14628 14958 14684 14992
rect 14718 14958 14774 14992
rect 14808 14958 14864 14992
rect 14898 14958 14954 14992
rect 14988 14958 15119 14992
rect 14157 14939 15119 14958
rect 23031 13253 23127 13287
rect 23387 13253 23483 13287
rect 23031 13191 23065 13253
rect 19408 12660 19508 12690
rect 19408 12620 19438 12660
rect 19478 12620 19508 12660
rect 19408 12560 19508 12620
rect 19408 12520 19438 12560
rect 19478 12520 19508 12560
rect 19408 12460 19508 12520
rect 19408 12420 19438 12460
rect 19478 12420 19508 12460
rect 19408 12360 19508 12420
rect 19408 12320 19438 12360
rect 19478 12320 19508 12360
rect 19408 12260 19508 12320
rect 19408 12220 19438 12260
rect 19478 12220 19508 12260
rect 19408 12190 19508 12220
rect 21608 12660 21708 12690
rect 21608 12620 21638 12660
rect 21678 12620 21708 12660
rect 21608 12560 21708 12620
rect 21608 12520 21638 12560
rect 21678 12520 21708 12560
rect 21608 12460 21708 12520
rect 21608 12420 21638 12460
rect 21678 12420 21708 12460
rect 21608 12360 21708 12420
rect 21608 12320 21638 12360
rect 21678 12320 21708 12360
rect 21608 12260 21708 12320
rect 21608 12220 21638 12260
rect 21678 12220 21708 12260
rect 21608 12190 21708 12220
rect 23449 13191 23483 13253
rect 23031 11983 23065 12045
rect 23449 11983 23483 12045
rect 23031 11949 23127 11983
rect 23387 11949 23483 11983
rect 10438 11790 10518 11820
rect 10438 11750 10458 11790
rect 10498 11750 10518 11790
rect 10438 11690 10518 11750
rect 10438 11650 10458 11690
rect 10498 11650 10518 11690
rect 10438 11620 10518 11650
rect 12998 11790 13078 11820
rect 12998 11750 13018 11790
rect 13058 11750 13078 11790
rect 12998 11690 13078 11750
rect 12998 11650 13018 11690
rect 13058 11650 13078 11690
rect 12998 11620 13078 11650
rect 13478 11790 13558 11820
rect 13478 11750 13498 11790
rect 13538 11750 13558 11790
rect 13478 11690 13558 11750
rect 13478 11650 13498 11690
rect 13538 11650 13558 11690
rect 13478 11620 13558 11650
rect 16038 11790 16118 11820
rect 16038 11750 16058 11790
rect 16098 11750 16118 11790
rect 16038 11690 16118 11750
rect 16038 11650 16058 11690
rect 16098 11650 16118 11690
rect 16038 11620 16118 11650
rect 20478 11710 20578 11740
rect 20478 11670 20508 11710
rect 20548 11670 20578 11710
rect 20478 11610 20578 11670
rect 20478 11570 20508 11610
rect 20548 11570 20578 11610
rect 20478 11540 20578 11570
rect 21458 11710 21558 11740
rect 21458 11670 21488 11710
rect 21528 11670 21558 11710
rect 21458 11610 21558 11670
rect 21458 11570 21488 11610
rect 21528 11570 21558 11610
rect 21458 11540 21558 11570
rect 21618 11710 21718 11740
rect 21618 11670 21648 11710
rect 21688 11670 21718 11710
rect 21618 11610 21718 11670
rect 21618 11570 21648 11610
rect 21688 11570 21718 11610
rect 21618 11540 21718 11570
rect 22598 11710 22698 11740
rect 22598 11670 22628 11710
rect 22668 11670 22698 11710
rect 22598 11610 22698 11670
rect 22598 11570 22628 11610
rect 22668 11570 22698 11610
rect 22598 11540 22698 11570
rect 23031 10733 23127 10767
rect 23387 10733 23483 10767
rect 23031 10671 23065 10733
rect 11538 10630 11618 10660
rect 11538 10590 11558 10630
rect 11598 10590 11618 10630
rect 11538 10530 11618 10590
rect 11538 10490 11558 10530
rect 11598 10490 11618 10530
rect 11538 10430 11618 10490
rect 11538 10390 11558 10430
rect 11598 10390 11618 10430
rect 11538 10330 11618 10390
rect 11538 10290 11558 10330
rect 11598 10290 11618 10330
rect 11538 10230 11618 10290
rect 11538 10190 11558 10230
rect 11598 10190 11618 10230
rect 11538 10130 11618 10190
rect 11538 10090 11558 10130
rect 11598 10090 11618 10130
rect 11538 10060 11618 10090
rect 14938 10630 15018 10660
rect 14938 10590 14958 10630
rect 14998 10590 15018 10630
rect 14938 10530 15018 10590
rect 14938 10490 14958 10530
rect 14998 10490 15018 10530
rect 14938 10430 15018 10490
rect 14938 10390 14958 10430
rect 14998 10390 15018 10430
rect 14938 10330 15018 10390
rect 14938 10290 14958 10330
rect 14998 10290 15018 10330
rect 14938 10230 15018 10290
rect 15398 10430 15478 10460
rect 15398 10390 15418 10430
rect 15458 10390 15478 10430
rect 15398 10330 15478 10390
rect 15398 10290 15418 10330
rect 15458 10290 15478 10330
rect 15398 10260 15478 10290
rect 16008 10430 16088 10460
rect 16008 10390 16028 10430
rect 16068 10390 16088 10430
rect 16008 10330 16088 10390
rect 16008 10290 16028 10330
rect 16068 10290 16088 10330
rect 16008 10260 16088 10290
rect 14938 10190 14958 10230
rect 14998 10190 15018 10230
rect 14938 10130 15018 10190
rect 14938 10090 14958 10130
rect 14998 10090 15018 10130
rect 14938 10060 15018 10090
rect 11548 9630 11628 9660
rect 11548 9590 11568 9630
rect 11608 9590 11628 9630
rect 11548 9530 11628 9590
rect 11548 9490 11568 9530
rect 11608 9490 11628 9530
rect 11548 9460 11628 9490
rect 13028 9630 13108 9660
rect 13028 9590 13048 9630
rect 13088 9590 13108 9630
rect 13028 9530 13108 9590
rect 13028 9490 13048 9530
rect 13088 9490 13108 9530
rect 13028 9460 13108 9490
rect 13448 9630 13528 9660
rect 13448 9590 13468 9630
rect 13508 9590 13528 9630
rect 13448 9530 13528 9590
rect 13448 9490 13468 9530
rect 13508 9490 13528 9530
rect 13448 9460 13528 9490
rect 14928 9630 15008 9660
rect 14928 9590 14948 9630
rect 14988 9590 15008 9630
rect 14928 9530 15008 9590
rect 14928 9490 14948 9530
rect 14988 9490 15008 9530
rect 14928 9460 15008 9490
rect 23449 10671 23483 10733
rect 23031 9519 23065 9581
rect 23449 9519 23483 9581
rect 23031 9485 23127 9519
rect 23387 9485 23483 9519
rect 13168 7640 13248 7670
rect 13168 7600 13188 7640
rect 13228 7600 13248 7640
rect 13168 7540 13248 7600
rect 13168 7500 13188 7540
rect 13228 7500 13248 7540
rect 13168 7440 13248 7500
rect 13168 7400 13188 7440
rect 13228 7400 13248 7440
rect 13168 7340 13248 7400
rect 13168 7300 13188 7340
rect 13228 7300 13248 7340
rect 13168 7270 13248 7300
rect 14068 7640 14148 7670
rect 14068 7600 14088 7640
rect 14128 7600 14148 7640
rect 14068 7540 14148 7600
rect 14068 7500 14088 7540
rect 14128 7500 14148 7540
rect 14068 7440 14148 7500
rect 14068 7400 14088 7440
rect 14128 7400 14148 7440
rect 14068 7340 14148 7400
rect 14068 7300 14088 7340
rect 14128 7300 14148 7340
rect 14068 7270 14148 7300
rect 14968 7640 15048 7670
rect 14968 7600 14988 7640
rect 15028 7600 15048 7640
rect 14968 7540 15048 7600
rect 14968 7500 14988 7540
rect 15028 7500 15048 7540
rect 14968 7440 15048 7500
rect 14968 7400 14988 7440
rect 15028 7400 15048 7440
rect 14968 7340 15048 7400
rect 14968 7300 14988 7340
rect 15028 7300 15048 7340
rect 14968 7270 15048 7300
rect 15368 7640 15448 7670
rect 15368 7600 15388 7640
rect 15428 7600 15448 7640
rect 15368 7540 15448 7600
rect 15368 7500 15388 7540
rect 15428 7500 15448 7540
rect 15368 7440 15448 7500
rect 15368 7400 15388 7440
rect 15428 7400 15448 7440
rect 15368 7340 15448 7400
rect 15368 7300 15388 7340
rect 15428 7300 15448 7340
rect 15368 7270 15448 7300
rect 15698 7640 15778 7670
rect 15698 7600 15718 7640
rect 15758 7600 15778 7640
rect 15698 7540 15778 7600
rect 15698 7500 15718 7540
rect 15758 7500 15778 7540
rect 15698 7440 15778 7500
rect 15698 7400 15718 7440
rect 15758 7400 15778 7440
rect 15698 7340 15778 7400
rect 15698 7300 15718 7340
rect 15758 7300 15778 7340
rect 15698 7270 15778 7300
rect 16028 7640 16108 7670
rect 16028 7600 16048 7640
rect 16088 7600 16108 7640
rect 16028 7540 16108 7600
rect 16028 7500 16048 7540
rect 16088 7500 16108 7540
rect 16028 7440 16108 7500
rect 16028 7400 16048 7440
rect 16088 7400 16108 7440
rect 16028 7340 16108 7400
rect 16028 7300 16048 7340
rect 16088 7300 16108 7340
rect 16028 7270 16108 7300
rect 16278 7640 16378 7670
rect 16278 7600 16308 7640
rect 16348 7600 16378 7640
rect 16278 7540 16378 7600
rect 16278 7500 16308 7540
rect 16348 7500 16378 7540
rect 16278 7440 16378 7500
rect 16278 7400 16308 7440
rect 16348 7400 16378 7440
rect 16278 7340 16378 7400
rect 16278 7300 16308 7340
rect 16348 7300 16378 7340
rect 16278 7270 16378 7300
rect 17058 7640 17158 7670
rect 17058 7600 17088 7640
rect 17128 7600 17158 7640
rect 17058 7540 17158 7600
rect 17058 7500 17088 7540
rect 17128 7500 17158 7540
rect 17058 7440 17158 7500
rect 17058 7400 17088 7440
rect 17128 7400 17158 7440
rect 17058 7340 17158 7400
rect 17058 7300 17088 7340
rect 17128 7300 17158 7340
rect 17058 7270 17158 7300
rect 19428 6910 19528 6940
rect 13168 6880 13248 6910
rect 13168 6840 13188 6880
rect 13228 6840 13248 6880
rect 13168 6780 13248 6840
rect 13168 6740 13188 6780
rect 13228 6740 13248 6780
rect 13168 6680 13248 6740
rect 13168 6640 13188 6680
rect 13228 6640 13248 6680
rect 13168 6580 13248 6640
rect 13168 6540 13188 6580
rect 13228 6540 13248 6580
rect 13168 6510 13248 6540
rect 14068 6880 14148 6910
rect 14068 6840 14088 6880
rect 14128 6840 14148 6880
rect 14068 6780 14148 6840
rect 14068 6740 14088 6780
rect 14128 6740 14148 6780
rect 14068 6680 14148 6740
rect 14068 6640 14088 6680
rect 14128 6640 14148 6680
rect 14068 6580 14148 6640
rect 14068 6540 14088 6580
rect 14128 6540 14148 6580
rect 14068 6510 14148 6540
rect 14968 6880 15048 6910
rect 14968 6840 14988 6880
rect 15028 6840 15048 6880
rect 14968 6780 15048 6840
rect 14968 6740 14988 6780
rect 15028 6740 15048 6780
rect 14968 6680 15048 6740
rect 14968 6640 14988 6680
rect 15028 6640 15048 6680
rect 14968 6580 15048 6640
rect 14968 6540 14988 6580
rect 15028 6540 15048 6580
rect 14968 6510 15048 6540
rect 15108 6900 15168 6910
rect 15108 6880 15188 6900
rect 15108 6840 15128 6880
rect 15168 6840 15188 6880
rect 15108 6780 15188 6840
rect 15108 6740 15128 6780
rect 15168 6740 15188 6780
rect 15108 6680 15188 6740
rect 15108 6640 15128 6680
rect 15168 6640 15188 6680
rect 15108 6580 15188 6640
rect 15108 6540 15128 6580
rect 15168 6540 15188 6580
rect 15108 6510 15188 6540
rect 15548 6880 15628 6910
rect 15548 6840 15568 6880
rect 15608 6840 15628 6880
rect 15548 6780 15628 6840
rect 15548 6740 15568 6780
rect 15608 6740 15628 6780
rect 15548 6680 15628 6740
rect 15548 6640 15568 6680
rect 15608 6640 15628 6680
rect 15548 6580 15628 6640
rect 15548 6540 15568 6580
rect 15608 6540 15628 6580
rect 15548 6510 15628 6540
rect 15878 6880 15958 6910
rect 15878 6840 15898 6880
rect 15938 6840 15958 6880
rect 15878 6780 15958 6840
rect 15878 6740 15898 6780
rect 15938 6740 15958 6780
rect 15878 6680 15958 6740
rect 15878 6640 15898 6680
rect 15938 6640 15958 6680
rect 15878 6580 15958 6640
rect 15878 6540 15898 6580
rect 15938 6540 15958 6580
rect 15878 6510 15958 6540
rect 16278 6880 16378 6910
rect 16278 6840 16308 6880
rect 16348 6840 16378 6880
rect 16278 6780 16378 6840
rect 16278 6740 16308 6780
rect 16348 6740 16378 6780
rect 16278 6680 16378 6740
rect 16278 6640 16308 6680
rect 16348 6640 16378 6680
rect 16278 6580 16378 6640
rect 16278 6540 16308 6580
rect 16348 6540 16378 6580
rect 16278 6510 16378 6540
rect 16668 6880 16768 6910
rect 16668 6840 16698 6880
rect 16738 6840 16768 6880
rect 16668 6780 16768 6840
rect 16668 6740 16698 6780
rect 16738 6740 16768 6780
rect 16668 6680 16768 6740
rect 16668 6640 16698 6680
rect 16738 6640 16768 6680
rect 16668 6580 16768 6640
rect 16668 6540 16698 6580
rect 16738 6540 16768 6580
rect 16668 6510 16768 6540
rect 17058 6880 17158 6910
rect 17058 6840 17088 6880
rect 17128 6840 17158 6880
rect 17058 6780 17158 6840
rect 17058 6740 17088 6780
rect 17128 6740 17158 6780
rect 17058 6680 17158 6740
rect 17058 6640 17088 6680
rect 17128 6640 17158 6680
rect 17058 6580 17158 6640
rect 17058 6540 17088 6580
rect 17128 6540 17158 6580
rect 17058 6510 17158 6540
rect 17738 6880 17838 6910
rect 17738 6840 17768 6880
rect 17808 6840 17838 6880
rect 17738 6780 17838 6840
rect 17738 6740 17768 6780
rect 17808 6740 17838 6780
rect 17738 6680 17838 6740
rect 17738 6640 17768 6680
rect 17808 6640 17838 6680
rect 17738 6580 17838 6640
rect 17738 6540 17768 6580
rect 17808 6540 17838 6580
rect 17738 6510 17838 6540
rect 19428 6870 19458 6910
rect 19498 6870 19528 6910
rect 19428 6810 19528 6870
rect 19428 6770 19458 6810
rect 19498 6770 19528 6810
rect 19428 6710 19528 6770
rect 19428 6670 19458 6710
rect 19498 6670 19528 6710
rect 19428 6610 19528 6670
rect 19428 6570 19458 6610
rect 19498 6570 19528 6610
rect 19428 6540 19528 6570
rect 20948 6910 21048 6940
rect 20948 6870 20978 6910
rect 21018 6870 21048 6910
rect 20948 6810 21048 6870
rect 20948 6770 20978 6810
rect 21018 6770 21048 6810
rect 20948 6710 21048 6770
rect 20948 6670 20978 6710
rect 21018 6670 21048 6710
rect 20948 6610 21048 6670
rect 20948 6570 20978 6610
rect 21018 6570 21048 6610
rect 20948 6540 21048 6570
rect 22468 6910 22568 6940
rect 22468 6870 22498 6910
rect 22538 6870 22568 6910
rect 22468 6810 22568 6870
rect 22468 6770 22498 6810
rect 22538 6770 22568 6810
rect 22468 6710 22568 6770
rect 22468 6670 22498 6710
rect 22538 6670 22568 6710
rect 22468 6610 22568 6670
rect 22468 6570 22498 6610
rect 22538 6570 22568 6610
rect 22468 6540 22568 6570
rect 23088 5490 24108 5530
rect 24268 5490 25148 5530
rect 25218 5490 25318 5530
rect 23088 5060 23128 5490
rect 25278 5060 25318 5490
rect 12778 3500 12858 3530
rect 12778 3460 12798 3500
rect 12838 3460 12858 3500
rect 12778 3430 12858 3460
rect 15148 3500 15228 3530
rect 15148 3460 15168 3500
rect 15208 3460 15228 3500
rect 15148 3430 15228 3460
rect 18018 3500 18098 3530
rect 18018 3460 18038 3500
rect 18078 3460 18098 3500
rect 18018 3430 18098 3460
rect 19318 3500 19398 3530
rect 19318 3460 19338 3500
rect 19378 3460 19398 3500
rect 19318 3430 19398 3460
rect 20618 3500 20698 3530
rect 20618 3460 20638 3500
rect 20678 3460 20698 3500
rect 20618 3430 20698 3460
rect 21918 3500 21998 3530
rect 21918 3460 21938 3500
rect 21978 3460 21998 3500
rect 21918 3430 21998 3460
rect 23088 3420 23128 4730
rect 25278 3420 25318 4730
rect 23088 3380 24108 3420
rect 24268 3380 25318 3420
<< psubdiffcont >>
rect 13258 19030 13298 19070
rect 13258 18950 13298 18990
rect 13258 18870 13298 18910
rect 11408 18718 11442 18752
rect 11498 18718 11532 18752
rect 11588 18718 11622 18752
rect 11678 18718 11712 18752
rect 11768 18718 11802 18752
rect 11858 18718 11892 18752
rect 11948 18718 11982 18752
rect 12038 18718 12072 18752
rect 12128 18718 12162 18752
rect 12218 18718 12252 18752
rect 12308 18718 12342 18752
rect 12398 18718 12432 18752
rect 11307 18634 11341 18668
rect 12494 18634 12528 18668
rect 11307 18544 11341 18578
rect 11307 18454 11341 18488
rect 11307 18364 11341 18398
rect 11307 18274 11341 18308
rect 11307 18184 11341 18218
rect 11307 18094 11341 18128
rect 11307 18004 11341 18038
rect 11307 17914 11341 17948
rect 11307 17824 11341 17858
rect 11307 17734 11341 17768
rect 11307 17644 11341 17678
rect 12494 18544 12528 18578
rect 12494 18454 12528 18488
rect 12494 18364 12528 18398
rect 12494 18274 12528 18308
rect 12494 18184 12528 18218
rect 12494 18094 12528 18128
rect 12494 18004 12528 18038
rect 12494 17914 12528 17948
rect 12494 17824 12528 17858
rect 12494 17734 12528 17768
rect 12494 17644 12528 17678
rect 11307 17554 11341 17588
rect 11408 17531 11442 17565
rect 11498 17531 11532 17565
rect 11588 17531 11622 17565
rect 11678 17531 11712 17565
rect 11768 17531 11802 17565
rect 11858 17531 11892 17565
rect 11948 17531 11982 17565
rect 12038 17531 12072 17565
rect 12128 17531 12162 17565
rect 12218 17531 12252 17565
rect 12308 17531 12342 17565
rect 12398 17531 12432 17565
rect 12494 17554 12528 17588
rect 12768 18718 12802 18752
rect 12858 18718 12892 18752
rect 12948 18718 12982 18752
rect 13038 18718 13072 18752
rect 13128 18718 13162 18752
rect 13218 18718 13252 18752
rect 13308 18718 13342 18752
rect 13398 18718 13432 18752
rect 13488 18718 13522 18752
rect 13578 18718 13612 18752
rect 13668 18718 13702 18752
rect 13758 18718 13792 18752
rect 12667 18634 12701 18668
rect 13854 18634 13888 18668
rect 12667 18544 12701 18578
rect 12667 18454 12701 18488
rect 12667 18364 12701 18398
rect 12667 18274 12701 18308
rect 12667 18184 12701 18218
rect 12667 18094 12701 18128
rect 12667 18004 12701 18038
rect 12667 17914 12701 17948
rect 12667 17824 12701 17858
rect 12667 17734 12701 17768
rect 12667 17644 12701 17678
rect 13854 18544 13888 18578
rect 13854 18454 13888 18488
rect 13854 18364 13888 18398
rect 13854 18274 13888 18308
rect 13854 18184 13888 18218
rect 13854 18094 13888 18128
rect 13854 18004 13888 18038
rect 13854 17914 13888 17948
rect 13854 17824 13888 17858
rect 13854 17734 13888 17768
rect 13854 17644 13888 17678
rect 12667 17554 12701 17588
rect 12768 17531 12802 17565
rect 12858 17531 12892 17565
rect 12948 17531 12982 17565
rect 13038 17531 13072 17565
rect 13128 17531 13162 17565
rect 13218 17531 13252 17565
rect 13308 17531 13342 17565
rect 13398 17531 13432 17565
rect 13488 17531 13522 17565
rect 13578 17531 13612 17565
rect 13668 17531 13702 17565
rect 13758 17531 13792 17565
rect 13854 17554 13888 17588
rect 14128 18718 14162 18752
rect 14218 18718 14252 18752
rect 14308 18718 14342 18752
rect 14398 18718 14432 18752
rect 14488 18718 14522 18752
rect 14578 18718 14612 18752
rect 14668 18718 14702 18752
rect 14758 18718 14792 18752
rect 14848 18718 14882 18752
rect 14938 18718 14972 18752
rect 15028 18718 15062 18752
rect 15118 18718 15152 18752
rect 14027 18634 14061 18668
rect 15214 18634 15248 18668
rect 14027 18544 14061 18578
rect 14027 18454 14061 18488
rect 14027 18364 14061 18398
rect 14027 18274 14061 18308
rect 14027 18184 14061 18218
rect 14027 18094 14061 18128
rect 14027 18004 14061 18038
rect 14027 17914 14061 17948
rect 14027 17824 14061 17858
rect 14027 17734 14061 17768
rect 14027 17644 14061 17678
rect 15214 18544 15248 18578
rect 15214 18454 15248 18488
rect 15214 18364 15248 18398
rect 15214 18274 15248 18308
rect 15214 18184 15248 18218
rect 15214 18094 15248 18128
rect 15214 18004 15248 18038
rect 15214 17914 15248 17948
rect 15214 17824 15248 17858
rect 15214 17734 15248 17768
rect 15214 17644 15248 17678
rect 14027 17554 14061 17588
rect 14128 17531 14162 17565
rect 14218 17531 14252 17565
rect 14308 17531 14342 17565
rect 14398 17531 14432 17565
rect 14488 17531 14522 17565
rect 14578 17531 14612 17565
rect 14668 17531 14702 17565
rect 14758 17531 14792 17565
rect 14848 17531 14882 17565
rect 14938 17531 14972 17565
rect 15028 17531 15062 17565
rect 15118 17531 15152 17565
rect 15214 17554 15248 17588
rect 11408 17358 11442 17392
rect 11498 17358 11532 17392
rect 11588 17358 11622 17392
rect 11678 17358 11712 17392
rect 11768 17358 11802 17392
rect 11858 17358 11892 17392
rect 11948 17358 11982 17392
rect 12038 17358 12072 17392
rect 12128 17358 12162 17392
rect 12218 17358 12252 17392
rect 12308 17358 12342 17392
rect 12398 17358 12432 17392
rect 11307 17274 11341 17308
rect 12494 17274 12528 17308
rect 11307 17184 11341 17218
rect 11307 17094 11341 17128
rect 11307 17004 11341 17038
rect 11307 16914 11341 16948
rect 11307 16824 11341 16858
rect 11307 16734 11341 16768
rect 11307 16644 11341 16678
rect 11307 16554 11341 16588
rect 11307 16464 11341 16498
rect 11307 16374 11341 16408
rect 11307 16284 11341 16318
rect 12494 17184 12528 17218
rect 12494 17094 12528 17128
rect 12494 17004 12528 17038
rect 12494 16914 12528 16948
rect 12494 16824 12528 16858
rect 12494 16734 12528 16768
rect 12494 16644 12528 16678
rect 12494 16554 12528 16588
rect 12494 16464 12528 16498
rect 12494 16374 12528 16408
rect 12494 16284 12528 16318
rect 11307 16194 11341 16228
rect 11408 16171 11442 16205
rect 11498 16171 11532 16205
rect 11588 16171 11622 16205
rect 11678 16171 11712 16205
rect 11768 16171 11802 16205
rect 11858 16171 11892 16205
rect 11948 16171 11982 16205
rect 12038 16171 12072 16205
rect 12128 16171 12162 16205
rect 12218 16171 12252 16205
rect 12308 16171 12342 16205
rect 12398 16171 12432 16205
rect 12494 16194 12528 16228
rect 12768 17358 12802 17392
rect 12858 17358 12892 17392
rect 12948 17358 12982 17392
rect 13038 17358 13072 17392
rect 13128 17358 13162 17392
rect 13218 17358 13252 17392
rect 13308 17358 13342 17392
rect 13398 17358 13432 17392
rect 13488 17358 13522 17392
rect 13578 17358 13612 17392
rect 13668 17358 13702 17392
rect 13758 17358 13792 17392
rect 12667 17274 12701 17308
rect 13854 17274 13888 17308
rect 12667 17184 12701 17218
rect 12667 17094 12701 17128
rect 12667 17004 12701 17038
rect 12667 16914 12701 16948
rect 12667 16824 12701 16858
rect 12667 16734 12701 16768
rect 12667 16644 12701 16678
rect 12667 16554 12701 16588
rect 12667 16464 12701 16498
rect 12667 16374 12701 16408
rect 12667 16284 12701 16318
rect 13854 17184 13888 17218
rect 13854 17094 13888 17128
rect 13854 17004 13888 17038
rect 13854 16914 13888 16948
rect 13854 16824 13888 16858
rect 13854 16734 13888 16768
rect 13854 16644 13888 16678
rect 13854 16554 13888 16588
rect 13854 16464 13888 16498
rect 13854 16374 13888 16408
rect 13854 16284 13888 16318
rect 12667 16194 12701 16228
rect 12768 16171 12802 16205
rect 12858 16171 12892 16205
rect 12948 16171 12982 16205
rect 13038 16171 13072 16205
rect 13128 16171 13162 16205
rect 13218 16171 13252 16205
rect 13308 16171 13342 16205
rect 13398 16171 13432 16205
rect 13488 16171 13522 16205
rect 13578 16171 13612 16205
rect 13668 16171 13702 16205
rect 13758 16171 13792 16205
rect 13854 16194 13888 16228
rect 14128 17358 14162 17392
rect 14218 17358 14252 17392
rect 14308 17358 14342 17392
rect 14398 17358 14432 17392
rect 14488 17358 14522 17392
rect 14578 17358 14612 17392
rect 14668 17358 14702 17392
rect 14758 17358 14792 17392
rect 14848 17358 14882 17392
rect 14938 17358 14972 17392
rect 15028 17358 15062 17392
rect 15118 17358 15152 17392
rect 14027 17274 14061 17308
rect 15214 17274 15248 17308
rect 14027 17184 14061 17218
rect 14027 17094 14061 17128
rect 14027 17004 14061 17038
rect 14027 16914 14061 16948
rect 14027 16824 14061 16858
rect 14027 16734 14061 16768
rect 14027 16644 14061 16678
rect 14027 16554 14061 16588
rect 14027 16464 14061 16498
rect 14027 16374 14061 16408
rect 14027 16284 14061 16318
rect 15214 17184 15248 17218
rect 15214 17094 15248 17128
rect 15214 17004 15248 17038
rect 15214 16914 15248 16948
rect 15214 16824 15248 16858
rect 15214 16734 15248 16768
rect 15214 16644 15248 16678
rect 15214 16554 15248 16588
rect 15214 16464 15248 16498
rect 15214 16374 15248 16408
rect 15214 16284 15248 16318
rect 14027 16194 14061 16228
rect 14128 16171 14162 16205
rect 14218 16171 14252 16205
rect 14308 16171 14342 16205
rect 14398 16171 14432 16205
rect 14488 16171 14522 16205
rect 14578 16171 14612 16205
rect 14668 16171 14702 16205
rect 14758 16171 14792 16205
rect 14848 16171 14882 16205
rect 14938 16171 14972 16205
rect 15028 16171 15062 16205
rect 15118 16171 15152 16205
rect 15214 16194 15248 16228
rect 11408 15998 11442 16032
rect 11498 15998 11532 16032
rect 11588 15998 11622 16032
rect 11678 15998 11712 16032
rect 11768 15998 11802 16032
rect 11858 15998 11892 16032
rect 11948 15998 11982 16032
rect 12038 15998 12072 16032
rect 12128 15998 12162 16032
rect 12218 15998 12252 16032
rect 12308 15998 12342 16032
rect 12398 15998 12432 16032
rect 11307 15914 11341 15948
rect 12494 15914 12528 15948
rect 11307 15824 11341 15858
rect 11307 15734 11341 15768
rect 11307 15644 11341 15678
rect 11307 15554 11341 15588
rect 11307 15464 11341 15498
rect 11307 15374 11341 15408
rect 11307 15284 11341 15318
rect 11307 15194 11341 15228
rect 11307 15104 11341 15138
rect 11307 15014 11341 15048
rect 11307 14924 11341 14958
rect 12494 15824 12528 15858
rect 12494 15734 12528 15768
rect 12494 15644 12528 15678
rect 12494 15554 12528 15588
rect 12494 15464 12528 15498
rect 12494 15374 12528 15408
rect 12494 15284 12528 15318
rect 12494 15194 12528 15228
rect 12494 15104 12528 15138
rect 12494 15014 12528 15048
rect 12494 14924 12528 14958
rect 11307 14834 11341 14868
rect 11408 14811 11442 14845
rect 11498 14811 11532 14845
rect 11588 14811 11622 14845
rect 11678 14811 11712 14845
rect 11768 14811 11802 14845
rect 11858 14811 11892 14845
rect 11948 14811 11982 14845
rect 12038 14811 12072 14845
rect 12128 14811 12162 14845
rect 12218 14811 12252 14845
rect 12308 14811 12342 14845
rect 12398 14811 12432 14845
rect 12494 14834 12528 14868
rect 12768 15998 12802 16032
rect 12858 15998 12892 16032
rect 12948 15998 12982 16032
rect 13038 15998 13072 16032
rect 13128 15998 13162 16032
rect 13218 15998 13252 16032
rect 13308 15998 13342 16032
rect 13398 15998 13432 16032
rect 13488 15998 13522 16032
rect 13578 15998 13612 16032
rect 13668 15998 13702 16032
rect 13758 15998 13792 16032
rect 12667 15914 12701 15948
rect 13854 15914 13888 15948
rect 12667 15824 12701 15858
rect 12667 15734 12701 15768
rect 12667 15644 12701 15678
rect 12667 15554 12701 15588
rect 12667 15464 12701 15498
rect 12667 15374 12701 15408
rect 12667 15284 12701 15318
rect 12667 15194 12701 15228
rect 12667 15104 12701 15138
rect 12667 15014 12701 15048
rect 12667 14924 12701 14958
rect 13854 15824 13888 15858
rect 13854 15734 13888 15768
rect 13854 15644 13888 15678
rect 13854 15554 13888 15588
rect 13854 15464 13888 15498
rect 13854 15374 13888 15408
rect 13854 15284 13888 15318
rect 13854 15194 13888 15228
rect 13854 15104 13888 15138
rect 13854 15014 13888 15048
rect 13854 14924 13888 14958
rect 12667 14834 12701 14868
rect 12768 14811 12802 14845
rect 12858 14811 12892 14845
rect 12948 14811 12982 14845
rect 13038 14811 13072 14845
rect 13128 14811 13162 14845
rect 13218 14811 13252 14845
rect 13308 14811 13342 14845
rect 13398 14811 13432 14845
rect 13488 14811 13522 14845
rect 13578 14811 13612 14845
rect 13668 14811 13702 14845
rect 13758 14811 13792 14845
rect 13854 14834 13888 14868
rect 14128 15998 14162 16032
rect 14218 15998 14252 16032
rect 14308 15998 14342 16032
rect 14398 15998 14432 16032
rect 14488 15998 14522 16032
rect 14578 15998 14612 16032
rect 14668 15998 14702 16032
rect 14758 15998 14792 16032
rect 14848 15998 14882 16032
rect 14938 15998 14972 16032
rect 15028 15998 15062 16032
rect 15118 15998 15152 16032
rect 14027 15914 14061 15948
rect 15214 15914 15248 15948
rect 14027 15824 14061 15858
rect 14027 15734 14061 15768
rect 14027 15644 14061 15678
rect 14027 15554 14061 15588
rect 14027 15464 14061 15498
rect 14027 15374 14061 15408
rect 14027 15284 14061 15318
rect 14027 15194 14061 15228
rect 14027 15104 14061 15138
rect 14027 15014 14061 15048
rect 14027 14924 14061 14958
rect 15214 15824 15248 15858
rect 15214 15734 15248 15768
rect 15214 15644 15248 15678
rect 15214 15554 15248 15588
rect 15214 15464 15248 15498
rect 15214 15374 15248 15408
rect 15214 15284 15248 15318
rect 15214 15194 15248 15228
rect 15214 15104 15248 15138
rect 15214 15014 15248 15048
rect 15214 14924 15248 14958
rect 14027 14834 14061 14868
rect 14128 14811 14162 14845
rect 14218 14811 14252 14845
rect 14308 14811 14342 14845
rect 14398 14811 14432 14845
rect 14488 14811 14522 14845
rect 14578 14811 14612 14845
rect 14668 14811 14702 14845
rect 14758 14811 14792 14845
rect 14848 14811 14882 14845
rect 14938 14811 14972 14845
rect 15028 14811 15062 14845
rect 15118 14811 15152 14845
rect 15214 14834 15248 14868
rect 15418 14210 15458 14250
rect 15418 14110 15458 14150
rect 11918 13600 11958 13640
rect 11918 13500 11958 13540
rect 11918 13400 11958 13440
rect 11918 13300 11958 13340
rect 11918 13200 11958 13240
rect 14598 13600 14638 13640
rect 14598 13500 14638 13540
rect 14598 13400 14638 13440
rect 14598 13300 14638 13340
rect 14598 13200 14638 13240
rect 12818 12680 12858 12720
rect 12818 12600 12858 12640
rect 12818 12520 12858 12560
rect 13698 12680 13738 12720
rect 13698 12600 13738 12640
rect 13698 12520 13738 12560
rect 19368 10990 19408 11030
rect 20348 10990 20388 11030
rect 21648 10990 21688 11030
rect 22628 10990 22668 11030
rect 19318 10440 19358 10490
rect 19318 10300 19358 10350
rect 21518 10440 21558 10490
rect 21518 10300 21558 10350
rect 13188 8020 13228 8060
rect 13188 7920 13228 7960
rect 14088 8020 14128 8060
rect 14088 7920 14128 7960
rect 14988 8020 15028 8060
rect 14988 7920 15028 7960
rect 15388 8020 15428 8060
rect 15388 7920 15428 7960
rect 15718 8020 15758 8060
rect 15718 7920 15758 7960
rect 16048 8020 16088 8060
rect 16048 7920 16088 7960
rect 16308 8020 16348 8060
rect 16308 7920 16348 7960
rect 17088 8020 17128 8060
rect 17088 7920 17128 7960
rect 17768 8020 17808 8060
rect 17768 7920 17808 7960
rect 19258 7970 19298 8010
rect 19258 7870 19298 7910
rect 19258 7770 19298 7810
rect 19258 7670 19298 7710
rect 20338 7970 20378 8010
rect 20338 7870 20378 7910
rect 20338 7770 20378 7810
rect 20338 7670 20378 7710
rect 21418 7970 21458 8010
rect 21418 7870 21458 7910
rect 21418 7770 21458 7810
rect 21418 7670 21458 7710
rect 22498 7970 22538 8010
rect 22498 7870 22538 7910
rect 22498 7770 22538 7810
rect 22498 7670 22538 7710
rect 13188 6220 13228 6260
rect 13188 6120 13228 6160
rect 14088 6220 14128 6260
rect 14088 6120 14128 6160
rect 14988 6220 15028 6260
rect 14988 6120 15028 6160
rect 15128 6220 15168 6260
rect 15128 6120 15168 6160
rect 15568 6220 15608 6260
rect 15568 6120 15608 6160
rect 15898 6220 15938 6260
rect 15898 6120 15938 6160
rect 16318 6220 16358 6260
rect 16318 6120 16358 6160
rect 16708 6220 16748 6260
rect 16708 6120 16748 6160
rect 17098 6220 17138 6260
rect 17098 6120 17138 6160
rect 15698 3140 15738 3180
rect 17148 3140 17188 3180
rect 24228 3180 24368 3220
rect 18938 3050 18978 3090
rect 20238 3050 20278 3090
rect 21538 3050 21578 3090
rect 23088 2450 23128 2660
rect 25088 2450 25128 2660
rect 24228 1880 24368 1920
<< nsubdiffcont >>
rect 14947 19663 17369 19697
rect 14851 19341 14885 19601
rect 17431 19341 17465 19601
rect 14947 19245 17369 19279
rect 8357 18563 8617 18597
rect 8261 17173 8295 18501
rect 8679 17173 8713 18501
rect 8357 17077 8617 17111
rect 9144 18566 9736 18600
rect 9048 16774 9082 18504
rect 9798 16774 9832 18504
rect 9144 16678 9736 16712
rect 10257 18563 10849 18597
rect 10161 16243 10195 18501
rect 10911 16243 10945 18501
rect 11548 18568 11582 18602
rect 11638 18568 11672 18602
rect 11728 18568 11762 18602
rect 11818 18568 11852 18602
rect 11908 18568 11942 18602
rect 11998 18568 12032 18602
rect 12088 18568 12122 18602
rect 12178 18568 12212 18602
rect 12268 18568 12302 18602
rect 11456 18474 11490 18508
rect 11456 18384 11490 18418
rect 11456 18294 11490 18328
rect 11456 18204 11490 18238
rect 11456 18114 11490 18148
rect 11456 18024 11490 18058
rect 11456 17934 11490 17968
rect 11456 17844 11490 17878
rect 12346 18455 12380 18489
rect 12346 18365 12380 18399
rect 12346 18275 12380 18309
rect 12346 18185 12380 18219
rect 12346 18095 12380 18129
rect 12346 18005 12380 18039
rect 12346 17915 12380 17949
rect 12346 17825 12380 17859
rect 11456 17754 11490 17788
rect 12346 17735 12380 17769
rect 11514 17678 11548 17712
rect 11604 17678 11638 17712
rect 11694 17678 11728 17712
rect 11784 17678 11818 17712
rect 11874 17678 11908 17712
rect 11964 17678 11998 17712
rect 12054 17678 12088 17712
rect 12144 17678 12178 17712
rect 12234 17678 12268 17712
rect 12908 18568 12942 18602
rect 12998 18568 13032 18602
rect 13088 18568 13122 18602
rect 13178 18568 13212 18602
rect 13268 18568 13302 18602
rect 13358 18568 13392 18602
rect 13448 18568 13482 18602
rect 13538 18568 13572 18602
rect 13628 18568 13662 18602
rect 12816 18474 12850 18508
rect 12816 18384 12850 18418
rect 12816 18294 12850 18328
rect 12816 18204 12850 18238
rect 12816 18114 12850 18148
rect 12816 18024 12850 18058
rect 12816 17934 12850 17968
rect 12816 17844 12850 17878
rect 13706 18455 13740 18489
rect 13706 18365 13740 18399
rect 13706 18275 13740 18309
rect 13706 18185 13740 18219
rect 13706 18095 13740 18129
rect 13706 18005 13740 18039
rect 13706 17915 13740 17949
rect 13706 17825 13740 17859
rect 12816 17754 12850 17788
rect 13706 17735 13740 17769
rect 12874 17678 12908 17712
rect 12964 17678 12998 17712
rect 13054 17678 13088 17712
rect 13144 17678 13178 17712
rect 13234 17678 13268 17712
rect 13324 17678 13358 17712
rect 13414 17678 13448 17712
rect 13504 17678 13538 17712
rect 13594 17678 13628 17712
rect 14268 18568 14302 18602
rect 14358 18568 14392 18602
rect 14448 18568 14482 18602
rect 14538 18568 14572 18602
rect 14628 18568 14662 18602
rect 14718 18568 14752 18602
rect 14808 18568 14842 18602
rect 14898 18568 14932 18602
rect 14988 18568 15022 18602
rect 14176 18474 14210 18508
rect 14176 18384 14210 18418
rect 14176 18294 14210 18328
rect 14176 18204 14210 18238
rect 14176 18114 14210 18148
rect 14176 18024 14210 18058
rect 14176 17934 14210 17968
rect 14176 17844 14210 17878
rect 15066 18455 15100 18489
rect 15066 18365 15100 18399
rect 15066 18275 15100 18309
rect 15066 18185 15100 18219
rect 15066 18095 15100 18129
rect 15066 18005 15100 18039
rect 15066 17915 15100 17949
rect 15066 17825 15100 17859
rect 14176 17754 14210 17788
rect 15066 17735 15100 17769
rect 14234 17678 14268 17712
rect 14324 17678 14358 17712
rect 14414 17678 14448 17712
rect 14504 17678 14538 17712
rect 14594 17678 14628 17712
rect 14684 17678 14718 17712
rect 14774 17678 14808 17712
rect 14864 17678 14898 17712
rect 14954 17678 14988 17712
rect 15577 18563 16169 18597
rect 10257 16147 10849 16181
rect 11548 17208 11582 17242
rect 11638 17208 11672 17242
rect 11728 17208 11762 17242
rect 11818 17208 11852 17242
rect 11908 17208 11942 17242
rect 11998 17208 12032 17242
rect 12088 17208 12122 17242
rect 12178 17208 12212 17242
rect 12268 17208 12302 17242
rect 11456 17114 11490 17148
rect 11456 17024 11490 17058
rect 11456 16934 11490 16968
rect 11456 16844 11490 16878
rect 11456 16754 11490 16788
rect 11456 16664 11490 16698
rect 11456 16574 11490 16608
rect 11456 16484 11490 16518
rect 12346 17095 12380 17129
rect 12346 17005 12380 17039
rect 12346 16915 12380 16949
rect 12346 16825 12380 16859
rect 12346 16735 12380 16769
rect 12346 16645 12380 16679
rect 12346 16555 12380 16589
rect 12346 16465 12380 16499
rect 11456 16394 11490 16428
rect 12346 16375 12380 16409
rect 11514 16318 11548 16352
rect 11604 16318 11638 16352
rect 11694 16318 11728 16352
rect 11784 16318 11818 16352
rect 11874 16318 11908 16352
rect 11964 16318 11998 16352
rect 12054 16318 12088 16352
rect 12144 16318 12178 16352
rect 12234 16318 12268 16352
rect 12908 17208 12942 17242
rect 12998 17208 13032 17242
rect 13088 17208 13122 17242
rect 13178 17208 13212 17242
rect 13268 17208 13302 17242
rect 13358 17208 13392 17242
rect 13448 17208 13482 17242
rect 13538 17208 13572 17242
rect 13628 17208 13662 17242
rect 12816 17114 12850 17148
rect 12816 17024 12850 17058
rect 12816 16934 12850 16968
rect 12816 16844 12850 16878
rect 12816 16754 12850 16788
rect 12816 16664 12850 16698
rect 12816 16574 12850 16608
rect 12816 16484 12850 16518
rect 13706 17095 13740 17129
rect 13706 17005 13740 17039
rect 13706 16915 13740 16949
rect 13706 16825 13740 16859
rect 13706 16735 13740 16769
rect 13706 16645 13740 16679
rect 13706 16555 13740 16589
rect 13706 16465 13740 16499
rect 12816 16394 12850 16428
rect 13706 16375 13740 16409
rect 12874 16318 12908 16352
rect 12964 16318 12998 16352
rect 13054 16318 13088 16352
rect 13144 16318 13178 16352
rect 13234 16318 13268 16352
rect 13324 16318 13358 16352
rect 13414 16318 13448 16352
rect 13504 16318 13538 16352
rect 13594 16318 13628 16352
rect 14268 17208 14302 17242
rect 14358 17208 14392 17242
rect 14448 17208 14482 17242
rect 14538 17208 14572 17242
rect 14628 17208 14662 17242
rect 14718 17208 14752 17242
rect 14808 17208 14842 17242
rect 14898 17208 14932 17242
rect 14988 17208 15022 17242
rect 14176 17114 14210 17148
rect 14176 17024 14210 17058
rect 14176 16934 14210 16968
rect 14176 16844 14210 16878
rect 14176 16754 14210 16788
rect 14176 16664 14210 16698
rect 14176 16574 14210 16608
rect 14176 16484 14210 16518
rect 15066 17095 15100 17129
rect 15066 17005 15100 17039
rect 15066 16915 15100 16949
rect 15066 16825 15100 16859
rect 15066 16735 15100 16769
rect 15066 16645 15100 16679
rect 15066 16555 15100 16589
rect 15066 16465 15100 16499
rect 14176 16394 14210 16428
rect 15066 16375 15100 16409
rect 14234 16318 14268 16352
rect 14324 16318 14358 16352
rect 14414 16318 14448 16352
rect 14504 16318 14538 16352
rect 14594 16318 14628 16352
rect 14684 16318 14718 16352
rect 14774 16318 14808 16352
rect 14864 16318 14898 16352
rect 14954 16318 14988 16352
rect 15481 16243 15515 18501
rect 16231 16243 16265 18501
rect 16690 18560 16950 18594
rect 16594 17380 16628 18498
rect 17012 17380 17046 18498
rect 16690 17284 16950 17318
rect 17477 18563 17737 18597
rect 17381 17173 17415 18501
rect 17799 17173 17833 18501
rect 17477 17077 17737 17111
rect 15577 16147 16169 16181
rect 11548 15848 11582 15882
rect 11638 15848 11672 15882
rect 11728 15848 11762 15882
rect 11818 15848 11852 15882
rect 11908 15848 11942 15882
rect 11998 15848 12032 15882
rect 12088 15848 12122 15882
rect 12178 15848 12212 15882
rect 12268 15848 12302 15882
rect 11456 15754 11490 15788
rect 11456 15664 11490 15698
rect 11456 15574 11490 15608
rect 11456 15484 11490 15518
rect 11456 15394 11490 15428
rect 11456 15304 11490 15338
rect 11456 15214 11490 15248
rect 11456 15124 11490 15158
rect 12346 15735 12380 15769
rect 12346 15645 12380 15679
rect 12346 15555 12380 15589
rect 12346 15465 12380 15499
rect 12346 15375 12380 15409
rect 12346 15285 12380 15319
rect 12346 15195 12380 15229
rect 12346 15105 12380 15139
rect 11456 15034 11490 15068
rect 12346 15015 12380 15049
rect 11514 14958 11548 14992
rect 11604 14958 11638 14992
rect 11694 14958 11728 14992
rect 11784 14958 11818 14992
rect 11874 14958 11908 14992
rect 11964 14958 11998 14992
rect 12054 14958 12088 14992
rect 12144 14958 12178 14992
rect 12234 14958 12268 14992
rect 12908 15848 12942 15882
rect 12998 15848 13032 15882
rect 13088 15848 13122 15882
rect 13178 15848 13212 15882
rect 13268 15848 13302 15882
rect 13358 15848 13392 15882
rect 13448 15848 13482 15882
rect 13538 15848 13572 15882
rect 13628 15848 13662 15882
rect 12816 15754 12850 15788
rect 12816 15664 12850 15698
rect 12816 15574 12850 15608
rect 12816 15484 12850 15518
rect 12816 15394 12850 15428
rect 12816 15304 12850 15338
rect 12816 15214 12850 15248
rect 12816 15124 12850 15158
rect 13706 15735 13740 15769
rect 13706 15645 13740 15679
rect 13706 15555 13740 15589
rect 13706 15465 13740 15499
rect 13706 15375 13740 15409
rect 13706 15285 13740 15319
rect 13706 15195 13740 15229
rect 13706 15105 13740 15139
rect 12816 15034 12850 15068
rect 13706 15015 13740 15049
rect 12874 14958 12908 14992
rect 12964 14958 12998 14992
rect 13054 14958 13088 14992
rect 13144 14958 13178 14992
rect 13234 14958 13268 14992
rect 13324 14958 13358 14992
rect 13414 14958 13448 14992
rect 13504 14958 13538 14992
rect 13594 14958 13628 14992
rect 14268 15848 14302 15882
rect 14358 15848 14392 15882
rect 14448 15848 14482 15882
rect 14538 15848 14572 15882
rect 14628 15848 14662 15882
rect 14718 15848 14752 15882
rect 14808 15848 14842 15882
rect 14898 15848 14932 15882
rect 14988 15848 15022 15882
rect 14176 15754 14210 15788
rect 14176 15664 14210 15698
rect 14176 15574 14210 15608
rect 14176 15484 14210 15518
rect 14176 15394 14210 15428
rect 14176 15304 14210 15338
rect 14176 15214 14210 15248
rect 14176 15124 14210 15158
rect 15066 15735 15100 15769
rect 15066 15645 15100 15679
rect 15066 15555 15100 15589
rect 15066 15465 15100 15499
rect 15066 15375 15100 15409
rect 15066 15285 15100 15319
rect 15066 15195 15100 15229
rect 15066 15105 15100 15139
rect 14176 15034 14210 15068
rect 15066 15015 15100 15049
rect 14234 14958 14268 14992
rect 14324 14958 14358 14992
rect 14414 14958 14448 14992
rect 14504 14958 14538 14992
rect 14594 14958 14628 14992
rect 14684 14958 14718 14992
rect 14774 14958 14808 14992
rect 14864 14958 14898 14992
rect 14954 14958 14988 14992
rect 23127 13253 23387 13287
rect 19438 12620 19478 12660
rect 19438 12520 19478 12560
rect 19438 12420 19478 12460
rect 19438 12320 19478 12360
rect 19438 12220 19478 12260
rect 21638 12620 21678 12660
rect 21638 12520 21678 12560
rect 21638 12420 21678 12460
rect 21638 12320 21678 12360
rect 21638 12220 21678 12260
rect 23031 12045 23065 13191
rect 23449 12045 23483 13191
rect 23127 11949 23387 11983
rect 10458 11750 10498 11790
rect 10458 11650 10498 11690
rect 13018 11750 13058 11790
rect 13018 11650 13058 11690
rect 13498 11750 13538 11790
rect 13498 11650 13538 11690
rect 16058 11750 16098 11790
rect 16058 11650 16098 11690
rect 20508 11670 20548 11710
rect 20508 11570 20548 11610
rect 21488 11670 21528 11710
rect 21488 11570 21528 11610
rect 21648 11670 21688 11710
rect 21648 11570 21688 11610
rect 22628 11670 22668 11710
rect 22628 11570 22668 11610
rect 23127 10733 23387 10767
rect 11558 10590 11598 10630
rect 11558 10490 11598 10530
rect 11558 10390 11598 10430
rect 11558 10290 11598 10330
rect 11558 10190 11598 10230
rect 11558 10090 11598 10130
rect 14958 10590 14998 10630
rect 14958 10490 14998 10530
rect 14958 10390 14998 10430
rect 14958 10290 14998 10330
rect 15418 10390 15458 10430
rect 15418 10290 15458 10330
rect 16028 10390 16068 10430
rect 16028 10290 16068 10330
rect 14958 10190 14998 10230
rect 14958 10090 14998 10130
rect 11568 9590 11608 9630
rect 11568 9490 11608 9530
rect 13048 9590 13088 9630
rect 13048 9490 13088 9530
rect 13468 9590 13508 9630
rect 13468 9490 13508 9530
rect 14948 9590 14988 9630
rect 14948 9490 14988 9530
rect 23031 9581 23065 10671
rect 23449 9581 23483 10671
rect 23127 9485 23387 9519
rect 13188 7600 13228 7640
rect 13188 7500 13228 7540
rect 13188 7400 13228 7440
rect 13188 7300 13228 7340
rect 14088 7600 14128 7640
rect 14088 7500 14128 7540
rect 14088 7400 14128 7440
rect 14088 7300 14128 7340
rect 14988 7600 15028 7640
rect 14988 7500 15028 7540
rect 14988 7400 15028 7440
rect 14988 7300 15028 7340
rect 15388 7600 15428 7640
rect 15388 7500 15428 7540
rect 15388 7400 15428 7440
rect 15388 7300 15428 7340
rect 15718 7600 15758 7640
rect 15718 7500 15758 7540
rect 15718 7400 15758 7440
rect 15718 7300 15758 7340
rect 16048 7600 16088 7640
rect 16048 7500 16088 7540
rect 16048 7400 16088 7440
rect 16048 7300 16088 7340
rect 16308 7600 16348 7640
rect 16308 7500 16348 7540
rect 16308 7400 16348 7440
rect 16308 7300 16348 7340
rect 17088 7600 17128 7640
rect 17088 7500 17128 7540
rect 17088 7400 17128 7440
rect 17088 7300 17128 7340
rect 13188 6840 13228 6880
rect 13188 6740 13228 6780
rect 13188 6640 13228 6680
rect 13188 6540 13228 6580
rect 14088 6840 14128 6880
rect 14088 6740 14128 6780
rect 14088 6640 14128 6680
rect 14088 6540 14128 6580
rect 14988 6840 15028 6880
rect 14988 6740 15028 6780
rect 14988 6640 15028 6680
rect 14988 6540 15028 6580
rect 15128 6840 15168 6880
rect 15128 6740 15168 6780
rect 15128 6640 15168 6680
rect 15128 6540 15168 6580
rect 15568 6840 15608 6880
rect 15568 6740 15608 6780
rect 15568 6640 15608 6680
rect 15568 6540 15608 6580
rect 15898 6840 15938 6880
rect 15898 6740 15938 6780
rect 15898 6640 15938 6680
rect 15898 6540 15938 6580
rect 16308 6840 16348 6880
rect 16308 6740 16348 6780
rect 16308 6640 16348 6680
rect 16308 6540 16348 6580
rect 16698 6840 16738 6880
rect 16698 6740 16738 6780
rect 16698 6640 16738 6680
rect 16698 6540 16738 6580
rect 17088 6840 17128 6880
rect 17088 6740 17128 6780
rect 17088 6640 17128 6680
rect 17088 6540 17128 6580
rect 17768 6840 17808 6880
rect 17768 6740 17808 6780
rect 17768 6640 17808 6680
rect 17768 6540 17808 6580
rect 19458 6870 19498 6910
rect 19458 6770 19498 6810
rect 19458 6670 19498 6710
rect 19458 6570 19498 6610
rect 20978 6870 21018 6910
rect 20978 6770 21018 6810
rect 20978 6670 21018 6710
rect 20978 6570 21018 6610
rect 22498 6870 22538 6910
rect 22498 6770 22538 6810
rect 22498 6670 22538 6710
rect 22498 6570 22538 6610
rect 24108 5490 24268 5530
rect 25148 5490 25218 5530
rect 23088 4730 23128 5060
rect 12798 3460 12838 3500
rect 15168 3460 15208 3500
rect 18038 3460 18078 3500
rect 19338 3460 19378 3500
rect 20638 3460 20678 3500
rect 21938 3460 21978 3500
rect 25278 4730 25318 5060
rect 24108 3380 24268 3420
<< poly >>
rect 11238 14280 13238 14310
rect 13318 14280 15318 14310
rect 11238 14050 13238 14080
rect 13318 14050 15318 14080
rect 11318 14030 11398 14050
rect 11318 13990 11338 14030
rect 11378 13990 11398 14030
rect 11318 13970 11398 13990
rect 11478 14030 11558 14050
rect 11478 13990 11498 14030
rect 11538 13990 11558 14030
rect 11478 13970 11558 13990
rect 11638 14030 11718 14050
rect 11638 13990 11658 14030
rect 11698 13990 11718 14030
rect 11638 13970 11718 13990
rect 11798 14030 11878 14050
rect 11798 13990 11818 14030
rect 11858 13990 11878 14030
rect 11798 13970 11878 13990
rect 11958 14030 12038 14050
rect 11958 13990 11978 14030
rect 12018 13990 12038 14030
rect 11958 13970 12038 13990
rect 12118 14030 12198 14050
rect 12118 13990 12138 14030
rect 12178 13990 12198 14030
rect 12118 13970 12198 13990
rect 12278 14030 12358 14050
rect 12278 13990 12298 14030
rect 12338 13990 12358 14030
rect 12278 13970 12358 13990
rect 12438 14030 12518 14050
rect 12438 13990 12458 14030
rect 12498 13990 12518 14030
rect 12438 13970 12518 13990
rect 12598 14030 12678 14050
rect 12598 13990 12618 14030
rect 12658 13990 12678 14030
rect 12598 13970 12678 13990
rect 12758 14030 12838 14050
rect 12758 13990 12778 14030
rect 12818 13990 12838 14030
rect 12758 13970 12838 13990
rect 12918 14030 12998 14050
rect 12918 13990 12938 14030
rect 12978 13990 12998 14030
rect 12918 13970 12998 13990
rect 13078 14030 13158 14050
rect 13078 13990 13098 14030
rect 13138 13990 13158 14030
rect 13078 13970 13158 13990
rect 13398 14030 13478 14050
rect 13398 13990 13418 14030
rect 13458 13990 13478 14030
rect 13398 13970 13478 13990
rect 13558 14030 13638 14050
rect 13558 13990 13578 14030
rect 13618 13990 13638 14030
rect 13558 13970 13638 13990
rect 13718 14030 13798 14050
rect 13718 13990 13738 14030
rect 13778 13990 13798 14030
rect 13718 13970 13798 13990
rect 13878 14030 13958 14050
rect 13878 13990 13898 14030
rect 13938 13990 13958 14030
rect 13878 13970 13958 13990
rect 14038 14030 14118 14050
rect 14038 13990 14058 14030
rect 14098 13990 14118 14030
rect 14038 13970 14118 13990
rect 14198 14030 14278 14050
rect 14198 13990 14218 14030
rect 14258 13990 14278 14030
rect 14198 13970 14278 13990
rect 14358 14030 14438 14050
rect 14358 13990 14378 14030
rect 14418 13990 14438 14030
rect 14358 13970 14438 13990
rect 14518 14030 14598 14050
rect 14518 13990 14538 14030
rect 14578 13990 14598 14030
rect 14518 13970 14598 13990
rect 14678 14030 14758 14050
rect 14678 13990 14698 14030
rect 14738 13990 14758 14030
rect 14678 13970 14758 13990
rect 14838 14030 14918 14050
rect 14838 13990 14858 14030
rect 14898 13990 14918 14030
rect 14838 13970 14918 13990
rect 14998 14030 15078 14050
rect 14998 13990 15018 14030
rect 15058 13990 15078 14030
rect 14998 13970 15078 13990
rect 15158 14030 15238 14050
rect 15158 13990 15178 14030
rect 15218 13990 15238 14030
rect 15158 13970 15238 13990
rect 10818 13670 11818 13700
rect 12058 13670 13058 13700
rect 13498 13670 14498 13700
rect 14738 13670 15738 13700
rect 10818 13140 11818 13170
rect 12058 13140 13058 13170
rect 13498 13140 14498 13170
rect 14738 13140 15738 13170
rect 10918 13120 10998 13140
rect 10918 13080 10938 13120
rect 10978 13080 10998 13120
rect 10918 13060 10998 13080
rect 11158 13120 11238 13140
rect 11158 13080 11178 13120
rect 11218 13080 11238 13120
rect 11158 13060 11238 13080
rect 11398 13120 11478 13140
rect 11398 13080 11418 13120
rect 11458 13080 11478 13120
rect 11398 13060 11478 13080
rect 11638 13120 11718 13140
rect 11638 13080 11658 13120
rect 11698 13080 11718 13120
rect 11638 13060 11718 13080
rect 12278 13120 12358 13140
rect 12278 13080 12298 13120
rect 12338 13080 12358 13120
rect 12278 13060 12358 13080
rect 12518 13120 12598 13140
rect 12518 13080 12538 13120
rect 12578 13080 12598 13120
rect 12518 13060 12598 13080
rect 12758 13120 12838 13140
rect 12758 13080 12778 13120
rect 12818 13080 12838 13120
rect 12758 13060 12838 13080
rect 13718 13120 13798 13140
rect 13718 13080 13738 13120
rect 13778 13080 13798 13120
rect 13718 13060 13798 13080
rect 13958 13120 14038 13140
rect 13958 13080 13978 13120
rect 14018 13080 14038 13120
rect 13958 13060 14038 13080
rect 14198 13120 14278 13140
rect 14198 13080 14218 13120
rect 14258 13080 14278 13120
rect 14198 13060 14278 13080
rect 14838 13120 14918 13140
rect 14838 13080 14858 13120
rect 14898 13080 14918 13120
rect 14838 13060 14918 13080
rect 15078 13120 15158 13140
rect 15078 13080 15098 13120
rect 15138 13080 15158 13120
rect 15078 13060 15158 13080
rect 15318 13120 15398 13140
rect 15318 13080 15338 13120
rect 15378 13080 15398 13120
rect 15318 13060 15398 13080
rect 15558 13120 15638 13140
rect 15558 13080 15578 13120
rect 15618 13080 15638 13120
rect 15558 13060 15638 13080
rect 20318 12780 20398 12800
rect 11429 12742 11487 12760
rect 11429 12708 11441 12742
rect 11475 12708 11487 12742
rect 11429 12690 11487 12708
rect 11789 12742 11847 12760
rect 11789 12708 11801 12742
rect 11835 12708 11847 12742
rect 11789 12690 11847 12708
rect 11909 12742 11967 12760
rect 11909 12708 11921 12742
rect 11955 12708 11967 12742
rect 11909 12690 11967 12708
rect 12269 12742 12327 12760
rect 12269 12708 12281 12742
rect 12315 12708 12327 12742
rect 12269 12690 12327 12708
rect 12389 12742 12447 12760
rect 12389 12708 12401 12742
rect 12435 12708 12447 12742
rect 12389 12690 12447 12708
rect 11438 12660 11478 12690
rect 11558 12660 11598 12690
rect 11678 12660 11718 12690
rect 11798 12660 11838 12690
rect 11918 12660 11958 12690
rect 12038 12660 12078 12690
rect 12158 12660 12198 12690
rect 12278 12660 12318 12690
rect 12398 12660 12438 12690
rect 12518 12660 12558 12690
rect 11438 12530 11478 12560
rect 11558 12530 11598 12560
rect 11530 12512 11598 12530
rect 11530 12478 11542 12512
rect 11576 12478 11598 12512
rect 11530 12460 11598 12478
rect 11678 12530 11718 12560
rect 11798 12530 11838 12560
rect 11918 12530 11958 12560
rect 12038 12530 12078 12560
rect 11678 12512 11746 12530
rect 11678 12478 11700 12512
rect 11734 12478 11746 12512
rect 11678 12460 11746 12478
rect 12012 12512 12078 12530
rect 12012 12478 12024 12512
rect 12058 12478 12078 12512
rect 12012 12460 12078 12478
rect 12158 12530 12198 12560
rect 12278 12530 12318 12560
rect 12398 12530 12438 12560
rect 12518 12530 12558 12560
rect 12158 12512 12224 12530
rect 12158 12478 12178 12512
rect 12212 12478 12224 12512
rect 12158 12460 12224 12478
rect 12490 12512 12558 12530
rect 12490 12478 12502 12512
rect 12536 12478 12558 12512
rect 14109 12742 14167 12760
rect 14109 12708 14121 12742
rect 14155 12708 14167 12742
rect 14109 12690 14167 12708
rect 14229 12742 14287 12760
rect 14229 12708 14241 12742
rect 14275 12708 14287 12742
rect 14229 12690 14287 12708
rect 14589 12742 14647 12760
rect 14589 12708 14601 12742
rect 14635 12708 14647 12742
rect 14589 12690 14647 12708
rect 14709 12742 14767 12760
rect 14709 12708 14721 12742
rect 14755 12708 14767 12742
rect 14709 12690 14767 12708
rect 15069 12742 15127 12760
rect 15069 12708 15081 12742
rect 15115 12708 15127 12742
rect 20318 12740 20338 12780
rect 20378 12740 20398 12780
rect 20718 12780 20798 12800
rect 20718 12740 20738 12780
rect 20778 12740 20798 12780
rect 15069 12690 15127 12708
rect 19608 12690 19708 12720
rect 19808 12710 21308 12740
rect 19808 12690 19908 12710
rect 20008 12690 20108 12710
rect 20208 12690 20308 12710
rect 20408 12690 20508 12710
rect 20608 12690 20708 12710
rect 20808 12690 20908 12710
rect 21008 12690 21108 12710
rect 21208 12690 21308 12710
rect 21408 12690 21508 12720
rect 13998 12660 14038 12690
rect 14118 12660 14158 12690
rect 14238 12660 14278 12690
rect 14358 12660 14398 12690
rect 14478 12660 14518 12690
rect 14598 12660 14638 12690
rect 14718 12660 14758 12690
rect 14838 12660 14878 12690
rect 14958 12660 14998 12690
rect 15078 12660 15118 12690
rect 13998 12530 14038 12560
rect 14118 12530 14158 12560
rect 14238 12530 14278 12560
rect 14358 12530 14398 12560
rect 13998 12512 14066 12530
rect 12490 12460 12558 12478
rect 13998 12478 14020 12512
rect 14054 12478 14066 12512
rect 13998 12460 14066 12478
rect 14332 12512 14398 12530
rect 14332 12478 14344 12512
rect 14378 12478 14398 12512
rect 14332 12460 14398 12478
rect 14478 12530 14518 12560
rect 14598 12530 14638 12560
rect 14718 12530 14758 12560
rect 14838 12530 14878 12560
rect 14478 12512 14544 12530
rect 14478 12478 14498 12512
rect 14532 12478 14544 12512
rect 14478 12460 14544 12478
rect 14810 12512 14878 12530
rect 14810 12478 14822 12512
rect 14856 12478 14878 12512
rect 14810 12460 14878 12478
rect 14958 12530 14998 12560
rect 15078 12530 15118 12560
rect 14958 12512 15026 12530
rect 14958 12478 14980 12512
rect 15014 12478 15026 12512
rect 14958 12460 15026 12478
rect 19608 12160 19708 12190
rect 19808 12160 19908 12190
rect 20008 12160 20108 12190
rect 20208 12160 20308 12190
rect 20408 12160 20508 12190
rect 20608 12160 20708 12190
rect 20808 12160 20908 12190
rect 21008 12160 21108 12190
rect 21208 12160 21308 12190
rect 21408 12160 21508 12190
rect 19518 12140 19708 12160
rect 19518 12100 19538 12140
rect 19578 12130 19708 12140
rect 21408 12140 21598 12160
rect 21408 12130 21538 12140
rect 19578 12100 19598 12130
rect 19518 12080 19598 12100
rect 21518 12100 21538 12130
rect 21578 12100 21598 12140
rect 21518 12080 21598 12100
rect 10708 11920 10768 11940
rect 10708 11880 10718 11920
rect 10758 11880 10768 11920
rect 10708 11860 10768 11880
rect 10878 11910 10958 11930
rect 10878 11870 10898 11910
rect 10938 11870 10958 11910
rect 11368 11910 11428 11930
rect 11368 11870 11378 11910
rect 11418 11870 11428 11910
rect 11598 11910 11678 11930
rect 11598 11870 11618 11910
rect 11658 11870 11678 11910
rect 12088 11910 12148 11930
rect 12088 11870 12098 11910
rect 12138 11870 12148 11910
rect 12318 11910 12398 11930
rect 12318 11870 12338 11910
rect 12378 11870 12398 11910
rect 12748 11910 12808 11930
rect 12748 11870 12758 11910
rect 12798 11870 12808 11910
rect 10598 11820 10638 11850
rect 10718 11820 10758 11860
rect 10838 11840 11238 11870
rect 10838 11820 10878 11840
rect 10958 11820 10998 11840
rect 11078 11820 11118 11840
rect 11198 11820 11238 11840
rect 11318 11840 11478 11870
rect 11318 11820 11358 11840
rect 11438 11820 11478 11840
rect 11558 11840 11958 11870
rect 11558 11820 11598 11840
rect 11678 11820 11718 11840
rect 11798 11820 11838 11840
rect 11918 11820 11958 11840
rect 12038 11840 12198 11870
rect 12038 11820 12078 11840
rect 12158 11820 12198 11840
rect 12278 11840 12678 11870
rect 12748 11850 12808 11870
rect 13748 11910 13808 11930
rect 13748 11870 13758 11910
rect 13798 11870 13808 11910
rect 14158 11910 14238 11930
rect 14158 11870 14178 11910
rect 14218 11870 14238 11910
rect 14408 11910 14468 11930
rect 14408 11870 14418 11910
rect 14458 11870 14468 11910
rect 14878 11910 14958 11930
rect 14878 11870 14898 11910
rect 14938 11870 14958 11910
rect 15128 11910 15188 11930
rect 15128 11870 15138 11910
rect 15178 11870 15188 11910
rect 15598 11910 15678 11930
rect 15598 11870 15618 11910
rect 15658 11870 15678 11910
rect 15788 11920 15848 11940
rect 15788 11880 15798 11920
rect 15838 11880 15848 11920
rect 13748 11850 13808 11870
rect 12278 11820 12318 11840
rect 12398 11820 12438 11840
rect 12518 11820 12558 11840
rect 12638 11820 12678 11840
rect 12758 11820 12798 11850
rect 12878 11820 12918 11850
rect 13638 11820 13678 11850
rect 13758 11820 13798 11850
rect 13878 11840 14278 11870
rect 13878 11820 13918 11840
rect 13998 11820 14038 11840
rect 14118 11820 14158 11840
rect 14238 11820 14278 11840
rect 14358 11840 14518 11870
rect 14358 11820 14398 11840
rect 14478 11820 14518 11840
rect 14598 11840 14998 11870
rect 14598 11820 14638 11840
rect 14718 11820 14758 11840
rect 14838 11820 14878 11840
rect 14958 11820 14998 11840
rect 15078 11840 15238 11870
rect 15078 11820 15118 11840
rect 15198 11820 15238 11840
rect 15318 11840 15718 11870
rect 15788 11860 15848 11880
rect 15318 11820 15358 11840
rect 15438 11820 15478 11840
rect 15558 11820 15598 11840
rect 15678 11820 15718 11840
rect 15798 11820 15838 11860
rect 15918 11820 15958 11850
rect 19508 11830 19588 11850
rect 19508 11790 19528 11830
rect 19568 11790 19588 11830
rect 19508 11770 19588 11790
rect 20168 11830 20248 11850
rect 20168 11790 20188 11830
rect 20228 11790 20248 11830
rect 20168 11770 20248 11790
rect 20648 11830 20728 11850
rect 20648 11790 20668 11830
rect 20708 11790 20728 11830
rect 20648 11770 20728 11790
rect 21308 11830 21388 11850
rect 21308 11790 21328 11830
rect 21368 11790 21388 11830
rect 21308 11770 21388 11790
rect 21788 11830 21868 11850
rect 21788 11790 21808 11830
rect 21848 11790 21868 11830
rect 21788 11770 21868 11790
rect 22448 11830 22528 11850
rect 22448 11790 22468 11830
rect 22508 11790 22528 11830
rect 22448 11770 22528 11790
rect 19538 11740 19568 11770
rect 19668 11740 19698 11770
rect 19798 11740 19828 11770
rect 19928 11740 19958 11770
rect 20058 11740 20088 11770
rect 20188 11740 20218 11770
rect 20678 11740 20708 11770
rect 20808 11740 20838 11770
rect 20938 11740 20968 11770
rect 21068 11740 21098 11770
rect 21198 11740 21228 11770
rect 21328 11740 21358 11770
rect 21818 11740 21848 11770
rect 21948 11740 21978 11770
rect 22078 11740 22108 11770
rect 22208 11740 22238 11770
rect 22338 11740 22368 11770
rect 22468 11740 22498 11770
rect 10598 11590 10638 11620
rect 10718 11590 10758 11620
rect 10838 11590 10878 11620
rect 10958 11590 10998 11620
rect 11078 11590 11118 11620
rect 11198 11590 11238 11620
rect 11318 11590 11358 11620
rect 11438 11590 11478 11620
rect 11558 11590 11598 11620
rect 11678 11590 11718 11620
rect 11798 11590 11838 11620
rect 11918 11590 11958 11620
rect 12038 11590 12078 11620
rect 12158 11590 12198 11620
rect 12278 11590 12318 11620
rect 12398 11590 12438 11620
rect 12518 11590 12558 11620
rect 12638 11590 12678 11620
rect 12758 11590 12798 11620
rect 12878 11590 12918 11620
rect 13638 11590 13678 11620
rect 13758 11590 13798 11620
rect 13878 11590 13918 11620
rect 13998 11590 14038 11620
rect 14118 11590 14158 11620
rect 14238 11590 14278 11620
rect 14358 11590 14398 11620
rect 14478 11590 14518 11620
rect 14598 11590 14638 11620
rect 14718 11590 14758 11620
rect 14838 11590 14878 11620
rect 14958 11590 14998 11620
rect 15078 11590 15118 11620
rect 15198 11590 15238 11620
rect 15318 11590 15358 11620
rect 15438 11590 15478 11620
rect 15558 11590 15598 11620
rect 15678 11590 15718 11620
rect 15798 11590 15838 11620
rect 15918 11590 15958 11620
rect 10528 11570 10638 11590
rect 10528 11530 10538 11570
rect 10578 11560 10638 11570
rect 12878 11570 12988 11590
rect 12878 11560 12938 11570
rect 10578 11530 10588 11560
rect 10528 11510 10588 11530
rect 12928 11530 12938 11560
rect 12978 11530 12988 11570
rect 12928 11510 12988 11530
rect 13568 11570 13678 11590
rect 13568 11530 13578 11570
rect 13618 11560 13678 11570
rect 15918 11570 16028 11590
rect 15918 11560 15978 11570
rect 13618 11530 13628 11560
rect 13568 11510 13628 11530
rect 15968 11530 15978 11560
rect 16018 11530 16028 11570
rect 15968 11510 16028 11530
rect 19538 11510 19568 11540
rect 19668 11520 19698 11540
rect 19798 11520 19828 11540
rect 19668 11510 19828 11520
rect 19618 11490 19828 11510
rect 19928 11520 19958 11540
rect 20058 11520 20088 11540
rect 19928 11510 20088 11520
rect 20188 11510 20218 11540
rect 20678 11510 20708 11540
rect 20808 11520 20838 11540
rect 20938 11520 20968 11540
rect 21068 11520 21098 11540
rect 21198 11520 21228 11540
rect 19928 11490 20138 11510
rect 20808 11490 21228 11520
rect 21328 11510 21358 11540
rect 21818 11510 21848 11540
rect 21948 11510 21978 11540
rect 21898 11490 21978 11510
rect 19618 11450 19638 11490
rect 19678 11450 19698 11490
rect 19618 11430 19698 11450
rect 20058 11450 20078 11490
rect 20118 11450 20138 11490
rect 20058 11430 20138 11450
rect 20848 11480 20928 11490
rect 20848 11440 20868 11480
rect 20908 11440 20928 11480
rect 20848 11420 20928 11440
rect 21898 11450 21918 11490
rect 21958 11460 21978 11490
rect 22078 11460 22108 11540
rect 22208 11460 22238 11540
rect 22338 11460 22368 11540
rect 22468 11510 22498 11540
rect 22738 11490 22818 11510
rect 22738 11460 22758 11490
rect 21958 11450 22758 11460
rect 22798 11450 22818 11490
rect 21898 11430 22818 11450
rect 21898 11270 21978 11290
rect 21898 11230 21918 11270
rect 21958 11230 21978 11270
rect 21898 11210 21978 11230
rect 21948 11170 21978 11210
rect 19708 11150 19788 11170
rect 19708 11110 19728 11150
rect 19768 11110 19788 11150
rect 20758 11150 20838 11170
rect 20758 11110 20778 11150
rect 20818 11110 20838 11150
rect 21198 11150 21278 11170
rect 21198 11110 21218 11150
rect 21258 11110 21278 11150
rect 19538 11060 19568 11090
rect 19668 11080 20088 11110
rect 20758 11090 20968 11110
rect 19668 11060 19698 11080
rect 19798 11060 19828 11080
rect 19928 11060 19958 11080
rect 20058 11060 20088 11080
rect 20188 11060 20218 11090
rect 20678 11060 20708 11090
rect 20808 11080 20968 11090
rect 20808 11060 20838 11080
rect 20938 11060 20968 11080
rect 21068 11090 21278 11110
rect 21948 11150 22818 11170
rect 21948 11140 22758 11150
rect 21068 11080 21228 11090
rect 21068 11060 21098 11080
rect 21198 11060 21228 11080
rect 21328 11060 21358 11090
rect 21818 11060 21848 11090
rect 21948 11060 21978 11140
rect 22078 11060 22108 11140
rect 22208 11060 22238 11140
rect 22338 11060 22368 11140
rect 22738 11110 22758 11140
rect 22798 11110 22818 11150
rect 22738 11090 22818 11110
rect 22468 11060 22498 11090
rect 19538 10930 19568 10960
rect 19668 10930 19698 10960
rect 19798 10930 19828 10960
rect 19928 10930 19958 10960
rect 20058 10930 20088 10960
rect 20188 10930 20218 10960
rect 20678 10930 20708 10960
rect 20808 10930 20838 10960
rect 20938 10930 20968 10960
rect 21068 10930 21098 10960
rect 21198 10930 21228 10960
rect 21328 10930 21358 10960
rect 21818 10930 21848 10960
rect 21948 10930 21978 10960
rect 22078 10930 22108 10960
rect 22208 10930 22238 10960
rect 22338 10930 22368 10960
rect 22468 10930 22498 10960
rect 19508 10910 19598 10930
rect 19508 10860 19528 10910
rect 19578 10860 19598 10910
rect 19508 10840 19598 10860
rect 20158 10910 20248 10930
rect 20158 10860 20178 10910
rect 20228 10860 20248 10910
rect 20158 10840 20248 10860
rect 20648 10910 20728 10930
rect 20648 10870 20668 10910
rect 20708 10870 20728 10910
rect 20648 10850 20728 10870
rect 21308 10910 21388 10930
rect 21308 10870 21328 10910
rect 21368 10870 21388 10910
rect 21308 10850 21388 10870
rect 21788 10910 21868 10930
rect 21788 10870 21808 10910
rect 21848 10870 21868 10910
rect 21788 10850 21868 10870
rect 22448 10910 22528 10930
rect 22448 10870 22468 10910
rect 22508 10870 22528 10910
rect 22448 10850 22528 10870
rect 11898 10750 11968 10770
rect 11898 10710 11908 10750
rect 11948 10710 11968 10750
rect 11898 10690 11968 10710
rect 12068 10750 12148 10770
rect 12068 10710 12088 10750
rect 12128 10710 12148 10750
rect 12068 10690 12148 10710
rect 12248 10750 12328 10770
rect 12248 10710 12268 10750
rect 12308 10710 12328 10750
rect 12248 10690 12328 10710
rect 12428 10750 12508 10770
rect 12428 10710 12448 10750
rect 12488 10710 12508 10750
rect 12428 10690 12508 10710
rect 12608 10750 12688 10770
rect 12608 10710 12628 10750
rect 12668 10710 12688 10750
rect 12608 10690 12688 10710
rect 12788 10750 12868 10770
rect 12788 10710 12808 10750
rect 12848 10710 12868 10750
rect 12788 10690 12868 10710
rect 12968 10750 13048 10770
rect 12968 10710 12988 10750
rect 13028 10710 13048 10750
rect 12968 10690 13048 10710
rect 13148 10750 13218 10770
rect 13148 10710 13168 10750
rect 13208 10710 13218 10750
rect 13148 10690 13218 10710
rect 13338 10750 13408 10770
rect 13338 10710 13348 10750
rect 13388 10710 13408 10750
rect 13338 10690 13408 10710
rect 13508 10750 13588 10770
rect 13508 10710 13528 10750
rect 13568 10710 13588 10750
rect 13508 10690 13588 10710
rect 13688 10750 13768 10770
rect 13688 10710 13708 10750
rect 13748 10710 13768 10750
rect 13688 10690 13768 10710
rect 13868 10750 13948 10770
rect 13868 10710 13888 10750
rect 13928 10710 13948 10750
rect 13868 10690 13948 10710
rect 14048 10750 14128 10770
rect 14048 10710 14068 10750
rect 14108 10710 14128 10750
rect 14048 10690 14128 10710
rect 14228 10750 14308 10770
rect 14228 10710 14248 10750
rect 14288 10710 14308 10750
rect 14228 10690 14308 10710
rect 14408 10750 14488 10770
rect 14408 10710 14428 10750
rect 14468 10710 14488 10750
rect 14408 10690 14488 10710
rect 14588 10750 14658 10770
rect 14588 10710 14608 10750
rect 14648 10710 14658 10750
rect 14588 10700 14658 10710
rect 11698 10660 11798 10690
rect 11878 10660 11978 10690
rect 12058 10660 12158 10690
rect 12238 10660 12338 10690
rect 12418 10660 12518 10690
rect 12598 10660 12698 10690
rect 12778 10660 12878 10690
rect 12958 10660 13058 10690
rect 13138 10660 13238 10690
rect 13318 10660 13418 10690
rect 13498 10660 13598 10690
rect 13678 10660 13778 10690
rect 13858 10660 13958 10690
rect 14038 10660 14138 10690
rect 14218 10660 14318 10690
rect 14398 10660 14498 10690
rect 14578 10660 14678 10700
rect 14758 10660 14858 10690
rect 19398 10610 19478 10630
rect 19398 10570 19418 10610
rect 19458 10580 19478 10610
rect 21398 10610 21478 10630
rect 21398 10580 21418 10610
rect 19458 10570 19588 10580
rect 15708 10550 15788 10570
rect 19398 10550 19588 10570
rect 21288 10570 21418 10580
rect 21458 10570 21478 10610
rect 21288 10550 21478 10570
rect 15708 10510 15728 10550
rect 15768 10510 15788 10550
rect 19488 10520 19588 10550
rect 19688 10520 19788 10550
rect 19888 10520 19988 10550
rect 20088 10520 20188 10550
rect 20288 10520 20388 10550
rect 20488 10520 20588 10550
rect 20688 10520 20788 10550
rect 20888 10520 20988 10550
rect 21088 10520 21188 10550
rect 21288 10520 21388 10550
rect 15568 10460 15598 10490
rect 15678 10480 15818 10510
rect 15678 10460 15708 10480
rect 15788 10460 15818 10480
rect 15898 10460 15928 10490
rect 15568 10240 15598 10260
rect 15498 10210 15598 10240
rect 15678 10230 15708 10260
rect 15788 10230 15818 10260
rect 15898 10240 15928 10260
rect 19488 10240 19588 10270
rect 19688 10250 19788 10270
rect 19888 10250 19988 10270
rect 20088 10250 20188 10270
rect 20288 10250 20388 10270
rect 20488 10250 20588 10270
rect 20688 10250 20788 10270
rect 20888 10250 20988 10270
rect 21088 10250 21188 10270
rect 15898 10210 15998 10240
rect 19688 10220 21188 10250
rect 21288 10240 21388 10270
rect 15498 10170 15508 10210
rect 15548 10170 15558 10210
rect 15498 10150 15558 10170
rect 15938 10170 15948 10210
rect 15988 10170 15998 10210
rect 15938 10150 15998 10170
rect 20198 10180 20218 10220
rect 20258 10180 20278 10220
rect 20198 10160 20278 10180
rect 20598 10180 20618 10220
rect 20658 10180 20678 10220
rect 20598 10160 20678 10180
rect 11698 10030 11798 10060
rect 11878 10030 11978 10060
rect 12058 10030 12158 10060
rect 12238 10030 12338 10060
rect 12418 10030 12518 10060
rect 12598 10030 12698 10060
rect 12778 10030 12878 10060
rect 12958 10030 13058 10060
rect 13138 10030 13238 10060
rect 13318 10030 13418 10060
rect 13498 10030 13598 10060
rect 13678 10030 13778 10060
rect 13858 10030 13958 10060
rect 14038 10030 14138 10060
rect 14218 10030 14318 10060
rect 14398 10030 14498 10060
rect 14578 10030 14678 10060
rect 14758 10030 14858 10060
rect 11618 10010 11798 10030
rect 11618 9970 11638 10010
rect 11678 10000 11798 10010
rect 14758 10010 14938 10030
rect 14758 10000 14878 10010
rect 11678 9970 11698 10000
rect 11618 9950 11698 9970
rect 14858 9970 14878 10000
rect 14918 9970 14938 10010
rect 19242 10024 19672 10040
rect 19242 9990 19258 10024
rect 19292 9990 19672 10024
rect 19242 9974 19672 9990
rect 20152 10024 20582 10040
rect 20152 9990 20532 10024
rect 20566 9990 20582 10024
rect 20152 9974 20582 9990
rect 14858 9950 14938 9970
rect 11804 9742 11862 9760
rect 11804 9708 11816 9742
rect 11850 9708 11862 9742
rect 11804 9690 11862 9708
rect 11914 9742 11972 9760
rect 11914 9708 11926 9742
rect 11960 9708 11972 9742
rect 11914 9690 11972 9708
rect 12024 9742 12082 9760
rect 12024 9708 12036 9742
rect 12070 9708 12082 9742
rect 12024 9690 12082 9708
rect 12134 9742 12192 9760
rect 12134 9708 12146 9742
rect 12180 9708 12192 9742
rect 12134 9690 12192 9708
rect 12244 9742 12302 9760
rect 12244 9708 12256 9742
rect 12290 9708 12302 9742
rect 12244 9690 12302 9708
rect 12354 9742 12412 9760
rect 12354 9708 12366 9742
rect 12400 9708 12412 9742
rect 12354 9690 12412 9708
rect 12464 9742 12522 9760
rect 12464 9708 12476 9742
rect 12510 9708 12522 9742
rect 12464 9690 12522 9708
rect 12574 9742 12632 9760
rect 12574 9708 12586 9742
rect 12620 9708 12632 9742
rect 12574 9690 12632 9708
rect 12684 9742 12742 9760
rect 12684 9708 12696 9742
rect 12730 9708 12742 9742
rect 12684 9690 12742 9708
rect 12794 9742 12852 9760
rect 12794 9708 12806 9742
rect 12840 9708 12852 9742
rect 12794 9690 12852 9708
rect 13704 9742 13762 9760
rect 13704 9708 13716 9742
rect 13750 9708 13762 9742
rect 13704 9690 13762 9708
rect 13814 9742 13872 9760
rect 13814 9708 13826 9742
rect 13860 9708 13872 9742
rect 13814 9690 13872 9708
rect 13924 9742 13982 9760
rect 13924 9708 13936 9742
rect 13970 9708 13982 9742
rect 13924 9690 13982 9708
rect 14034 9742 14092 9760
rect 14034 9708 14046 9742
rect 14080 9708 14092 9742
rect 14034 9690 14092 9708
rect 14144 9742 14202 9760
rect 14144 9708 14156 9742
rect 14190 9708 14202 9742
rect 14144 9690 14202 9708
rect 14254 9742 14312 9760
rect 14254 9708 14266 9742
rect 14300 9708 14312 9742
rect 14254 9690 14312 9708
rect 14364 9742 14422 9760
rect 14364 9708 14376 9742
rect 14410 9708 14422 9742
rect 14364 9690 14422 9708
rect 14474 9742 14532 9760
rect 14474 9708 14486 9742
rect 14520 9708 14532 9742
rect 14474 9690 14532 9708
rect 14584 9742 14642 9760
rect 14584 9708 14596 9742
rect 14630 9708 14642 9742
rect 14584 9690 14642 9708
rect 14694 9742 14752 9760
rect 14694 9708 14706 9742
rect 14740 9708 14752 9742
rect 14694 9690 14752 9708
rect 11708 9660 11738 9690
rect 11818 9660 11848 9690
rect 11928 9660 11958 9690
rect 12038 9660 12068 9690
rect 12148 9660 12178 9690
rect 12258 9660 12288 9690
rect 12368 9660 12398 9690
rect 12478 9660 12508 9690
rect 12588 9660 12618 9690
rect 12698 9660 12728 9690
rect 12808 9660 12838 9690
rect 12918 9660 12948 9690
rect 13608 9660 13638 9690
rect 13718 9660 13748 9690
rect 13828 9660 13858 9690
rect 13938 9660 13968 9690
rect 14048 9660 14078 9690
rect 14158 9660 14188 9690
rect 14268 9660 14298 9690
rect 14378 9660 14408 9690
rect 14488 9660 14518 9690
rect 14598 9660 14628 9690
rect 14708 9660 14738 9690
rect 14818 9660 14848 9690
rect 11708 9430 11738 9460
rect 11818 9430 11848 9460
rect 11928 9430 11958 9460
rect 12038 9430 12068 9460
rect 12148 9430 12178 9460
rect 12258 9430 12288 9460
rect 12368 9430 12398 9460
rect 12478 9430 12508 9460
rect 12588 9430 12618 9460
rect 12698 9430 12728 9460
rect 12808 9430 12838 9460
rect 12918 9430 12948 9460
rect 13608 9430 13638 9460
rect 13718 9430 13748 9460
rect 13828 9430 13858 9460
rect 13938 9430 13968 9460
rect 14048 9430 14078 9460
rect 14158 9430 14188 9460
rect 14268 9430 14298 9460
rect 14378 9430 14408 9460
rect 14488 9430 14518 9460
rect 14598 9430 14628 9460
rect 14708 9430 14738 9460
rect 14818 9430 14848 9460
rect 11628 9410 11738 9430
rect 11628 9370 11648 9410
rect 11688 9400 11738 9410
rect 12918 9410 13028 9430
rect 12918 9400 12968 9410
rect 11688 9370 11708 9400
rect 11628 9350 11708 9370
rect 12948 9370 12968 9400
rect 13008 9370 13028 9410
rect 12948 9350 13028 9370
rect 13528 9410 13638 9430
rect 13528 9370 13548 9410
rect 13588 9400 13638 9410
rect 14818 9410 14928 9430
rect 14818 9400 14868 9410
rect 13588 9370 13608 9400
rect 13528 9350 13608 9370
rect 14848 9370 14868 9400
rect 14908 9370 14928 9410
rect 14848 9350 14928 9370
rect 13848 8170 14258 8200
rect 13328 8090 13358 8120
rect 13438 8090 13468 8120
rect 13848 8090 13878 8170
rect 13958 8090 13988 8120
rect 14228 8090 14258 8170
rect 16868 8180 16978 8200
rect 16868 8140 16918 8180
rect 16958 8140 16978 8180
rect 16868 8120 16978 8140
rect 17528 8180 17608 8200
rect 17528 8140 17548 8180
rect 17588 8140 17608 8180
rect 17528 8120 17608 8140
rect 19338 8130 19418 8150
rect 14338 8090 14368 8120
rect 14748 8090 14778 8120
rect 14858 8090 14888 8120
rect 15258 8090 15288 8120
rect 15588 8090 15618 8120
rect 15918 8090 15948 8120
rect 16478 8090 16508 8120
rect 16868 8090 16898 8120
rect 17258 8090 17288 8120
rect 17548 8090 17578 8120
rect 17938 8090 17968 8120
rect 19338 8090 19358 8130
rect 19398 8100 19418 8130
rect 19868 8120 20848 8150
rect 19868 8100 19988 8120
rect 19398 8090 19548 8100
rect 19338 8070 19548 8090
rect 19428 8040 19548 8070
rect 19648 8060 19988 8100
rect 20728 8100 20848 8120
rect 22378 8130 22458 8150
rect 22378 8100 22398 8130
rect 19648 8040 19768 8060
rect 19868 8040 19988 8060
rect 20088 8040 20208 8070
rect 20508 8040 20628 8070
rect 20728 8060 21068 8100
rect 20728 8040 20848 8060
rect 20948 8040 21068 8060
rect 21168 8040 21288 8070
rect 21588 8040 21708 8070
rect 21808 8060 22148 8100
rect 21808 8040 21928 8060
rect 22028 8040 22148 8060
rect 22248 8090 22398 8100
rect 22438 8090 22458 8130
rect 22248 8070 22458 8090
rect 22248 8040 22368 8070
rect 13328 7820 13358 7890
rect 13128 7800 13358 7820
rect 13128 7760 13148 7800
rect 13188 7790 13358 7800
rect 13188 7760 13208 7790
rect 13128 7740 13208 7760
rect 13328 7670 13358 7790
rect 13438 7860 13468 7890
rect 13438 7840 13538 7860
rect 13848 7850 13878 7890
rect 13438 7800 13478 7840
rect 13518 7800 13538 7840
rect 13438 7780 13538 7800
rect 13628 7820 13878 7850
rect 13438 7670 13468 7780
rect 13628 7360 13658 7820
rect 13848 7670 13878 7820
rect 13958 7780 13988 7890
rect 13958 7760 14058 7780
rect 13958 7720 13998 7760
rect 14038 7720 14058 7760
rect 13958 7700 14058 7720
rect 13958 7670 13988 7700
rect 14228 7670 14258 7890
rect 14338 7860 14368 7890
rect 14338 7840 14438 7860
rect 14748 7850 14778 7890
rect 14338 7800 14378 7840
rect 14418 7800 14438 7840
rect 14338 7780 14438 7800
rect 14528 7820 14778 7850
rect 14338 7670 14368 7780
rect 13578 7340 13658 7360
rect 13578 7300 13598 7340
rect 13638 7300 13658 7340
rect 13578 7280 13658 7300
rect 14528 7360 14558 7820
rect 14748 7670 14778 7820
rect 14858 7760 14888 7890
rect 15048 7790 15208 7810
rect 15048 7760 15068 7790
rect 14858 7750 15068 7760
rect 15108 7750 15148 7790
rect 15188 7750 15208 7790
rect 14858 7730 15208 7750
rect 15258 7790 15288 7890
rect 15458 7790 15538 7810
rect 15258 7760 15478 7790
rect 14858 7670 14888 7730
rect 15258 7670 15288 7760
rect 15458 7750 15478 7760
rect 15518 7750 15538 7790
rect 15458 7730 15538 7750
rect 15588 7790 15618 7890
rect 15788 7790 15868 7810
rect 15588 7760 15808 7790
rect 15588 7670 15618 7760
rect 15788 7750 15808 7760
rect 15848 7750 15868 7790
rect 15788 7730 15868 7750
rect 15918 7790 15948 7890
rect 16478 7820 16508 7890
rect 16868 7860 16898 7890
rect 16078 7790 16158 7810
rect 15918 7760 16098 7790
rect 15918 7670 15948 7760
rect 16078 7750 16098 7760
rect 16138 7750 16158 7790
rect 16078 7730 16158 7750
rect 16228 7800 16508 7820
rect 16228 7760 16248 7800
rect 16288 7790 16508 7800
rect 16288 7760 16308 7790
rect 16228 7740 16308 7760
rect 16478 7670 16508 7790
rect 16948 7770 17028 7790
rect 16948 7730 16968 7770
rect 17008 7740 17028 7770
rect 17258 7740 17288 7890
rect 17548 7870 17578 7890
rect 17338 7850 17578 7870
rect 17338 7810 17358 7850
rect 17398 7840 17578 7850
rect 17398 7810 17418 7840
rect 17338 7800 17418 7810
rect 17938 7740 17968 7890
rect 17008 7730 17968 7740
rect 16948 7710 17968 7730
rect 16868 7670 16898 7700
rect 17258 7670 17288 7710
rect 17548 7670 17578 7710
rect 14478 7340 14558 7360
rect 14478 7300 14498 7340
rect 14538 7300 14558 7340
rect 14478 7280 14558 7300
rect 19428 7610 19548 7640
rect 19648 7620 19768 7640
rect 19868 7620 19988 7640
rect 19648 7600 19988 7620
rect 19648 7590 19798 7600
rect 19778 7560 19798 7590
rect 19838 7590 19988 7600
rect 20088 7620 20208 7640
rect 20508 7620 20628 7640
rect 20088 7590 20628 7620
rect 20728 7620 20848 7640
rect 20948 7620 21068 7640
rect 20728 7590 21068 7620
rect 21168 7620 21288 7640
rect 21588 7620 21708 7640
rect 21168 7590 21708 7620
rect 21808 7610 21928 7640
rect 22028 7610 22148 7640
rect 22248 7610 22368 7640
rect 19838 7560 19858 7590
rect 19778 7540 19858 7560
rect 20318 7550 20338 7590
rect 20378 7550 20398 7590
rect 20318 7530 20398 7550
rect 21398 7550 21418 7590
rect 21458 7550 21478 7590
rect 21398 7530 21478 7550
rect 21808 7580 22148 7610
rect 21808 7560 21888 7580
rect 21808 7520 21828 7560
rect 21868 7520 21888 7560
rect 21808 7500 21888 7520
rect 22068 7560 22148 7580
rect 22068 7520 22088 7560
rect 22128 7520 22148 7560
rect 22068 7500 22148 7520
rect 13328 7240 13358 7270
rect 13438 7240 13468 7270
rect 13848 7240 13878 7270
rect 13958 7240 13988 7270
rect 14228 7240 14258 7270
rect 14338 7240 14368 7270
rect 14748 7240 14778 7270
rect 14858 7240 14888 7270
rect 15258 7240 15288 7270
rect 15588 7240 15618 7270
rect 15918 7240 15948 7270
rect 16478 7240 16508 7270
rect 16868 7240 16898 7270
rect 17258 7240 17288 7270
rect 17548 7240 17578 7270
rect 13698 7220 13778 7240
rect 13698 7180 13718 7220
rect 13758 7180 13778 7220
rect 13698 7160 13778 7180
rect 16818 7220 16898 7240
rect 16818 7180 16838 7220
rect 16878 7180 16898 7220
rect 16818 7170 16898 7180
rect 21368 7060 21448 7080
rect 20198 7030 20278 7050
rect 15248 7000 15328 7010
rect 20198 7000 20218 7030
rect 15248 6960 15268 7000
rect 15308 6960 15328 7000
rect 19848 6990 20218 7000
rect 20258 7000 20278 7030
rect 20958 7030 21038 7050
rect 20258 6990 20628 7000
rect 20958 6990 20978 7030
rect 21018 6990 21038 7030
rect 21368 7020 21388 7060
rect 21428 7020 21448 7060
rect 21368 7000 21448 7020
rect 22068 7060 22148 7080
rect 22068 7020 22088 7060
rect 22128 7020 22148 7060
rect 22068 7000 22148 7020
rect 15248 6940 15328 6960
rect 19628 6940 19748 6970
rect 19848 6960 20628 6990
rect 19848 6940 19968 6960
rect 20068 6940 20188 6960
rect 20288 6940 20408 6960
rect 20508 6940 20628 6960
rect 20728 6960 21268 6990
rect 20728 6940 20848 6960
rect 21148 6940 21268 6960
rect 21368 6970 22148 7000
rect 21368 6940 21488 6970
rect 21588 6940 21708 6970
rect 21808 6940 21928 6970
rect 22028 6940 22148 6970
rect 22248 6940 22368 6970
rect 13328 6910 13358 6940
rect 13438 6910 13468 6940
rect 13848 6910 13878 6940
rect 13958 6910 13988 6940
rect 14228 6910 14258 6940
rect 14338 6910 14368 6940
rect 14748 6910 14778 6940
rect 14858 6910 14888 6940
rect 15268 6910 15298 6940
rect 15378 6910 15408 6940
rect 15708 6910 15738 6940
rect 16038 6910 16068 6940
rect 16478 6910 16508 6940
rect 16868 6910 16898 6940
rect 17258 6910 17288 6940
rect 17548 6910 17578 6940
rect 17938 6910 17968 6940
rect 13578 6880 13658 6900
rect 13578 6840 13598 6880
rect 13638 6840 13658 6880
rect 13578 6820 13658 6840
rect 13128 6420 13208 6440
rect 13128 6380 13148 6420
rect 13188 6390 13208 6420
rect 13328 6390 13358 6510
rect 13188 6380 13358 6390
rect 13128 6360 13358 6380
rect 13328 6290 13358 6360
rect 13438 6400 13468 6510
rect 13438 6380 13538 6400
rect 13438 6340 13478 6380
rect 13518 6340 13538 6380
rect 13438 6320 13538 6340
rect 13628 6360 13658 6820
rect 14478 6880 14558 6900
rect 14478 6840 14498 6880
rect 14538 6840 14558 6880
rect 14478 6820 14558 6840
rect 13848 6360 13878 6510
rect 13628 6330 13878 6360
rect 13438 6290 13468 6320
rect 13848 6290 13878 6330
rect 13958 6480 13988 6510
rect 13958 6460 14058 6480
rect 13958 6420 13998 6460
rect 14038 6420 14058 6460
rect 13958 6400 14058 6420
rect 13958 6290 13988 6400
rect 14228 6290 14258 6510
rect 14338 6400 14368 6510
rect 14338 6380 14438 6400
rect 14338 6340 14378 6380
rect 14418 6340 14438 6380
rect 14338 6320 14438 6340
rect 14528 6360 14558 6820
rect 19628 6510 19748 6540
rect 14748 6360 14778 6510
rect 14528 6330 14778 6360
rect 14338 6290 14368 6320
rect 14748 6290 14778 6330
rect 14858 6360 14888 6510
rect 15028 6390 15108 6410
rect 15028 6360 15048 6390
rect 14858 6350 15048 6360
rect 15088 6350 15108 6390
rect 14858 6330 15108 6350
rect 14858 6290 14888 6330
rect 15268 6290 15298 6510
rect 15378 6290 15408 6510
rect 15458 6430 15538 6450
rect 15458 6390 15478 6430
rect 15518 6420 15538 6430
rect 15708 6420 15738 6510
rect 15518 6390 15738 6420
rect 15458 6370 15538 6390
rect 15708 6290 15738 6390
rect 15788 6430 15868 6450
rect 15788 6390 15808 6430
rect 15848 6420 15868 6430
rect 16038 6420 16068 6510
rect 15848 6390 16068 6420
rect 15788 6370 15868 6390
rect 16038 6290 16068 6390
rect 16118 6430 16198 6450
rect 16118 6390 16138 6430
rect 16178 6390 16198 6430
rect 16478 6420 16508 6510
rect 16868 6450 16898 6510
rect 16118 6370 16198 6390
rect 16248 6400 16508 6420
rect 16248 6360 16268 6400
rect 16308 6390 16508 6400
rect 16308 6360 16328 6390
rect 16248 6340 16328 6360
rect 16478 6290 16508 6390
rect 16818 6430 16898 6450
rect 16818 6390 16838 6430
rect 16878 6390 16898 6430
rect 17258 6400 17288 6510
rect 17548 6480 17578 6510
rect 17338 6460 17768 6480
rect 17338 6420 17358 6460
rect 17398 6450 17708 6460
rect 17398 6420 17418 6450
rect 17338 6400 17418 6420
rect 17688 6420 17708 6450
rect 17748 6420 17768 6460
rect 17688 6400 17768 6420
rect 16818 6370 16898 6390
rect 16868 6290 16898 6370
rect 17208 6380 17288 6400
rect 17208 6340 17228 6380
rect 17268 6350 17288 6380
rect 17938 6350 17968 6510
rect 19538 6490 19748 6510
rect 19538 6450 19558 6490
rect 19598 6480 19748 6490
rect 19848 6520 19968 6540
rect 20068 6520 20188 6540
rect 20288 6520 20408 6540
rect 20508 6520 20628 6540
rect 19848 6480 20628 6520
rect 20728 6510 20848 6540
rect 21148 6510 21268 6540
rect 21368 6520 21488 6540
rect 21588 6520 21708 6540
rect 21808 6520 21928 6540
rect 22028 6520 22148 6540
rect 21368 6480 22148 6520
rect 22248 6510 22368 6540
rect 22248 6490 22458 6510
rect 22248 6480 22398 6490
rect 19598 6450 19618 6480
rect 19538 6430 19618 6450
rect 22378 6450 22398 6480
rect 22438 6450 22458 6490
rect 22378 6430 22458 6450
rect 17268 6340 17968 6350
rect 17208 6320 17968 6340
rect 17258 6290 17288 6320
rect 17548 6290 17578 6320
rect 13328 6060 13358 6090
rect 13438 6060 13468 6090
rect 13848 6010 13878 6090
rect 13958 6060 13988 6090
rect 14228 6010 14258 6090
rect 14338 6060 14368 6090
rect 14748 6060 14778 6090
rect 14858 6060 14888 6090
rect 15268 6060 15298 6090
rect 15378 6060 15408 6090
rect 15708 6060 15738 6090
rect 16038 6060 16068 6090
rect 16478 6060 16508 6090
rect 16868 6060 16898 6090
rect 17258 6060 17288 6090
rect 17548 6060 17578 6090
rect 13848 5980 14258 6010
rect 15378 6040 15458 6060
rect 15378 6000 15398 6040
rect 15438 6000 15458 6040
rect 15378 5980 15458 6000
rect 23278 5430 23578 5460
rect 23798 5430 24098 5460
rect 24318 5430 24618 5460
rect 24838 5430 25138 5460
rect 23278 5000 23578 5030
rect 23798 5000 24098 5030
rect 24318 5000 24618 5030
rect 24838 5000 25138 5030
rect 23388 4980 23468 5000
rect 23388 4940 23408 4980
rect 23448 4940 23468 4980
rect 23388 4920 23468 4940
rect 23908 4980 23988 5000
rect 23908 4940 23928 4980
rect 23968 4940 23988 4980
rect 23908 4920 23988 4940
rect 24428 4980 24508 5000
rect 24428 4940 24448 4980
rect 24488 4940 24508 4980
rect 24428 4920 24508 4940
rect 24958 4980 25018 5000
rect 24958 4940 24968 4980
rect 25008 4940 25018 4980
rect 24958 4920 25018 4940
rect 23278 4740 23308 4770
rect 23798 4740 23828 4770
rect 24318 4740 24348 4770
rect 13018 3620 13118 3640
rect 14138 3620 14228 3640
rect 13018 3580 13038 3620
rect 13078 3580 13118 3620
rect 13018 3560 13118 3580
rect 13328 3600 13408 3620
rect 13328 3560 13348 3600
rect 13388 3560 13408 3600
rect 14138 3580 14158 3620
rect 14198 3580 14228 3620
rect 14138 3560 14228 3580
rect 14278 3620 14338 3640
rect 14278 3580 14288 3620
rect 14328 3580 14338 3620
rect 14278 3560 14338 3580
rect 15398 3620 15488 3640
rect 15398 3580 15418 3620
rect 15458 3580 15488 3620
rect 15398 3560 15488 3580
rect 17158 3630 17238 3640
rect 17158 3590 17178 3630
rect 17218 3600 17238 3630
rect 19658 3620 19768 3640
rect 17218 3590 17318 3600
rect 17158 3570 17318 3590
rect 19658 3580 19708 3620
rect 19748 3580 19768 3620
rect 20958 3620 21068 3640
rect 20958 3580 21008 3620
rect 21048 3580 21068 3620
rect 22258 3620 22368 3640
rect 22258 3580 22308 3620
rect 22348 3580 22368 3620
rect 12668 3530 12698 3560
rect 13088 3530 13118 3560
rect 13198 3530 13228 3560
rect 13328 3540 13408 3560
rect 12358 3500 12438 3520
rect 12358 3460 12378 3500
rect 12418 3460 12438 3500
rect 12358 3440 12438 3460
rect 12488 3300 12568 3320
rect 12488 3260 12508 3300
rect 12548 3260 12568 3300
rect 12668 3260 12698 3430
rect 13088 3400 13118 3430
rect 13198 3370 13228 3430
rect 13328 3370 13358 3540
rect 13758 3530 13788 3560
rect 13868 3530 13898 3560
rect 14198 3530 14228 3560
rect 14308 3530 14338 3560
rect 14418 3530 14448 3560
rect 15038 3530 15068 3560
rect 15458 3530 15488 3560
rect 15568 3530 15598 3560
rect 15908 3530 15938 3560
rect 16018 3530 16048 3560
rect 16268 3530 16298 3560
rect 16378 3530 16408 3560
rect 16848 3530 16878 3560
rect 16958 3530 16988 3560
rect 17288 3530 17318 3570
rect 17398 3530 17428 3560
rect 17908 3530 17938 3560
rect 18248 3530 18278 3560
rect 18358 3530 18388 3560
rect 18608 3550 18748 3580
rect 19658 3560 19768 3580
rect 18608 3530 18638 3550
rect 18718 3530 18748 3550
rect 19208 3530 19238 3560
rect 19548 3530 19578 3560
rect 19658 3530 19688 3560
rect 19908 3550 20048 3580
rect 20958 3560 21068 3580
rect 19908 3530 19938 3550
rect 20018 3530 20048 3550
rect 20508 3530 20538 3560
rect 20848 3530 20878 3560
rect 20958 3530 20988 3560
rect 21208 3550 21348 3580
rect 22258 3560 22368 3580
rect 21208 3530 21238 3550
rect 21318 3530 21348 3550
rect 21808 3530 21838 3560
rect 22148 3530 22178 3560
rect 22258 3530 22288 3560
rect 22508 3550 22648 3580
rect 22508 3530 22538 3550
rect 22618 3530 22648 3550
rect 13198 3340 13358 3370
rect 13608 3380 13688 3400
rect 13608 3350 13628 3380
rect 13068 3300 13148 3320
rect 13068 3260 13088 3300
rect 13128 3260 13148 3300
rect 12488 3240 12568 3260
rect 12618 3240 13148 3260
rect 12508 3210 12538 3240
rect 12618 3230 13118 3240
rect 12618 3210 12648 3230
rect 12728 3210 12758 3230
rect 12838 3210 12868 3230
rect 13088 3210 13118 3230
rect 13198 3210 13228 3340
rect 12508 3080 12538 3110
rect 12618 3080 12648 3110
rect 12728 3080 12758 3110
rect 12838 3080 12868 3110
rect 13088 3080 13118 3110
rect 13198 3080 13228 3110
rect 13328 3100 13358 3340
rect 13538 3340 13628 3350
rect 13668 3340 13688 3380
rect 13538 3320 13688 3340
rect 13408 3300 13488 3320
rect 13408 3260 13428 3300
rect 13468 3260 13488 3300
rect 13408 3240 13488 3260
rect 13538 3210 13568 3320
rect 13758 3270 13788 3430
rect 13868 3400 13898 3430
rect 14008 3420 14088 3440
rect 14008 3400 14028 3420
rect 13868 3380 14028 3400
rect 14068 3380 14088 3420
rect 13868 3370 14088 3380
rect 14008 3360 14088 3370
rect 13988 3300 14068 3310
rect 13988 3270 14008 3300
rect 13648 3260 14008 3270
rect 14048 3260 14068 3300
rect 13648 3240 14068 3260
rect 13648 3210 13678 3240
rect 13758 3210 13788 3240
rect 13868 3210 13898 3240
rect 14198 3210 14228 3430
rect 14308 3210 14338 3430
rect 14418 3210 14448 3430
rect 15038 3390 15068 3430
rect 15458 3400 15488 3430
rect 14708 3360 15068 3390
rect 14508 3300 14588 3310
rect 14508 3260 14528 3300
rect 14568 3270 14588 3300
rect 14708 3270 14738 3360
rect 14568 3260 14738 3270
rect 14508 3240 14738 3260
rect 14858 3300 14938 3310
rect 14858 3260 14878 3300
rect 14918 3260 14938 3300
rect 15038 3260 15068 3360
rect 15568 3390 15598 3430
rect 15708 3420 15788 3440
rect 15708 3390 15728 3420
rect 15568 3380 15728 3390
rect 15768 3380 15788 3420
rect 15908 3410 15938 3430
rect 16018 3410 16048 3430
rect 15908 3380 16048 3410
rect 16268 3410 16298 3430
rect 16378 3410 16408 3430
rect 16268 3380 16408 3410
rect 15568 3360 15788 3380
rect 15438 3300 15518 3320
rect 15438 3260 15458 3300
rect 15498 3260 15518 3300
rect 14858 3240 14938 3260
rect 14988 3240 15518 3260
rect 14528 3210 14558 3240
rect 14878 3210 14908 3240
rect 14988 3230 15488 3240
rect 14988 3210 15018 3230
rect 15098 3210 15128 3230
rect 15208 3210 15238 3230
rect 15458 3210 15488 3230
rect 15568 3210 15598 3360
rect 15648 3300 15728 3310
rect 15888 3300 15968 3320
rect 15648 3260 15668 3300
rect 15708 3270 15908 3300
rect 15708 3260 15728 3270
rect 15648 3240 15728 3260
rect 15888 3260 15908 3270
rect 15948 3260 15968 3300
rect 15888 3240 15968 3260
rect 16018 3210 16048 3380
rect 16378 3340 16408 3380
rect 16698 3380 16778 3400
rect 16498 3350 16578 3370
rect 16698 3350 16718 3380
rect 16498 3340 16518 3350
rect 16228 3310 16308 3330
rect 16228 3270 16248 3310
rect 16288 3270 16308 3310
rect 16228 3250 16308 3270
rect 16378 3310 16518 3340
rect 16558 3310 16578 3350
rect 16378 3210 16408 3310
rect 16498 3290 16578 3310
rect 16628 3340 16718 3350
rect 16758 3340 16778 3380
rect 16628 3320 16778 3340
rect 16628 3210 16658 3320
rect 16848 3270 16878 3430
rect 16958 3400 16988 3430
rect 17098 3420 17178 3440
rect 17688 3500 17768 3520
rect 17688 3470 17708 3500
rect 17528 3460 17708 3470
rect 17748 3460 17768 3500
rect 17528 3440 17768 3460
rect 17098 3400 17118 3420
rect 16958 3380 17118 3400
rect 17158 3380 17178 3420
rect 16958 3370 17178 3380
rect 17098 3360 17178 3370
rect 17128 3300 17208 3310
rect 17128 3270 17148 3300
rect 16738 3260 17148 3270
rect 17188 3260 17208 3300
rect 16738 3240 17208 3260
rect 16738 3210 16768 3240
rect 16848 3210 16878 3240
rect 16958 3210 16988 3240
rect 17288 3210 17318 3430
rect 17398 3390 17428 3430
rect 17528 3390 17558 3440
rect 17908 3390 17938 3430
rect 18248 3400 18278 3430
rect 18358 3410 18388 3430
rect 17398 3360 17558 3390
rect 17668 3360 17978 3390
rect 17398 3210 17428 3360
rect 17488 3300 17568 3310
rect 17488 3260 17508 3300
rect 17548 3270 17568 3300
rect 17668 3270 17698 3360
rect 17548 3260 17698 3270
rect 17488 3240 17698 3260
rect 17818 3300 17898 3310
rect 17818 3260 17838 3300
rect 17878 3260 17898 3300
rect 17818 3240 17898 3260
rect 17948 3260 17978 3360
rect 18228 3380 18308 3400
rect 18358 3380 18558 3410
rect 18608 3400 18638 3430
rect 18228 3340 18248 3380
rect 18288 3340 18308 3380
rect 18228 3320 18308 3340
rect 18528 3350 18558 3380
rect 18528 3320 18638 3350
rect 18398 3300 18478 3320
rect 18398 3260 18418 3300
rect 18458 3260 18478 3300
rect 17508 3210 17538 3240
rect 17838 3210 17868 3240
rect 17948 3230 18528 3260
rect 17948 3210 17978 3230
rect 18058 3210 18088 3230
rect 18168 3210 18198 3230
rect 18498 3210 18528 3230
rect 18608 3210 18638 3320
rect 18718 3320 18748 3430
rect 19208 3400 19238 3430
rect 19548 3400 19578 3430
rect 19208 3370 19278 3400
rect 18868 3320 18948 3340
rect 18718 3290 18888 3320
rect 18718 3210 18748 3290
rect 18868 3280 18888 3290
rect 18928 3280 18948 3320
rect 18868 3260 18948 3280
rect 19118 3210 19198 3230
rect 19118 3170 19138 3210
rect 19178 3170 19198 3210
rect 19118 3150 19198 3170
rect 19248 3170 19278 3370
rect 19528 3380 19608 3400
rect 19528 3340 19548 3380
rect 19588 3340 19608 3380
rect 19528 3320 19608 3340
rect 19658 3320 19688 3430
rect 19908 3400 19938 3430
rect 20018 3320 20048 3430
rect 20508 3400 20538 3430
rect 20848 3400 20878 3430
rect 20508 3370 20578 3400
rect 20168 3320 20248 3340
rect 19658 3290 19938 3320
rect 19698 3210 19778 3230
rect 19698 3170 19718 3210
rect 19758 3170 19778 3210
rect 19138 3120 19168 3150
rect 19248 3140 19828 3170
rect 19248 3120 19278 3140
rect 19358 3120 19388 3140
rect 19468 3120 19498 3140
rect 19798 3120 19828 3140
rect 19908 3120 19938 3290
rect 20018 3290 20188 3320
rect 20018 3120 20048 3290
rect 20168 3280 20188 3290
rect 20228 3280 20248 3320
rect 20168 3260 20248 3280
rect 20418 3210 20498 3230
rect 20418 3170 20438 3210
rect 20478 3170 20498 3210
rect 20418 3150 20498 3170
rect 20548 3170 20578 3370
rect 20828 3380 20908 3400
rect 20828 3340 20848 3380
rect 20888 3340 20908 3380
rect 20828 3320 20908 3340
rect 20958 3320 20988 3430
rect 21208 3400 21238 3430
rect 21318 3320 21348 3430
rect 21808 3400 21838 3430
rect 22148 3400 22178 3430
rect 21808 3370 21878 3400
rect 21468 3320 21548 3340
rect 20958 3290 21238 3320
rect 20998 3210 21078 3230
rect 20998 3170 21018 3210
rect 21058 3170 21078 3210
rect 20438 3120 20468 3150
rect 20548 3140 21128 3170
rect 20548 3120 20578 3140
rect 20658 3120 20688 3140
rect 20768 3120 20798 3140
rect 21098 3120 21128 3140
rect 21208 3120 21238 3290
rect 21318 3290 21488 3320
rect 21318 3120 21348 3290
rect 21468 3280 21488 3290
rect 21528 3280 21548 3320
rect 21468 3260 21548 3280
rect 21718 3210 21798 3230
rect 21718 3170 21738 3210
rect 21778 3170 21798 3210
rect 21718 3150 21798 3170
rect 21848 3170 21878 3370
rect 22128 3380 22208 3400
rect 22128 3340 22148 3380
rect 22188 3340 22208 3380
rect 22128 3320 22208 3340
rect 22258 3320 22288 3430
rect 22508 3400 22538 3430
rect 22618 3320 22648 3430
rect 23278 4110 23308 4140
rect 23798 4110 23828 4140
rect 24318 4110 24348 4140
rect 23278 4092 23336 4110
rect 23278 4058 23290 4092
rect 23324 4058 23336 4092
rect 23278 4040 23336 4058
rect 23798 4092 23856 4110
rect 23798 4058 23810 4092
rect 23844 4058 23856 4092
rect 23798 4040 23856 4058
rect 24318 4092 24376 4110
rect 24318 4058 24330 4092
rect 24364 4058 24376 4092
rect 24318 4040 24376 4058
rect 23276 3960 23308 3990
rect 23796 3960 23828 3990
rect 24316 3960 24348 3990
rect 23276 3530 23308 3560
rect 23796 3530 23828 3560
rect 24316 3530 24348 3560
rect 23250 3512 23308 3530
rect 23250 3478 23262 3512
rect 23296 3478 23308 3512
rect 23250 3460 23308 3478
rect 23770 3512 23828 3530
rect 23770 3478 23782 3512
rect 23816 3478 23828 3512
rect 23770 3460 23828 3478
rect 24290 3512 24348 3530
rect 24290 3478 24302 3512
rect 24336 3478 24348 3512
rect 24290 3460 24348 3478
rect 22750 3322 22808 3340
rect 22750 3320 22762 3322
rect 22258 3290 22538 3320
rect 22298 3210 22378 3230
rect 22298 3170 22318 3210
rect 22358 3170 22378 3210
rect 21738 3120 21768 3150
rect 21848 3140 22428 3170
rect 21848 3120 21878 3140
rect 21958 3120 21988 3140
rect 22068 3120 22098 3140
rect 22398 3120 22428 3140
rect 22508 3120 22538 3290
rect 22618 3290 22762 3320
rect 22618 3120 22648 3290
rect 22750 3288 22762 3290
rect 22796 3288 22808 3322
rect 22750 3260 22808 3288
rect 13328 3080 13408 3100
rect 13538 3080 13568 3110
rect 13648 3080 13678 3110
rect 13758 3080 13788 3110
rect 13868 3080 13898 3110
rect 14198 3080 14228 3110
rect 14308 3080 14338 3110
rect 14418 3080 14448 3110
rect 14528 3080 14558 3110
rect 14878 3080 14908 3110
rect 14988 3080 15018 3110
rect 15098 3080 15128 3110
rect 15208 3080 15238 3110
rect 15458 3080 15488 3110
rect 15568 3080 15598 3110
rect 16018 3080 16048 3110
rect 16378 3080 16408 3110
rect 16628 3080 16658 3110
rect 16738 3080 16768 3110
rect 16848 3080 16878 3110
rect 16958 3080 16988 3110
rect 17288 3080 17318 3110
rect 17398 3080 17428 3110
rect 17508 3080 17538 3110
rect 17838 3080 17868 3110
rect 17948 3080 17978 3110
rect 18058 3080 18088 3110
rect 18168 3080 18198 3110
rect 18498 3080 18528 3110
rect 18608 3080 18638 3110
rect 18718 3080 18748 3110
rect 12378 3060 12458 3080
rect 12378 3020 12398 3060
rect 12438 3020 12458 3060
rect 13328 3040 13348 3080
rect 13388 3040 13408 3080
rect 13328 3020 13408 3040
rect 14398 3070 14478 3080
rect 14398 3030 14418 3070
rect 14458 3030 14478 3070
rect 12378 3000 12458 3020
rect 14398 3010 14478 3030
rect 15958 3070 16048 3080
rect 15958 3030 15978 3070
rect 16018 3030 16048 3070
rect 15958 3010 16048 3030
rect 18572 3060 18638 3080
rect 18572 3020 18582 3060
rect 18622 3020 18638 3060
rect 18572 3000 18638 3020
rect 19138 2990 19168 3020
rect 19248 2990 19278 3020
rect 19358 2990 19388 3020
rect 19468 2990 19498 3020
rect 19798 2990 19828 3020
rect 19908 2990 19938 3020
rect 20018 2990 20048 3020
rect 20438 2990 20468 3020
rect 20548 2990 20578 3020
rect 20658 2990 20688 3020
rect 20768 2990 20798 3020
rect 21098 2990 21128 3020
rect 21208 2990 21238 3020
rect 21318 2990 21348 3020
rect 21738 2990 21768 3020
rect 21848 2990 21878 3020
rect 21958 2990 21988 3020
rect 22068 2990 22098 3020
rect 22398 2990 22428 3020
rect 22508 2990 22538 3020
rect 22618 2990 22648 3020
rect 23250 3122 23308 3140
rect 23250 3088 23262 3122
rect 23296 3088 23308 3122
rect 23250 3070 23308 3088
rect 23770 3122 23828 3140
rect 23770 3088 23782 3122
rect 23816 3088 23828 3122
rect 23770 3070 23828 3088
rect 24290 3122 24348 3140
rect 24290 3088 24302 3122
rect 24336 3088 24348 3122
rect 24290 3070 24348 3088
rect 23276 3040 23308 3070
rect 23796 3040 23828 3070
rect 24316 3040 24348 3070
rect 23276 2810 23308 2840
rect 23796 2810 23828 2840
rect 24316 2810 24348 2840
rect 23278 2742 23336 2760
rect 23278 2708 23290 2742
rect 23324 2708 23336 2742
rect 23278 2690 23336 2708
rect 23798 2742 23856 2760
rect 23798 2708 23810 2742
rect 23844 2708 23856 2742
rect 23798 2690 23856 2708
rect 24318 2742 24376 2760
rect 24318 2708 24330 2742
rect 24364 2708 24376 2742
rect 24318 2690 24376 2708
rect 23278 2660 23308 2690
rect 23798 2660 23828 2690
rect 24318 2660 24348 2690
rect 23278 2330 23308 2360
rect 23798 2330 23828 2360
rect 24318 2330 24348 2360
rect 23264 2262 23322 2280
rect 23264 2228 23276 2262
rect 23310 2228 23322 2262
rect 23264 2210 23322 2228
rect 23784 2262 23842 2280
rect 23784 2228 23796 2262
rect 23830 2228 23842 2262
rect 23784 2210 23842 2228
rect 24304 2262 24362 2280
rect 24304 2228 24316 2262
rect 24350 2228 24362 2262
rect 24304 2210 24362 2228
rect 24872 2262 24948 2280
rect 24872 2228 24884 2262
rect 24918 2228 24948 2262
rect 24872 2210 24948 2228
rect 23278 2180 23308 2210
rect 23798 2180 23828 2210
rect 24318 2180 24348 2210
rect 24918 2180 24948 2210
rect 23278 1950 23308 1980
rect 23798 1950 23828 1980
rect 24318 1950 24348 1980
rect 24918 1950 24948 1980
<< polycont >>
rect 11338 13990 11378 14030
rect 11498 13990 11538 14030
rect 11658 13990 11698 14030
rect 11818 13990 11858 14030
rect 11978 13990 12018 14030
rect 12138 13990 12178 14030
rect 12298 13990 12338 14030
rect 12458 13990 12498 14030
rect 12618 13990 12658 14030
rect 12778 13990 12818 14030
rect 12938 13990 12978 14030
rect 13098 13990 13138 14030
rect 13418 13990 13458 14030
rect 13578 13990 13618 14030
rect 13738 13990 13778 14030
rect 13898 13990 13938 14030
rect 14058 13990 14098 14030
rect 14218 13990 14258 14030
rect 14378 13990 14418 14030
rect 14538 13990 14578 14030
rect 14698 13990 14738 14030
rect 14858 13990 14898 14030
rect 15018 13990 15058 14030
rect 15178 13990 15218 14030
rect 10938 13080 10978 13120
rect 11178 13080 11218 13120
rect 11418 13080 11458 13120
rect 11658 13080 11698 13120
rect 12298 13080 12338 13120
rect 12538 13080 12578 13120
rect 12778 13080 12818 13120
rect 13738 13080 13778 13120
rect 13978 13080 14018 13120
rect 14218 13080 14258 13120
rect 14858 13080 14898 13120
rect 15098 13080 15138 13120
rect 15338 13080 15378 13120
rect 15578 13080 15618 13120
rect 11441 12708 11475 12742
rect 11801 12708 11835 12742
rect 11921 12708 11955 12742
rect 12281 12708 12315 12742
rect 12401 12708 12435 12742
rect 11542 12478 11576 12512
rect 11700 12478 11734 12512
rect 12024 12478 12058 12512
rect 12178 12478 12212 12512
rect 12502 12478 12536 12512
rect 14121 12708 14155 12742
rect 14241 12708 14275 12742
rect 14601 12708 14635 12742
rect 14721 12708 14755 12742
rect 15081 12708 15115 12742
rect 20338 12740 20378 12780
rect 20738 12740 20778 12780
rect 14020 12478 14054 12512
rect 14344 12478 14378 12512
rect 14498 12478 14532 12512
rect 14822 12478 14856 12512
rect 14980 12478 15014 12512
rect 19538 12100 19578 12140
rect 21538 12100 21578 12140
rect 10718 11880 10758 11920
rect 10898 11870 10938 11910
rect 11378 11870 11418 11910
rect 11618 11870 11658 11910
rect 12098 11870 12138 11910
rect 12338 11870 12378 11910
rect 12758 11870 12798 11910
rect 13758 11870 13798 11910
rect 14178 11870 14218 11910
rect 14418 11870 14458 11910
rect 14898 11870 14938 11910
rect 15138 11870 15178 11910
rect 15618 11870 15658 11910
rect 15798 11880 15838 11920
rect 19528 11790 19568 11830
rect 20188 11790 20228 11830
rect 20668 11790 20708 11830
rect 21328 11790 21368 11830
rect 21808 11790 21848 11830
rect 22468 11790 22508 11830
rect 10538 11530 10578 11570
rect 12938 11530 12978 11570
rect 13578 11530 13618 11570
rect 15978 11530 16018 11570
rect 19638 11450 19678 11490
rect 20078 11450 20118 11490
rect 20868 11440 20908 11480
rect 21918 11450 21958 11490
rect 22758 11450 22798 11490
rect 21918 11230 21958 11270
rect 19728 11110 19768 11150
rect 20778 11110 20818 11150
rect 21218 11110 21258 11150
rect 22758 11110 22798 11150
rect 19528 10860 19578 10910
rect 20178 10860 20228 10910
rect 20668 10870 20708 10910
rect 21328 10870 21368 10910
rect 21808 10870 21848 10910
rect 22468 10870 22508 10910
rect 11908 10710 11948 10750
rect 12088 10710 12128 10750
rect 12268 10710 12308 10750
rect 12448 10710 12488 10750
rect 12628 10710 12668 10750
rect 12808 10710 12848 10750
rect 12988 10710 13028 10750
rect 13168 10710 13208 10750
rect 13348 10710 13388 10750
rect 13528 10710 13568 10750
rect 13708 10710 13748 10750
rect 13888 10710 13928 10750
rect 14068 10710 14108 10750
rect 14248 10710 14288 10750
rect 14428 10710 14468 10750
rect 14608 10710 14648 10750
rect 19418 10570 19458 10610
rect 21418 10570 21458 10610
rect 15728 10510 15768 10550
rect 15508 10170 15548 10210
rect 15948 10170 15988 10210
rect 20218 10180 20258 10220
rect 20618 10180 20658 10220
rect 11638 9970 11678 10010
rect 14878 9970 14918 10010
rect 19258 9990 19292 10024
rect 20532 9990 20566 10024
rect 11816 9708 11850 9742
rect 11926 9708 11960 9742
rect 12036 9708 12070 9742
rect 12146 9708 12180 9742
rect 12256 9708 12290 9742
rect 12366 9708 12400 9742
rect 12476 9708 12510 9742
rect 12586 9708 12620 9742
rect 12696 9708 12730 9742
rect 12806 9708 12840 9742
rect 13716 9708 13750 9742
rect 13826 9708 13860 9742
rect 13936 9708 13970 9742
rect 14046 9708 14080 9742
rect 14156 9708 14190 9742
rect 14266 9708 14300 9742
rect 14376 9708 14410 9742
rect 14486 9708 14520 9742
rect 14596 9708 14630 9742
rect 14706 9708 14740 9742
rect 11648 9370 11688 9410
rect 12968 9370 13008 9410
rect 13548 9370 13588 9410
rect 14868 9370 14908 9410
rect 16918 8140 16958 8180
rect 17548 8140 17588 8180
rect 19358 8090 19398 8130
rect 22398 8090 22438 8130
rect 13148 7760 13188 7800
rect 13478 7800 13518 7840
rect 13998 7720 14038 7760
rect 14378 7800 14418 7840
rect 13598 7300 13638 7340
rect 15068 7750 15108 7790
rect 15148 7750 15188 7790
rect 15478 7750 15518 7790
rect 15808 7750 15848 7790
rect 16098 7750 16138 7790
rect 16248 7760 16288 7800
rect 16968 7730 17008 7770
rect 17358 7810 17398 7850
rect 14498 7300 14538 7340
rect 19798 7560 19838 7600
rect 20338 7550 20378 7590
rect 21418 7550 21458 7590
rect 21828 7520 21868 7560
rect 22088 7520 22128 7560
rect 13718 7180 13758 7220
rect 16838 7180 16878 7220
rect 15268 6960 15308 7000
rect 20218 6990 20258 7030
rect 20978 6990 21018 7030
rect 21388 7020 21428 7060
rect 22088 7020 22128 7060
rect 13598 6840 13638 6880
rect 13148 6380 13188 6420
rect 13478 6340 13518 6380
rect 14498 6840 14538 6880
rect 13998 6420 14038 6460
rect 14378 6340 14418 6380
rect 15048 6350 15088 6390
rect 15478 6390 15518 6430
rect 15808 6390 15848 6430
rect 16138 6390 16178 6430
rect 16268 6360 16308 6400
rect 16838 6390 16878 6430
rect 17358 6420 17398 6460
rect 17708 6420 17748 6460
rect 17228 6340 17268 6380
rect 19558 6450 19598 6490
rect 22398 6450 22438 6490
rect 15398 6000 15438 6040
rect 23408 4940 23448 4980
rect 23928 4940 23968 4980
rect 24448 4940 24488 4980
rect 24968 4940 25008 4980
rect 13038 3580 13078 3620
rect 13348 3560 13388 3600
rect 14158 3580 14198 3620
rect 14288 3580 14328 3620
rect 15418 3580 15458 3620
rect 17178 3590 17218 3630
rect 19708 3580 19748 3620
rect 21008 3580 21048 3620
rect 22308 3580 22348 3620
rect 12378 3460 12418 3500
rect 12508 3260 12548 3300
rect 13088 3260 13128 3300
rect 13628 3340 13668 3380
rect 13428 3260 13468 3300
rect 14028 3380 14068 3420
rect 14008 3260 14048 3300
rect 14528 3260 14568 3300
rect 14878 3260 14918 3300
rect 15728 3380 15768 3420
rect 15458 3260 15498 3300
rect 15668 3260 15708 3300
rect 15908 3260 15948 3300
rect 16248 3270 16288 3310
rect 16518 3310 16558 3350
rect 16718 3340 16758 3380
rect 17708 3460 17748 3500
rect 17118 3380 17158 3420
rect 17148 3260 17188 3300
rect 17508 3260 17548 3300
rect 17838 3260 17878 3300
rect 18248 3340 18288 3380
rect 18418 3260 18458 3300
rect 18888 3280 18928 3320
rect 19138 3170 19178 3210
rect 19548 3340 19588 3380
rect 19718 3170 19758 3210
rect 20188 3280 20228 3320
rect 20438 3170 20478 3210
rect 20848 3340 20888 3380
rect 21018 3170 21058 3210
rect 21488 3280 21528 3320
rect 21738 3170 21778 3210
rect 22148 3340 22188 3380
rect 23290 4058 23324 4092
rect 23810 4058 23844 4092
rect 24330 4058 24364 4092
rect 23262 3478 23296 3512
rect 23782 3478 23816 3512
rect 24302 3478 24336 3512
rect 22318 3170 22358 3210
rect 22762 3288 22796 3322
rect 12398 3020 12438 3060
rect 13348 3040 13388 3080
rect 14418 3030 14458 3070
rect 15978 3030 16018 3070
rect 18582 3020 18622 3060
rect 23262 3088 23296 3122
rect 23782 3088 23816 3122
rect 24302 3088 24336 3122
rect 23290 2708 23324 2742
rect 23810 2708 23844 2742
rect 24330 2708 24364 2742
rect 23276 2228 23310 2262
rect 23796 2228 23830 2262
rect 24316 2228 24350 2262
rect 24884 2228 24918 2262
<< xpolycontact >>
rect 14990 19436 15422 19506
rect 16894 19436 17326 19506
rect 8452 18026 8522 18458
rect 8452 17216 8522 17648
rect 9239 18029 9309 18461
rect 9571 16817 9641 17249
rect 10684 18026 10754 18458
rect 10352 16286 10422 16718
rect 15672 18026 15742 18458
rect 16004 16286 16074 16718
rect 16785 18023 16855 18455
rect 16785 17423 16855 17855
rect 17572 18026 17642 18458
rect 17572 17216 17642 17648
rect 12630 14540 13070 14610
rect 13498 14540 13938 14610
rect 23222 12716 23292 13148
rect 23222 12088 23292 12520
rect 23222 10196 23292 10628
rect 23222 9624 23292 10056
<< npolyres >>
rect 19672 9974 20152 10040
<< ppolyres >>
rect 8452 17648 8522 18026
rect 17572 17648 17642 18026
<< xpolyres >>
rect 15422 19436 16894 19506
rect 9239 17423 9309 18029
rect 9405 17855 9641 17925
rect 9405 17423 9475 17855
rect 9239 17353 9475 17423
rect 9571 17249 9641 17855
rect 10352 17852 10588 17922
rect 10352 16718 10422 17852
rect 10518 16892 10588 17852
rect 10684 16892 10754 18026
rect 10518 16822 10754 16892
rect 15672 16892 15742 18026
rect 15838 17852 16074 17922
rect 15838 16892 15908 17852
rect 15672 16822 15908 16892
rect 16004 16718 16074 17852
rect 16785 17855 16855 18023
rect 13070 14540 13498 14610
rect 23222 12520 23292 12716
rect 23222 10056 23292 10196
<< locali >>
rect 16118 19697 16198 19700
rect 14851 19663 14947 19697
rect 17369 19663 17465 19697
rect 14851 19601 14885 19663
rect 16118 19640 16138 19663
rect 16178 19640 16198 19663
rect 16118 19620 16198 19640
rect 17431 19601 17465 19663
rect 14851 19279 14885 19341
rect 17431 19279 17465 19341
rect 14851 19245 14947 19279
rect 17369 19245 17465 19279
rect 13238 19070 13318 19090
rect 13238 19030 13258 19070
rect 13298 19030 13318 19070
rect 13238 18990 13318 19030
rect 13238 18950 13258 18990
rect 13298 18950 13318 18990
rect 13238 18910 13318 18950
rect 13238 18870 13258 18910
rect 13298 18870 13318 18910
rect 12558 18784 12638 18790
rect 13238 18784 13318 18870
rect 13918 18784 13998 18790
rect 11274 18752 15282 18784
rect 11274 18718 11408 18752
rect 11442 18718 11498 18752
rect 11532 18718 11588 18752
rect 11622 18718 11678 18752
rect 11712 18718 11768 18752
rect 11802 18718 11858 18752
rect 11892 18718 11948 18752
rect 11982 18718 12038 18752
rect 12072 18718 12128 18752
rect 12162 18718 12218 18752
rect 12252 18718 12308 18752
rect 12342 18718 12398 18752
rect 12432 18718 12768 18752
rect 12802 18718 12858 18752
rect 12892 18718 12948 18752
rect 12982 18718 13038 18752
rect 13072 18718 13128 18752
rect 13162 18718 13218 18752
rect 13252 18718 13308 18752
rect 13342 18718 13398 18752
rect 13432 18718 13488 18752
rect 13522 18718 13578 18752
rect 13612 18718 13668 18752
rect 13702 18718 13758 18752
rect 13792 18718 14128 18752
rect 14162 18718 14218 18752
rect 14252 18718 14308 18752
rect 14342 18718 14398 18752
rect 14432 18718 14488 18752
rect 14522 18718 14578 18752
rect 14612 18718 14668 18752
rect 14702 18718 14758 18752
rect 14792 18718 14848 18752
rect 14882 18718 14938 18752
rect 14972 18718 15028 18752
rect 15062 18718 15118 18752
rect 15152 18718 15282 18752
rect 11274 18685 15282 18718
rect 11274 18668 11373 18685
rect 11274 18634 11307 18668
rect 11341 18634 11373 18668
rect 8448 18610 8528 18630
rect 8448 18597 8468 18610
rect 8508 18597 8528 18610
rect 9238 18610 9318 18630
rect 9238 18600 9258 18610
rect 9298 18600 9318 18610
rect 10678 18610 10758 18630
rect 8261 18563 8357 18597
rect 8617 18563 8713 18597
rect 8261 18501 8295 18563
rect 8448 18550 8528 18563
rect 8679 18501 8713 18563
rect 8261 17111 8295 17173
rect 8679 17111 8713 17173
rect 8261 17077 8357 17111
rect 8617 17077 8713 17111
rect 9048 18566 9144 18600
rect 9736 18566 9832 18600
rect 10678 18597 10698 18610
rect 10738 18597 10758 18610
rect 9048 18504 9082 18566
rect 9238 18550 9318 18566
rect 9798 18504 9832 18566
rect 9048 16712 9082 16774
rect 9798 16712 9832 16774
rect 9048 16678 9144 16712
rect 9736 16678 9832 16712
rect 10161 18563 10257 18597
rect 10849 18563 10945 18597
rect 10161 18501 10195 18563
rect 10678 18550 10758 18563
rect 10911 18501 10945 18563
rect 10161 16181 10195 16243
rect 11274 18578 11373 18634
rect 12463 18668 12733 18685
rect 12463 18634 12494 18668
rect 12528 18634 12667 18668
rect 12701 18634 12733 18668
rect 11274 18544 11307 18578
rect 11341 18544 11373 18578
rect 11274 18488 11373 18544
rect 11274 18454 11307 18488
rect 11341 18454 11373 18488
rect 11274 18398 11373 18454
rect 11274 18364 11307 18398
rect 11341 18364 11373 18398
rect 11274 18308 11373 18364
rect 11274 18274 11307 18308
rect 11341 18274 11373 18308
rect 11274 18218 11373 18274
rect 11274 18184 11307 18218
rect 11341 18184 11373 18218
rect 11274 18128 11373 18184
rect 11274 18094 11307 18128
rect 11341 18094 11373 18128
rect 11274 18038 11373 18094
rect 11274 18004 11307 18038
rect 11341 18004 11373 18038
rect 11274 17948 11373 18004
rect 11274 17914 11307 17948
rect 11341 17914 11373 17948
rect 11274 17858 11373 17914
rect 11274 17824 11307 17858
rect 11341 17824 11373 17858
rect 11274 17768 11373 17824
rect 11274 17740 11307 17768
rect 11268 17734 11307 17740
rect 11341 17740 11373 17768
rect 11437 18602 12399 18621
rect 11437 18568 11548 18602
rect 11582 18568 11638 18602
rect 11672 18568 11728 18602
rect 11762 18568 11818 18602
rect 11852 18568 11908 18602
rect 11942 18568 11998 18602
rect 12032 18568 12088 18602
rect 12122 18568 12178 18602
rect 12212 18568 12268 18602
rect 12302 18568 12399 18602
rect 11437 18549 12399 18568
rect 11437 18508 11509 18549
rect 11437 18474 11456 18508
rect 11490 18474 11509 18508
rect 12327 18489 12399 18549
rect 11437 18418 11509 18474
rect 11437 18384 11456 18418
rect 11490 18384 11509 18418
rect 11437 18328 11509 18384
rect 11437 18294 11456 18328
rect 11490 18294 11509 18328
rect 11437 18238 11509 18294
rect 11437 18204 11456 18238
rect 11490 18204 11509 18238
rect 11437 18148 11509 18204
rect 11437 18114 11456 18148
rect 11490 18114 11509 18148
rect 11437 18058 11509 18114
rect 11437 18024 11456 18058
rect 11490 18024 11509 18058
rect 11437 17968 11509 18024
rect 11437 17934 11456 17968
rect 11490 17934 11509 17968
rect 11437 17878 11509 17934
rect 11437 17844 11456 17878
rect 11490 17844 11509 17878
rect 11437 17788 11509 17844
rect 11571 18426 12265 18487
rect 11571 18392 11630 18426
rect 11664 18414 11720 18426
rect 11692 18392 11720 18414
rect 11754 18414 11810 18426
rect 11754 18392 11758 18414
rect 11571 18380 11658 18392
rect 11692 18380 11758 18392
rect 11792 18392 11810 18414
rect 11844 18414 11900 18426
rect 11844 18392 11858 18414
rect 11792 18380 11858 18392
rect 11892 18392 11900 18414
rect 11934 18414 11990 18426
rect 12024 18414 12080 18426
rect 12114 18414 12170 18426
rect 11934 18392 11958 18414
rect 12024 18392 12058 18414
rect 12114 18392 12158 18414
rect 12204 18392 12265 18426
rect 11892 18380 11958 18392
rect 11992 18380 12058 18392
rect 12092 18380 12158 18392
rect 12192 18380 12265 18392
rect 11571 18336 12265 18380
rect 11571 18302 11630 18336
rect 11664 18314 11720 18336
rect 11692 18302 11720 18314
rect 11754 18314 11810 18336
rect 11754 18302 11758 18314
rect 11571 18280 11658 18302
rect 11692 18280 11758 18302
rect 11792 18302 11810 18314
rect 11844 18314 11900 18336
rect 11844 18302 11858 18314
rect 11792 18280 11858 18302
rect 11892 18302 11900 18314
rect 11934 18314 11990 18336
rect 12024 18314 12080 18336
rect 12114 18314 12170 18336
rect 11934 18302 11958 18314
rect 12024 18302 12058 18314
rect 12114 18302 12158 18314
rect 12204 18302 12265 18336
rect 11892 18280 11958 18302
rect 11992 18280 12058 18302
rect 12092 18280 12158 18302
rect 12192 18280 12265 18302
rect 11571 18246 12265 18280
rect 11571 18212 11630 18246
rect 11664 18214 11720 18246
rect 11692 18212 11720 18214
rect 11754 18214 11810 18246
rect 11754 18212 11758 18214
rect 11571 18180 11658 18212
rect 11692 18180 11758 18212
rect 11792 18212 11810 18214
rect 11844 18214 11900 18246
rect 11844 18212 11858 18214
rect 11792 18180 11858 18212
rect 11892 18212 11900 18214
rect 11934 18214 11990 18246
rect 12024 18214 12080 18246
rect 12114 18214 12170 18246
rect 11934 18212 11958 18214
rect 12024 18212 12058 18214
rect 12114 18212 12158 18214
rect 12204 18212 12265 18246
rect 11892 18180 11958 18212
rect 11992 18180 12058 18212
rect 12092 18180 12158 18212
rect 12192 18180 12265 18212
rect 11571 18156 12265 18180
rect 11571 18122 11630 18156
rect 11664 18122 11720 18156
rect 11754 18122 11810 18156
rect 11844 18122 11900 18156
rect 11934 18122 11990 18156
rect 12024 18122 12080 18156
rect 12114 18122 12170 18156
rect 12204 18122 12265 18156
rect 11571 18114 12265 18122
rect 11571 18080 11658 18114
rect 11692 18080 11758 18114
rect 11792 18080 11858 18114
rect 11892 18080 11958 18114
rect 11992 18080 12058 18114
rect 12092 18080 12158 18114
rect 12192 18080 12265 18114
rect 11571 18066 12265 18080
rect 11571 18032 11630 18066
rect 11664 18032 11720 18066
rect 11754 18032 11810 18066
rect 11844 18032 11900 18066
rect 11934 18032 11990 18066
rect 12024 18032 12080 18066
rect 12114 18032 12170 18066
rect 12204 18032 12265 18066
rect 11571 18014 12265 18032
rect 11571 17980 11658 18014
rect 11692 17980 11758 18014
rect 11792 17980 11858 18014
rect 11892 17980 11958 18014
rect 11992 17980 12058 18014
rect 12092 17980 12158 18014
rect 12192 17980 12265 18014
rect 11571 17976 12265 17980
rect 11571 17942 11630 17976
rect 11664 17942 11720 17976
rect 11754 17942 11810 17976
rect 11844 17942 11900 17976
rect 11934 17942 11990 17976
rect 12024 17942 12080 17976
rect 12114 17942 12170 17976
rect 12204 17942 12265 17976
rect 11571 17914 12265 17942
rect 11571 17886 11658 17914
rect 11692 17886 11758 17914
rect 11571 17852 11630 17886
rect 11692 17880 11720 17886
rect 11664 17852 11720 17880
rect 11754 17880 11758 17886
rect 11792 17886 11858 17914
rect 11792 17880 11810 17886
rect 11754 17852 11810 17880
rect 11844 17880 11858 17886
rect 11892 17886 11958 17914
rect 11992 17886 12058 17914
rect 12092 17886 12158 17914
rect 12192 17886 12265 17914
rect 11892 17880 11900 17886
rect 11844 17852 11900 17880
rect 11934 17880 11958 17886
rect 12024 17880 12058 17886
rect 12114 17880 12158 17886
rect 11934 17852 11990 17880
rect 12024 17852 12080 17880
rect 12114 17852 12170 17880
rect 12204 17852 12265 17886
rect 11571 17793 12265 17852
rect 12327 18455 12346 18489
rect 12380 18455 12399 18489
rect 12327 18399 12399 18455
rect 12327 18365 12346 18399
rect 12380 18365 12399 18399
rect 12327 18309 12399 18365
rect 12327 18275 12346 18309
rect 12380 18275 12399 18309
rect 12327 18219 12399 18275
rect 12327 18185 12346 18219
rect 12380 18185 12399 18219
rect 12327 18129 12399 18185
rect 12327 18095 12346 18129
rect 12380 18095 12399 18129
rect 12327 18039 12399 18095
rect 12327 18005 12346 18039
rect 12380 18005 12399 18039
rect 12327 17949 12399 18005
rect 12327 17915 12346 17949
rect 12380 17915 12399 17949
rect 12327 17859 12399 17915
rect 12327 17825 12346 17859
rect 12380 17825 12399 17859
rect 11437 17754 11456 17788
rect 11490 17754 11509 17788
rect 11437 17740 11509 17754
rect 12327 17769 12399 17825
rect 12327 17740 12346 17769
rect 11341 17735 12346 17740
rect 12380 17740 12399 17769
rect 12463 18578 12733 18634
rect 13823 18668 14093 18685
rect 13823 18634 13854 18668
rect 13888 18634 14027 18668
rect 14061 18634 14093 18668
rect 12463 18544 12494 18578
rect 12528 18544 12667 18578
rect 12701 18544 12733 18578
rect 12463 18488 12733 18544
rect 12463 18454 12494 18488
rect 12528 18454 12667 18488
rect 12701 18454 12733 18488
rect 12463 18398 12733 18454
rect 12463 18364 12494 18398
rect 12528 18364 12667 18398
rect 12701 18364 12733 18398
rect 12463 18308 12733 18364
rect 12463 18274 12494 18308
rect 12528 18274 12667 18308
rect 12701 18274 12733 18308
rect 12463 18218 12733 18274
rect 12463 18184 12494 18218
rect 12528 18184 12667 18218
rect 12701 18184 12733 18218
rect 12463 18128 12733 18184
rect 12463 18094 12494 18128
rect 12528 18094 12667 18128
rect 12701 18094 12733 18128
rect 12463 18038 12733 18094
rect 12463 18004 12494 18038
rect 12528 18004 12667 18038
rect 12701 18004 12733 18038
rect 12463 17948 12733 18004
rect 12463 17914 12494 17948
rect 12528 17914 12667 17948
rect 12701 17914 12733 17948
rect 12463 17858 12733 17914
rect 12463 17824 12494 17858
rect 12528 17824 12667 17858
rect 12701 17824 12733 17858
rect 12463 17768 12733 17824
rect 12463 17740 12494 17768
rect 12380 17735 12494 17740
rect 11341 17734 12494 17735
rect 12528 17734 12667 17768
rect 12701 17740 12733 17768
rect 12797 18602 13759 18621
rect 12797 18568 12908 18602
rect 12942 18568 12998 18602
rect 13032 18568 13088 18602
rect 13122 18568 13178 18602
rect 13212 18568 13268 18602
rect 13302 18568 13358 18602
rect 13392 18568 13448 18602
rect 13482 18568 13538 18602
rect 13572 18568 13628 18602
rect 13662 18568 13759 18602
rect 12797 18549 13759 18568
rect 12797 18508 12869 18549
rect 12797 18474 12816 18508
rect 12850 18474 12869 18508
rect 13687 18489 13759 18549
rect 12797 18418 12869 18474
rect 12797 18384 12816 18418
rect 12850 18384 12869 18418
rect 12797 18328 12869 18384
rect 12797 18294 12816 18328
rect 12850 18294 12869 18328
rect 12797 18238 12869 18294
rect 12797 18204 12816 18238
rect 12850 18204 12869 18238
rect 12797 18148 12869 18204
rect 12797 18114 12816 18148
rect 12850 18114 12869 18148
rect 12797 18058 12869 18114
rect 12797 18024 12816 18058
rect 12850 18024 12869 18058
rect 12797 17968 12869 18024
rect 12797 17934 12816 17968
rect 12850 17934 12869 17968
rect 12797 17878 12869 17934
rect 12797 17844 12816 17878
rect 12850 17844 12869 17878
rect 12797 17788 12869 17844
rect 12931 18426 13625 18487
rect 12931 18392 12990 18426
rect 13024 18414 13080 18426
rect 13052 18392 13080 18414
rect 13114 18414 13170 18426
rect 13114 18392 13118 18414
rect 12931 18380 13018 18392
rect 13052 18380 13118 18392
rect 13152 18392 13170 18414
rect 13204 18414 13260 18426
rect 13204 18392 13218 18414
rect 13152 18380 13218 18392
rect 13252 18392 13260 18414
rect 13294 18414 13350 18426
rect 13384 18414 13440 18426
rect 13474 18414 13530 18426
rect 13294 18392 13318 18414
rect 13384 18392 13418 18414
rect 13474 18392 13518 18414
rect 13564 18392 13625 18426
rect 13252 18380 13318 18392
rect 13352 18380 13418 18392
rect 13452 18380 13518 18392
rect 13552 18380 13625 18392
rect 12931 18336 13625 18380
rect 12931 18302 12990 18336
rect 13024 18314 13080 18336
rect 13052 18302 13080 18314
rect 13114 18314 13170 18336
rect 13114 18302 13118 18314
rect 12931 18280 13018 18302
rect 13052 18280 13118 18302
rect 13152 18302 13170 18314
rect 13204 18314 13260 18336
rect 13204 18302 13218 18314
rect 13152 18280 13218 18302
rect 13252 18302 13260 18314
rect 13294 18314 13350 18336
rect 13384 18314 13440 18336
rect 13474 18314 13530 18336
rect 13294 18302 13318 18314
rect 13384 18302 13418 18314
rect 13474 18302 13518 18314
rect 13564 18302 13625 18336
rect 13252 18280 13318 18302
rect 13352 18280 13418 18302
rect 13452 18280 13518 18302
rect 13552 18280 13625 18302
rect 12931 18246 13625 18280
rect 12931 18212 12990 18246
rect 13024 18214 13080 18246
rect 13052 18212 13080 18214
rect 13114 18214 13170 18246
rect 13114 18212 13118 18214
rect 12931 18180 13018 18212
rect 13052 18180 13118 18212
rect 13152 18212 13170 18214
rect 13204 18214 13260 18246
rect 13204 18212 13218 18214
rect 13152 18180 13218 18212
rect 13252 18212 13260 18214
rect 13294 18214 13350 18246
rect 13384 18214 13440 18246
rect 13474 18214 13530 18246
rect 13294 18212 13318 18214
rect 13384 18212 13418 18214
rect 13474 18212 13518 18214
rect 13564 18212 13625 18246
rect 13252 18180 13318 18212
rect 13352 18180 13418 18212
rect 13452 18180 13518 18212
rect 13552 18180 13625 18212
rect 12931 18156 13625 18180
rect 12931 18122 12990 18156
rect 13024 18122 13080 18156
rect 13114 18122 13170 18156
rect 13204 18122 13260 18156
rect 13294 18122 13350 18156
rect 13384 18122 13440 18156
rect 13474 18122 13530 18156
rect 13564 18122 13625 18156
rect 12931 18114 13625 18122
rect 12931 18080 13018 18114
rect 13052 18080 13118 18114
rect 13152 18080 13218 18114
rect 13252 18080 13318 18114
rect 13352 18080 13418 18114
rect 13452 18080 13518 18114
rect 13552 18080 13625 18114
rect 12931 18066 13625 18080
rect 12931 18032 12990 18066
rect 13024 18032 13080 18066
rect 13114 18032 13170 18066
rect 13204 18032 13260 18066
rect 13294 18032 13350 18066
rect 13384 18032 13440 18066
rect 13474 18032 13530 18066
rect 13564 18032 13625 18066
rect 12931 18014 13625 18032
rect 12931 17980 13018 18014
rect 13052 17980 13118 18014
rect 13152 17980 13218 18014
rect 13252 17980 13318 18014
rect 13352 17980 13418 18014
rect 13452 17980 13518 18014
rect 13552 17980 13625 18014
rect 12931 17976 13625 17980
rect 12931 17942 12990 17976
rect 13024 17942 13080 17976
rect 13114 17942 13170 17976
rect 13204 17942 13260 17976
rect 13294 17942 13350 17976
rect 13384 17942 13440 17976
rect 13474 17942 13530 17976
rect 13564 17942 13625 17976
rect 12931 17914 13625 17942
rect 12931 17886 13018 17914
rect 13052 17886 13118 17914
rect 12931 17852 12990 17886
rect 13052 17880 13080 17886
rect 13024 17852 13080 17880
rect 13114 17880 13118 17886
rect 13152 17886 13218 17914
rect 13152 17880 13170 17886
rect 13114 17852 13170 17880
rect 13204 17880 13218 17886
rect 13252 17886 13318 17914
rect 13352 17886 13418 17914
rect 13452 17886 13518 17914
rect 13552 17886 13625 17914
rect 13252 17880 13260 17886
rect 13204 17852 13260 17880
rect 13294 17880 13318 17886
rect 13384 17880 13418 17886
rect 13474 17880 13518 17886
rect 13294 17852 13350 17880
rect 13384 17852 13440 17880
rect 13474 17852 13530 17880
rect 13564 17852 13625 17886
rect 12931 17793 13625 17852
rect 13687 18455 13706 18489
rect 13740 18455 13759 18489
rect 13687 18399 13759 18455
rect 13687 18365 13706 18399
rect 13740 18365 13759 18399
rect 13687 18309 13759 18365
rect 13687 18275 13706 18309
rect 13740 18275 13759 18309
rect 13687 18219 13759 18275
rect 13687 18185 13706 18219
rect 13740 18185 13759 18219
rect 13687 18129 13759 18185
rect 13687 18095 13706 18129
rect 13740 18095 13759 18129
rect 13687 18039 13759 18095
rect 13687 18005 13706 18039
rect 13740 18005 13759 18039
rect 13687 17949 13759 18005
rect 13687 17915 13706 17949
rect 13740 17915 13759 17949
rect 13687 17859 13759 17915
rect 13687 17825 13706 17859
rect 13740 17825 13759 17859
rect 12797 17754 12816 17788
rect 12850 17754 12869 17788
rect 12797 17740 12869 17754
rect 13687 17769 13759 17825
rect 13687 17740 13706 17769
rect 12701 17735 13706 17740
rect 13740 17740 13759 17769
rect 13823 18578 14093 18634
rect 15183 18668 15282 18685
rect 15183 18634 15214 18668
rect 15248 18634 15282 18668
rect 13823 18544 13854 18578
rect 13888 18544 14027 18578
rect 14061 18544 14093 18578
rect 13823 18488 14093 18544
rect 13823 18454 13854 18488
rect 13888 18454 14027 18488
rect 14061 18454 14093 18488
rect 13823 18398 14093 18454
rect 13823 18364 13854 18398
rect 13888 18364 14027 18398
rect 14061 18364 14093 18398
rect 13823 18308 14093 18364
rect 13823 18274 13854 18308
rect 13888 18274 14027 18308
rect 14061 18274 14093 18308
rect 13823 18218 14093 18274
rect 13823 18184 13854 18218
rect 13888 18184 14027 18218
rect 14061 18184 14093 18218
rect 13823 18128 14093 18184
rect 13823 18094 13854 18128
rect 13888 18094 14027 18128
rect 14061 18094 14093 18128
rect 13823 18038 14093 18094
rect 13823 18004 13854 18038
rect 13888 18004 14027 18038
rect 14061 18004 14093 18038
rect 13823 17948 14093 18004
rect 13823 17914 13854 17948
rect 13888 17914 14027 17948
rect 14061 17914 14093 17948
rect 13823 17858 14093 17914
rect 13823 17824 13854 17858
rect 13888 17824 14027 17858
rect 14061 17824 14093 17858
rect 13823 17768 14093 17824
rect 13823 17740 13854 17768
rect 13740 17735 13854 17740
rect 12701 17734 13854 17735
rect 13888 17734 14027 17768
rect 14061 17740 14093 17768
rect 14157 18602 15119 18621
rect 14157 18568 14268 18602
rect 14302 18568 14358 18602
rect 14392 18568 14448 18602
rect 14482 18568 14538 18602
rect 14572 18568 14628 18602
rect 14662 18568 14718 18602
rect 14752 18568 14808 18602
rect 14842 18568 14898 18602
rect 14932 18568 14988 18602
rect 15022 18568 15119 18602
rect 14157 18549 15119 18568
rect 14157 18508 14229 18549
rect 14157 18474 14176 18508
rect 14210 18474 14229 18508
rect 15047 18489 15119 18549
rect 14157 18418 14229 18474
rect 14157 18384 14176 18418
rect 14210 18384 14229 18418
rect 14157 18328 14229 18384
rect 14157 18294 14176 18328
rect 14210 18294 14229 18328
rect 14157 18238 14229 18294
rect 14157 18204 14176 18238
rect 14210 18204 14229 18238
rect 14157 18148 14229 18204
rect 14157 18114 14176 18148
rect 14210 18114 14229 18148
rect 14157 18058 14229 18114
rect 14157 18024 14176 18058
rect 14210 18024 14229 18058
rect 14157 17968 14229 18024
rect 14157 17934 14176 17968
rect 14210 17934 14229 17968
rect 14157 17878 14229 17934
rect 14157 17844 14176 17878
rect 14210 17844 14229 17878
rect 14157 17788 14229 17844
rect 14291 18426 14985 18487
rect 14291 18392 14350 18426
rect 14384 18414 14440 18426
rect 14412 18392 14440 18414
rect 14474 18414 14530 18426
rect 14474 18392 14478 18414
rect 14291 18380 14378 18392
rect 14412 18380 14478 18392
rect 14512 18392 14530 18414
rect 14564 18414 14620 18426
rect 14564 18392 14578 18414
rect 14512 18380 14578 18392
rect 14612 18392 14620 18414
rect 14654 18414 14710 18426
rect 14744 18414 14800 18426
rect 14834 18414 14890 18426
rect 14654 18392 14678 18414
rect 14744 18392 14778 18414
rect 14834 18392 14878 18414
rect 14924 18392 14985 18426
rect 14612 18380 14678 18392
rect 14712 18380 14778 18392
rect 14812 18380 14878 18392
rect 14912 18380 14985 18392
rect 14291 18336 14985 18380
rect 14291 18302 14350 18336
rect 14384 18314 14440 18336
rect 14412 18302 14440 18314
rect 14474 18314 14530 18336
rect 14474 18302 14478 18314
rect 14291 18280 14378 18302
rect 14412 18280 14478 18302
rect 14512 18302 14530 18314
rect 14564 18314 14620 18336
rect 14564 18302 14578 18314
rect 14512 18280 14578 18302
rect 14612 18302 14620 18314
rect 14654 18314 14710 18336
rect 14744 18314 14800 18336
rect 14834 18314 14890 18336
rect 14654 18302 14678 18314
rect 14744 18302 14778 18314
rect 14834 18302 14878 18314
rect 14924 18302 14985 18336
rect 14612 18280 14678 18302
rect 14712 18280 14778 18302
rect 14812 18280 14878 18302
rect 14912 18280 14985 18302
rect 14291 18246 14985 18280
rect 14291 18212 14350 18246
rect 14384 18214 14440 18246
rect 14412 18212 14440 18214
rect 14474 18214 14530 18246
rect 14474 18212 14478 18214
rect 14291 18180 14378 18212
rect 14412 18180 14478 18212
rect 14512 18212 14530 18214
rect 14564 18214 14620 18246
rect 14564 18212 14578 18214
rect 14512 18180 14578 18212
rect 14612 18212 14620 18214
rect 14654 18214 14710 18246
rect 14744 18214 14800 18246
rect 14834 18214 14890 18246
rect 14654 18212 14678 18214
rect 14744 18212 14778 18214
rect 14834 18212 14878 18214
rect 14924 18212 14985 18246
rect 14612 18180 14678 18212
rect 14712 18180 14778 18212
rect 14812 18180 14878 18212
rect 14912 18180 14985 18212
rect 14291 18156 14985 18180
rect 14291 18122 14350 18156
rect 14384 18122 14440 18156
rect 14474 18122 14530 18156
rect 14564 18122 14620 18156
rect 14654 18122 14710 18156
rect 14744 18122 14800 18156
rect 14834 18122 14890 18156
rect 14924 18122 14985 18156
rect 14291 18114 14985 18122
rect 14291 18080 14378 18114
rect 14412 18080 14478 18114
rect 14512 18080 14578 18114
rect 14612 18080 14678 18114
rect 14712 18080 14778 18114
rect 14812 18080 14878 18114
rect 14912 18080 14985 18114
rect 14291 18066 14985 18080
rect 14291 18032 14350 18066
rect 14384 18032 14440 18066
rect 14474 18032 14530 18066
rect 14564 18032 14620 18066
rect 14654 18032 14710 18066
rect 14744 18032 14800 18066
rect 14834 18032 14890 18066
rect 14924 18032 14985 18066
rect 14291 18014 14985 18032
rect 14291 17980 14378 18014
rect 14412 17980 14478 18014
rect 14512 17980 14578 18014
rect 14612 17980 14678 18014
rect 14712 17980 14778 18014
rect 14812 17980 14878 18014
rect 14912 17980 14985 18014
rect 14291 17976 14985 17980
rect 14291 17942 14350 17976
rect 14384 17942 14440 17976
rect 14474 17942 14530 17976
rect 14564 17942 14620 17976
rect 14654 17942 14710 17976
rect 14744 17942 14800 17976
rect 14834 17942 14890 17976
rect 14924 17942 14985 17976
rect 14291 17914 14985 17942
rect 14291 17886 14378 17914
rect 14412 17886 14478 17914
rect 14291 17852 14350 17886
rect 14412 17880 14440 17886
rect 14384 17852 14440 17880
rect 14474 17880 14478 17886
rect 14512 17886 14578 17914
rect 14512 17880 14530 17886
rect 14474 17852 14530 17880
rect 14564 17880 14578 17886
rect 14612 17886 14678 17914
rect 14712 17886 14778 17914
rect 14812 17886 14878 17914
rect 14912 17886 14985 17914
rect 14612 17880 14620 17886
rect 14564 17852 14620 17880
rect 14654 17880 14678 17886
rect 14744 17880 14778 17886
rect 14834 17880 14878 17886
rect 14654 17852 14710 17880
rect 14744 17852 14800 17880
rect 14834 17852 14890 17880
rect 14924 17852 14985 17886
rect 14291 17793 14985 17852
rect 15047 18455 15066 18489
rect 15100 18455 15119 18489
rect 15047 18399 15119 18455
rect 15047 18365 15066 18399
rect 15100 18365 15119 18399
rect 15047 18309 15119 18365
rect 15047 18275 15066 18309
rect 15100 18275 15119 18309
rect 15047 18219 15119 18275
rect 15047 18185 15066 18219
rect 15100 18185 15119 18219
rect 15047 18129 15119 18185
rect 15047 18095 15066 18129
rect 15100 18095 15119 18129
rect 15047 18039 15119 18095
rect 15047 18005 15066 18039
rect 15100 18005 15119 18039
rect 15047 17949 15119 18005
rect 15047 17915 15066 17949
rect 15100 17915 15119 17949
rect 15047 17859 15119 17915
rect 15047 17825 15066 17859
rect 15100 17825 15119 17859
rect 14157 17754 14176 17788
rect 14210 17754 14229 17788
rect 14157 17740 14229 17754
rect 15047 17769 15119 17825
rect 15047 17740 15066 17769
rect 14061 17735 15066 17740
rect 15100 17740 15119 17769
rect 15183 18578 15282 18634
rect 15668 18610 15748 18630
rect 15668 18597 15688 18610
rect 15728 18597 15748 18610
rect 16778 18610 16858 18630
rect 15183 18544 15214 18578
rect 15248 18544 15282 18578
rect 15183 18488 15282 18544
rect 15183 18454 15214 18488
rect 15248 18454 15282 18488
rect 15183 18398 15282 18454
rect 15183 18364 15214 18398
rect 15248 18364 15282 18398
rect 15183 18308 15282 18364
rect 15183 18274 15214 18308
rect 15248 18274 15282 18308
rect 15183 18218 15282 18274
rect 15183 18184 15214 18218
rect 15248 18184 15282 18218
rect 15183 18128 15282 18184
rect 15183 18094 15214 18128
rect 15248 18094 15282 18128
rect 15183 18038 15282 18094
rect 15183 18004 15214 18038
rect 15248 18004 15282 18038
rect 15183 17948 15282 18004
rect 15183 17914 15214 17948
rect 15248 17914 15282 17948
rect 15183 17858 15282 17914
rect 15183 17824 15214 17858
rect 15248 17824 15282 17858
rect 15183 17768 15282 17824
rect 15183 17740 15214 17768
rect 15100 17735 15214 17740
rect 14061 17734 15214 17735
rect 15248 17740 15282 17768
rect 15481 18563 15577 18597
rect 16169 18563 16265 18597
rect 16778 18594 16798 18610
rect 16838 18594 16858 18610
rect 17568 18610 17648 18630
rect 17568 18597 17588 18610
rect 17628 18597 17648 18610
rect 15481 18501 15515 18563
rect 15668 18550 15748 18563
rect 15248 17734 15288 17740
rect 11268 17712 15288 17734
rect 11268 17678 11514 17712
rect 11548 17678 11604 17712
rect 11638 17678 11694 17712
rect 11728 17678 11784 17712
rect 11818 17678 11874 17712
rect 11908 17678 11964 17712
rect 11998 17678 12054 17712
rect 12088 17678 12144 17712
rect 12178 17678 12234 17712
rect 12268 17678 12874 17712
rect 12908 17678 12964 17712
rect 12998 17678 13054 17712
rect 13088 17678 13144 17712
rect 13178 17678 13234 17712
rect 13268 17678 13324 17712
rect 13358 17678 13414 17712
rect 13448 17678 13504 17712
rect 13538 17678 13594 17712
rect 13628 17678 14234 17712
rect 14268 17678 14324 17712
rect 14358 17678 14414 17712
rect 14448 17678 14504 17712
rect 14538 17678 14594 17712
rect 14628 17678 14684 17712
rect 14718 17678 14774 17712
rect 14808 17678 14864 17712
rect 14898 17678 14954 17712
rect 14988 17678 15288 17712
rect 11268 17644 11307 17678
rect 11341 17644 12494 17678
rect 12528 17644 12667 17678
rect 12701 17644 13854 17678
rect 13888 17644 14027 17678
rect 14061 17644 15214 17678
rect 15248 17644 15288 17678
rect 11268 17588 15288 17644
rect 11268 17554 11307 17588
rect 11341 17565 12494 17588
rect 11341 17554 11408 17565
rect 11268 17531 11408 17554
rect 11442 17531 11498 17565
rect 11532 17531 11588 17565
rect 11622 17531 11678 17565
rect 11712 17531 11768 17565
rect 11802 17531 11858 17565
rect 11892 17531 11948 17565
rect 11982 17531 12038 17565
rect 12072 17531 12128 17565
rect 12162 17531 12218 17565
rect 12252 17531 12308 17565
rect 12342 17531 12398 17565
rect 12432 17554 12494 17565
rect 12528 17554 12667 17588
rect 12701 17565 13854 17588
rect 12701 17554 12768 17565
rect 12432 17531 12768 17554
rect 12802 17531 12858 17565
rect 12892 17531 12948 17565
rect 12982 17531 13038 17565
rect 13072 17531 13128 17565
rect 13162 17531 13218 17565
rect 13252 17531 13308 17565
rect 13342 17531 13398 17565
rect 13432 17531 13488 17565
rect 13522 17531 13578 17565
rect 13612 17531 13668 17565
rect 13702 17531 13758 17565
rect 13792 17554 13854 17565
rect 13888 17554 14027 17588
rect 14061 17565 15214 17588
rect 14061 17554 14128 17565
rect 13792 17531 14128 17554
rect 14162 17531 14218 17565
rect 14252 17531 14308 17565
rect 14342 17531 14398 17565
rect 14432 17531 14488 17565
rect 14522 17531 14578 17565
rect 14612 17531 14668 17565
rect 14702 17531 14758 17565
rect 14792 17531 14848 17565
rect 14882 17531 14938 17565
rect 14972 17531 15028 17565
rect 15062 17531 15118 17565
rect 15152 17554 15214 17565
rect 15248 17554 15288 17588
rect 15152 17531 15288 17554
rect 11268 17490 15288 17531
rect 12558 17424 12638 17490
rect 13918 17424 13998 17490
rect 11274 17392 15282 17424
rect 11274 17358 11408 17392
rect 11442 17358 11498 17392
rect 11532 17358 11588 17392
rect 11622 17358 11678 17392
rect 11712 17358 11768 17392
rect 11802 17358 11858 17392
rect 11892 17358 11948 17392
rect 11982 17358 12038 17392
rect 12072 17358 12128 17392
rect 12162 17358 12218 17392
rect 12252 17358 12308 17392
rect 12342 17358 12398 17392
rect 12432 17358 12768 17392
rect 12802 17358 12858 17392
rect 12892 17358 12948 17392
rect 12982 17358 13038 17392
rect 13072 17358 13128 17392
rect 13162 17358 13218 17392
rect 13252 17358 13308 17392
rect 13342 17358 13398 17392
rect 13432 17358 13488 17392
rect 13522 17358 13578 17392
rect 13612 17358 13668 17392
rect 13702 17358 13758 17392
rect 13792 17358 14128 17392
rect 14162 17358 14218 17392
rect 14252 17358 14308 17392
rect 14342 17358 14398 17392
rect 14432 17358 14488 17392
rect 14522 17358 14578 17392
rect 14612 17358 14668 17392
rect 14702 17358 14758 17392
rect 14792 17358 14848 17392
rect 14882 17358 14938 17392
rect 14972 17358 15028 17392
rect 15062 17358 15118 17392
rect 15152 17358 15282 17392
rect 11274 17325 15282 17358
rect 11274 17308 11373 17325
rect 11274 17274 11307 17308
rect 11341 17274 11373 17308
rect 11274 17218 11373 17274
rect 12463 17308 12733 17325
rect 12463 17274 12494 17308
rect 12528 17274 12667 17308
rect 12701 17274 12733 17308
rect 11274 17184 11307 17218
rect 11341 17184 11373 17218
rect 11274 17128 11373 17184
rect 11274 17094 11307 17128
rect 11341 17094 11373 17128
rect 11274 17038 11373 17094
rect 11274 17004 11307 17038
rect 11341 17004 11373 17038
rect 11274 16948 11373 17004
rect 11274 16914 11307 16948
rect 11341 16914 11373 16948
rect 11274 16858 11373 16914
rect 11274 16824 11307 16858
rect 11341 16824 11373 16858
rect 11274 16768 11373 16824
rect 11274 16734 11307 16768
rect 11341 16734 11373 16768
rect 11274 16678 11373 16734
rect 11274 16644 11307 16678
rect 11341 16644 11373 16678
rect 11274 16588 11373 16644
rect 11274 16554 11307 16588
rect 11341 16554 11373 16588
rect 11274 16498 11373 16554
rect 11274 16464 11307 16498
rect 11341 16464 11373 16498
rect 11274 16408 11373 16464
rect 11274 16380 11307 16408
rect 10911 16181 10945 16243
rect 10161 16147 10257 16181
rect 10849 16147 10945 16181
rect 11268 16374 11307 16380
rect 11341 16380 11373 16408
rect 11437 17242 12399 17261
rect 11437 17208 11548 17242
rect 11582 17208 11638 17242
rect 11672 17208 11728 17242
rect 11762 17208 11818 17242
rect 11852 17208 11908 17242
rect 11942 17208 11998 17242
rect 12032 17208 12088 17242
rect 12122 17208 12178 17242
rect 12212 17208 12268 17242
rect 12302 17208 12399 17242
rect 11437 17189 12399 17208
rect 11437 17148 11509 17189
rect 11437 17114 11456 17148
rect 11490 17114 11509 17148
rect 12327 17129 12399 17189
rect 11437 17058 11509 17114
rect 11437 17024 11456 17058
rect 11490 17024 11509 17058
rect 11437 16968 11509 17024
rect 11437 16934 11456 16968
rect 11490 16934 11509 16968
rect 11437 16878 11509 16934
rect 11437 16844 11456 16878
rect 11490 16844 11509 16878
rect 11437 16788 11509 16844
rect 11437 16754 11456 16788
rect 11490 16754 11509 16788
rect 11437 16698 11509 16754
rect 11437 16664 11456 16698
rect 11490 16664 11509 16698
rect 11437 16608 11509 16664
rect 11437 16574 11456 16608
rect 11490 16574 11509 16608
rect 11437 16518 11509 16574
rect 11437 16484 11456 16518
rect 11490 16484 11509 16518
rect 11437 16428 11509 16484
rect 11571 17066 12265 17127
rect 11571 17032 11630 17066
rect 11664 17054 11720 17066
rect 11692 17032 11720 17054
rect 11754 17054 11810 17066
rect 11754 17032 11758 17054
rect 11571 17020 11658 17032
rect 11692 17020 11758 17032
rect 11792 17032 11810 17054
rect 11844 17054 11900 17066
rect 11844 17032 11858 17054
rect 11792 17020 11858 17032
rect 11892 17032 11900 17054
rect 11934 17054 11990 17066
rect 12024 17054 12080 17066
rect 12114 17054 12170 17066
rect 11934 17032 11958 17054
rect 12024 17032 12058 17054
rect 12114 17032 12158 17054
rect 12204 17032 12265 17066
rect 11892 17020 11958 17032
rect 11992 17020 12058 17032
rect 12092 17020 12158 17032
rect 12192 17020 12265 17032
rect 11571 16976 12265 17020
rect 11571 16942 11630 16976
rect 11664 16954 11720 16976
rect 11692 16942 11720 16954
rect 11754 16954 11810 16976
rect 11754 16942 11758 16954
rect 11571 16920 11658 16942
rect 11692 16920 11758 16942
rect 11792 16942 11810 16954
rect 11844 16954 11900 16976
rect 11844 16942 11858 16954
rect 11792 16920 11858 16942
rect 11892 16942 11900 16954
rect 11934 16954 11990 16976
rect 12024 16954 12080 16976
rect 12114 16954 12170 16976
rect 11934 16942 11958 16954
rect 12024 16942 12058 16954
rect 12114 16942 12158 16954
rect 12204 16942 12265 16976
rect 11892 16920 11958 16942
rect 11992 16920 12058 16942
rect 12092 16920 12158 16942
rect 12192 16920 12265 16942
rect 11571 16886 12265 16920
rect 11571 16852 11630 16886
rect 11664 16854 11720 16886
rect 11692 16852 11720 16854
rect 11754 16854 11810 16886
rect 11754 16852 11758 16854
rect 11571 16820 11658 16852
rect 11692 16820 11758 16852
rect 11792 16852 11810 16854
rect 11844 16854 11900 16886
rect 11844 16852 11858 16854
rect 11792 16820 11858 16852
rect 11892 16852 11900 16854
rect 11934 16854 11990 16886
rect 12024 16854 12080 16886
rect 12114 16854 12170 16886
rect 11934 16852 11958 16854
rect 12024 16852 12058 16854
rect 12114 16852 12158 16854
rect 12204 16852 12265 16886
rect 11892 16820 11958 16852
rect 11992 16820 12058 16852
rect 12092 16820 12158 16852
rect 12192 16820 12265 16852
rect 11571 16796 12265 16820
rect 11571 16762 11630 16796
rect 11664 16762 11720 16796
rect 11754 16762 11810 16796
rect 11844 16762 11900 16796
rect 11934 16762 11990 16796
rect 12024 16762 12080 16796
rect 12114 16762 12170 16796
rect 12204 16762 12265 16796
rect 11571 16754 12265 16762
rect 11571 16720 11658 16754
rect 11692 16720 11758 16754
rect 11792 16720 11858 16754
rect 11892 16720 11958 16754
rect 11992 16720 12058 16754
rect 12092 16720 12158 16754
rect 12192 16720 12265 16754
rect 11571 16706 12265 16720
rect 11571 16672 11630 16706
rect 11664 16672 11720 16706
rect 11754 16672 11810 16706
rect 11844 16672 11900 16706
rect 11934 16672 11990 16706
rect 12024 16672 12080 16706
rect 12114 16672 12170 16706
rect 12204 16672 12265 16706
rect 11571 16654 12265 16672
rect 11571 16620 11658 16654
rect 11692 16620 11758 16654
rect 11792 16620 11858 16654
rect 11892 16620 11958 16654
rect 11992 16620 12058 16654
rect 12092 16620 12158 16654
rect 12192 16620 12265 16654
rect 11571 16616 12265 16620
rect 11571 16582 11630 16616
rect 11664 16582 11720 16616
rect 11754 16582 11810 16616
rect 11844 16582 11900 16616
rect 11934 16582 11990 16616
rect 12024 16582 12080 16616
rect 12114 16582 12170 16616
rect 12204 16582 12265 16616
rect 11571 16554 12265 16582
rect 11571 16526 11658 16554
rect 11692 16526 11758 16554
rect 11571 16492 11630 16526
rect 11692 16520 11720 16526
rect 11664 16492 11720 16520
rect 11754 16520 11758 16526
rect 11792 16526 11858 16554
rect 11792 16520 11810 16526
rect 11754 16492 11810 16520
rect 11844 16520 11858 16526
rect 11892 16526 11958 16554
rect 11992 16526 12058 16554
rect 12092 16526 12158 16554
rect 12192 16526 12265 16554
rect 11892 16520 11900 16526
rect 11844 16492 11900 16520
rect 11934 16520 11958 16526
rect 12024 16520 12058 16526
rect 12114 16520 12158 16526
rect 11934 16492 11990 16520
rect 12024 16492 12080 16520
rect 12114 16492 12170 16520
rect 12204 16492 12265 16526
rect 11571 16433 12265 16492
rect 12327 17095 12346 17129
rect 12380 17095 12399 17129
rect 12327 17039 12399 17095
rect 12327 17005 12346 17039
rect 12380 17005 12399 17039
rect 12327 16949 12399 17005
rect 12327 16915 12346 16949
rect 12380 16915 12399 16949
rect 12327 16859 12399 16915
rect 12327 16825 12346 16859
rect 12380 16825 12399 16859
rect 12327 16769 12399 16825
rect 12327 16735 12346 16769
rect 12380 16735 12399 16769
rect 12327 16679 12399 16735
rect 12327 16645 12346 16679
rect 12380 16645 12399 16679
rect 12327 16589 12399 16645
rect 12327 16555 12346 16589
rect 12380 16555 12399 16589
rect 12327 16499 12399 16555
rect 12327 16465 12346 16499
rect 12380 16465 12399 16499
rect 11437 16394 11456 16428
rect 11490 16394 11509 16428
rect 11437 16380 11509 16394
rect 12327 16409 12399 16465
rect 12327 16380 12346 16409
rect 11341 16375 12346 16380
rect 12380 16380 12399 16409
rect 12463 17218 12733 17274
rect 13823 17308 14093 17325
rect 13823 17274 13854 17308
rect 13888 17274 14027 17308
rect 14061 17274 14093 17308
rect 12463 17184 12494 17218
rect 12528 17184 12667 17218
rect 12701 17184 12733 17218
rect 12463 17128 12733 17184
rect 12463 17094 12494 17128
rect 12528 17094 12667 17128
rect 12701 17094 12733 17128
rect 12463 17038 12733 17094
rect 12463 17004 12494 17038
rect 12528 17004 12667 17038
rect 12701 17004 12733 17038
rect 12463 16948 12733 17004
rect 12463 16914 12494 16948
rect 12528 16914 12667 16948
rect 12701 16914 12733 16948
rect 12463 16858 12733 16914
rect 12463 16824 12494 16858
rect 12528 16824 12667 16858
rect 12701 16824 12733 16858
rect 12463 16768 12733 16824
rect 12463 16734 12494 16768
rect 12528 16734 12667 16768
rect 12701 16734 12733 16768
rect 12463 16678 12733 16734
rect 12463 16644 12494 16678
rect 12528 16644 12667 16678
rect 12701 16644 12733 16678
rect 12463 16588 12733 16644
rect 12463 16554 12494 16588
rect 12528 16554 12667 16588
rect 12701 16554 12733 16588
rect 12463 16498 12733 16554
rect 12463 16464 12494 16498
rect 12528 16464 12667 16498
rect 12701 16464 12733 16498
rect 12463 16408 12733 16464
rect 12463 16380 12494 16408
rect 12380 16375 12494 16380
rect 11341 16374 12494 16375
rect 12528 16374 12667 16408
rect 12701 16380 12733 16408
rect 12797 17242 13759 17261
rect 12797 17208 12908 17242
rect 12942 17208 12998 17242
rect 13032 17208 13088 17242
rect 13122 17208 13178 17242
rect 13212 17208 13268 17242
rect 13302 17208 13358 17242
rect 13392 17208 13448 17242
rect 13482 17208 13538 17242
rect 13572 17208 13628 17242
rect 13662 17208 13759 17242
rect 12797 17189 13759 17208
rect 12797 17148 12869 17189
rect 12797 17114 12816 17148
rect 12850 17114 12869 17148
rect 13687 17129 13759 17189
rect 12797 17058 12869 17114
rect 12797 17024 12816 17058
rect 12850 17024 12869 17058
rect 12797 16968 12869 17024
rect 12797 16934 12816 16968
rect 12850 16934 12869 16968
rect 12797 16878 12869 16934
rect 12797 16844 12816 16878
rect 12850 16844 12869 16878
rect 12797 16788 12869 16844
rect 12797 16754 12816 16788
rect 12850 16754 12869 16788
rect 12797 16698 12869 16754
rect 12797 16664 12816 16698
rect 12850 16664 12869 16698
rect 12797 16608 12869 16664
rect 12797 16574 12816 16608
rect 12850 16574 12869 16608
rect 12797 16518 12869 16574
rect 12797 16484 12816 16518
rect 12850 16484 12869 16518
rect 12797 16428 12869 16484
rect 12931 17066 13625 17127
rect 12931 17032 12990 17066
rect 13024 17054 13080 17066
rect 13052 17032 13080 17054
rect 13114 17054 13170 17066
rect 13114 17032 13118 17054
rect 12931 17020 13018 17032
rect 13052 17020 13118 17032
rect 13152 17032 13170 17054
rect 13204 17054 13260 17066
rect 13204 17032 13218 17054
rect 13152 17020 13218 17032
rect 13252 17032 13260 17054
rect 13294 17054 13350 17066
rect 13384 17054 13440 17066
rect 13474 17054 13530 17066
rect 13294 17032 13318 17054
rect 13384 17032 13418 17054
rect 13474 17032 13518 17054
rect 13564 17032 13625 17066
rect 13252 17020 13318 17032
rect 13352 17020 13418 17032
rect 13452 17020 13518 17032
rect 13552 17020 13625 17032
rect 12931 16976 13625 17020
rect 12931 16942 12990 16976
rect 13024 16954 13080 16976
rect 13052 16942 13080 16954
rect 13114 16954 13170 16976
rect 13114 16942 13118 16954
rect 12931 16920 13018 16942
rect 13052 16920 13118 16942
rect 13152 16942 13170 16954
rect 13204 16954 13260 16976
rect 13204 16942 13218 16954
rect 13152 16920 13218 16942
rect 13252 16942 13260 16954
rect 13294 16954 13350 16976
rect 13384 16954 13440 16976
rect 13474 16954 13530 16976
rect 13294 16942 13318 16954
rect 13384 16942 13418 16954
rect 13474 16942 13518 16954
rect 13564 16942 13625 16976
rect 13252 16920 13318 16942
rect 13352 16920 13418 16942
rect 13452 16920 13518 16942
rect 13552 16920 13625 16942
rect 12931 16886 13625 16920
rect 12931 16852 12990 16886
rect 13024 16854 13080 16886
rect 13052 16852 13080 16854
rect 13114 16854 13170 16886
rect 13114 16852 13118 16854
rect 12931 16820 13018 16852
rect 13052 16820 13118 16852
rect 13152 16852 13170 16854
rect 13204 16854 13260 16886
rect 13204 16852 13218 16854
rect 13152 16820 13218 16852
rect 13252 16852 13260 16854
rect 13294 16854 13350 16886
rect 13384 16854 13440 16886
rect 13474 16854 13530 16886
rect 13294 16852 13318 16854
rect 13384 16852 13418 16854
rect 13474 16852 13518 16854
rect 13564 16852 13625 16886
rect 13252 16820 13318 16852
rect 13352 16820 13418 16852
rect 13452 16820 13518 16852
rect 13552 16820 13625 16852
rect 12931 16796 13625 16820
rect 12931 16762 12990 16796
rect 13024 16762 13080 16796
rect 13114 16762 13170 16796
rect 13204 16762 13260 16796
rect 13294 16762 13350 16796
rect 13384 16762 13440 16796
rect 13474 16762 13530 16796
rect 13564 16762 13625 16796
rect 12931 16754 13625 16762
rect 12931 16720 13018 16754
rect 13052 16720 13118 16754
rect 13152 16720 13218 16754
rect 13252 16720 13318 16754
rect 13352 16720 13418 16754
rect 13452 16720 13518 16754
rect 13552 16720 13625 16754
rect 12931 16706 13625 16720
rect 12931 16672 12990 16706
rect 13024 16672 13080 16706
rect 13114 16672 13170 16706
rect 13204 16672 13260 16706
rect 13294 16672 13350 16706
rect 13384 16672 13440 16706
rect 13474 16672 13530 16706
rect 13564 16672 13625 16706
rect 12931 16654 13625 16672
rect 12931 16620 13018 16654
rect 13052 16620 13118 16654
rect 13152 16620 13218 16654
rect 13252 16620 13318 16654
rect 13352 16620 13418 16654
rect 13452 16620 13518 16654
rect 13552 16620 13625 16654
rect 12931 16616 13625 16620
rect 12931 16582 12990 16616
rect 13024 16582 13080 16616
rect 13114 16582 13170 16616
rect 13204 16582 13260 16616
rect 13294 16582 13350 16616
rect 13384 16582 13440 16616
rect 13474 16582 13530 16616
rect 13564 16582 13625 16616
rect 12931 16554 13625 16582
rect 12931 16526 13018 16554
rect 13052 16526 13118 16554
rect 12931 16492 12990 16526
rect 13052 16520 13080 16526
rect 13024 16492 13080 16520
rect 13114 16520 13118 16526
rect 13152 16526 13218 16554
rect 13152 16520 13170 16526
rect 13114 16492 13170 16520
rect 13204 16520 13218 16526
rect 13252 16526 13318 16554
rect 13352 16526 13418 16554
rect 13452 16526 13518 16554
rect 13552 16526 13625 16554
rect 13252 16520 13260 16526
rect 13204 16492 13260 16520
rect 13294 16520 13318 16526
rect 13384 16520 13418 16526
rect 13474 16520 13518 16526
rect 13294 16492 13350 16520
rect 13384 16492 13440 16520
rect 13474 16492 13530 16520
rect 13564 16492 13625 16526
rect 12931 16433 13625 16492
rect 13687 17095 13706 17129
rect 13740 17095 13759 17129
rect 13687 17039 13759 17095
rect 13687 17005 13706 17039
rect 13740 17005 13759 17039
rect 13687 16949 13759 17005
rect 13687 16915 13706 16949
rect 13740 16915 13759 16949
rect 13687 16859 13759 16915
rect 13687 16825 13706 16859
rect 13740 16825 13759 16859
rect 13687 16769 13759 16825
rect 13687 16735 13706 16769
rect 13740 16735 13759 16769
rect 13687 16679 13759 16735
rect 13687 16645 13706 16679
rect 13740 16645 13759 16679
rect 13687 16589 13759 16645
rect 13687 16555 13706 16589
rect 13740 16555 13759 16589
rect 13687 16499 13759 16555
rect 13687 16465 13706 16499
rect 13740 16465 13759 16499
rect 12797 16394 12816 16428
rect 12850 16394 12869 16428
rect 12797 16380 12869 16394
rect 13687 16409 13759 16465
rect 13687 16380 13706 16409
rect 12701 16375 13706 16380
rect 13740 16380 13759 16409
rect 13823 17218 14093 17274
rect 15183 17308 15282 17325
rect 15183 17274 15214 17308
rect 15248 17274 15282 17308
rect 13823 17184 13854 17218
rect 13888 17184 14027 17218
rect 14061 17184 14093 17218
rect 13823 17128 14093 17184
rect 13823 17094 13854 17128
rect 13888 17094 14027 17128
rect 14061 17094 14093 17128
rect 13823 17038 14093 17094
rect 13823 17004 13854 17038
rect 13888 17004 14027 17038
rect 14061 17004 14093 17038
rect 13823 16948 14093 17004
rect 13823 16914 13854 16948
rect 13888 16914 14027 16948
rect 14061 16914 14093 16948
rect 13823 16858 14093 16914
rect 13823 16824 13854 16858
rect 13888 16824 14027 16858
rect 14061 16824 14093 16858
rect 13823 16768 14093 16824
rect 13823 16734 13854 16768
rect 13888 16734 14027 16768
rect 14061 16734 14093 16768
rect 13823 16678 14093 16734
rect 13823 16644 13854 16678
rect 13888 16644 14027 16678
rect 14061 16644 14093 16678
rect 13823 16588 14093 16644
rect 13823 16554 13854 16588
rect 13888 16554 14027 16588
rect 14061 16554 14093 16588
rect 13823 16498 14093 16554
rect 13823 16464 13854 16498
rect 13888 16464 14027 16498
rect 14061 16464 14093 16498
rect 13823 16408 14093 16464
rect 13823 16380 13854 16408
rect 13740 16375 13854 16380
rect 12701 16374 13854 16375
rect 13888 16374 14027 16408
rect 14061 16380 14093 16408
rect 14157 17242 15119 17261
rect 14157 17208 14268 17242
rect 14302 17208 14358 17242
rect 14392 17208 14448 17242
rect 14482 17208 14538 17242
rect 14572 17208 14628 17242
rect 14662 17208 14718 17242
rect 14752 17208 14808 17242
rect 14842 17208 14898 17242
rect 14932 17208 14988 17242
rect 15022 17208 15119 17242
rect 14157 17189 15119 17208
rect 14157 17148 14229 17189
rect 14157 17114 14176 17148
rect 14210 17114 14229 17148
rect 15047 17129 15119 17189
rect 14157 17058 14229 17114
rect 14157 17024 14176 17058
rect 14210 17024 14229 17058
rect 14157 16968 14229 17024
rect 14157 16934 14176 16968
rect 14210 16934 14229 16968
rect 14157 16878 14229 16934
rect 14157 16844 14176 16878
rect 14210 16844 14229 16878
rect 14157 16788 14229 16844
rect 14157 16754 14176 16788
rect 14210 16754 14229 16788
rect 14157 16698 14229 16754
rect 14157 16664 14176 16698
rect 14210 16664 14229 16698
rect 14157 16608 14229 16664
rect 14157 16574 14176 16608
rect 14210 16574 14229 16608
rect 14157 16518 14229 16574
rect 14157 16484 14176 16518
rect 14210 16484 14229 16518
rect 14157 16428 14229 16484
rect 14291 17066 14985 17127
rect 14291 17032 14350 17066
rect 14384 17054 14440 17066
rect 14412 17032 14440 17054
rect 14474 17054 14530 17066
rect 14474 17032 14478 17054
rect 14291 17020 14378 17032
rect 14412 17020 14478 17032
rect 14512 17032 14530 17054
rect 14564 17054 14620 17066
rect 14564 17032 14578 17054
rect 14512 17020 14578 17032
rect 14612 17032 14620 17054
rect 14654 17054 14710 17066
rect 14744 17054 14800 17066
rect 14834 17054 14890 17066
rect 14654 17032 14678 17054
rect 14744 17032 14778 17054
rect 14834 17032 14878 17054
rect 14924 17032 14985 17066
rect 14612 17020 14678 17032
rect 14712 17020 14778 17032
rect 14812 17020 14878 17032
rect 14912 17020 14985 17032
rect 14291 16976 14985 17020
rect 14291 16942 14350 16976
rect 14384 16954 14440 16976
rect 14412 16942 14440 16954
rect 14474 16954 14530 16976
rect 14474 16942 14478 16954
rect 14291 16920 14378 16942
rect 14412 16920 14478 16942
rect 14512 16942 14530 16954
rect 14564 16954 14620 16976
rect 14564 16942 14578 16954
rect 14512 16920 14578 16942
rect 14612 16942 14620 16954
rect 14654 16954 14710 16976
rect 14744 16954 14800 16976
rect 14834 16954 14890 16976
rect 14654 16942 14678 16954
rect 14744 16942 14778 16954
rect 14834 16942 14878 16954
rect 14924 16942 14985 16976
rect 14612 16920 14678 16942
rect 14712 16920 14778 16942
rect 14812 16920 14878 16942
rect 14912 16920 14985 16942
rect 14291 16886 14985 16920
rect 14291 16852 14350 16886
rect 14384 16854 14440 16886
rect 14412 16852 14440 16854
rect 14474 16854 14530 16886
rect 14474 16852 14478 16854
rect 14291 16820 14378 16852
rect 14412 16820 14478 16852
rect 14512 16852 14530 16854
rect 14564 16854 14620 16886
rect 14564 16852 14578 16854
rect 14512 16820 14578 16852
rect 14612 16852 14620 16854
rect 14654 16854 14710 16886
rect 14744 16854 14800 16886
rect 14834 16854 14890 16886
rect 14654 16852 14678 16854
rect 14744 16852 14778 16854
rect 14834 16852 14878 16854
rect 14924 16852 14985 16886
rect 14612 16820 14678 16852
rect 14712 16820 14778 16852
rect 14812 16820 14878 16852
rect 14912 16820 14985 16852
rect 14291 16796 14985 16820
rect 14291 16762 14350 16796
rect 14384 16762 14440 16796
rect 14474 16762 14530 16796
rect 14564 16762 14620 16796
rect 14654 16762 14710 16796
rect 14744 16762 14800 16796
rect 14834 16762 14890 16796
rect 14924 16762 14985 16796
rect 14291 16754 14985 16762
rect 14291 16720 14378 16754
rect 14412 16720 14478 16754
rect 14512 16720 14578 16754
rect 14612 16720 14678 16754
rect 14712 16720 14778 16754
rect 14812 16720 14878 16754
rect 14912 16720 14985 16754
rect 14291 16706 14985 16720
rect 14291 16672 14350 16706
rect 14384 16672 14440 16706
rect 14474 16672 14530 16706
rect 14564 16672 14620 16706
rect 14654 16672 14710 16706
rect 14744 16672 14800 16706
rect 14834 16672 14890 16706
rect 14924 16672 14985 16706
rect 14291 16654 14985 16672
rect 14291 16620 14378 16654
rect 14412 16620 14478 16654
rect 14512 16620 14578 16654
rect 14612 16620 14678 16654
rect 14712 16620 14778 16654
rect 14812 16620 14878 16654
rect 14912 16620 14985 16654
rect 14291 16616 14985 16620
rect 14291 16582 14350 16616
rect 14384 16582 14440 16616
rect 14474 16582 14530 16616
rect 14564 16582 14620 16616
rect 14654 16582 14710 16616
rect 14744 16582 14800 16616
rect 14834 16582 14890 16616
rect 14924 16582 14985 16616
rect 14291 16554 14985 16582
rect 14291 16526 14378 16554
rect 14412 16526 14478 16554
rect 14291 16492 14350 16526
rect 14412 16520 14440 16526
rect 14384 16492 14440 16520
rect 14474 16520 14478 16526
rect 14512 16526 14578 16554
rect 14512 16520 14530 16526
rect 14474 16492 14530 16520
rect 14564 16520 14578 16526
rect 14612 16526 14678 16554
rect 14712 16526 14778 16554
rect 14812 16526 14878 16554
rect 14912 16526 14985 16554
rect 14612 16520 14620 16526
rect 14564 16492 14620 16520
rect 14654 16520 14678 16526
rect 14744 16520 14778 16526
rect 14834 16520 14878 16526
rect 14654 16492 14710 16520
rect 14744 16492 14800 16520
rect 14834 16492 14890 16520
rect 14924 16492 14985 16526
rect 14291 16433 14985 16492
rect 15047 17095 15066 17129
rect 15100 17095 15119 17129
rect 15047 17039 15119 17095
rect 15047 17005 15066 17039
rect 15100 17005 15119 17039
rect 15047 16949 15119 17005
rect 15047 16915 15066 16949
rect 15100 16915 15119 16949
rect 15047 16859 15119 16915
rect 15047 16825 15066 16859
rect 15100 16825 15119 16859
rect 15047 16769 15119 16825
rect 15047 16735 15066 16769
rect 15100 16735 15119 16769
rect 15047 16679 15119 16735
rect 15047 16645 15066 16679
rect 15100 16645 15119 16679
rect 15047 16589 15119 16645
rect 15047 16555 15066 16589
rect 15100 16555 15119 16589
rect 15047 16499 15119 16555
rect 15047 16465 15066 16499
rect 15100 16465 15119 16499
rect 14157 16394 14176 16428
rect 14210 16394 14229 16428
rect 14157 16380 14229 16394
rect 15047 16409 15119 16465
rect 15047 16380 15066 16409
rect 14061 16375 15066 16380
rect 15100 16380 15119 16409
rect 15183 17218 15282 17274
rect 15183 17184 15214 17218
rect 15248 17184 15282 17218
rect 15183 17128 15282 17184
rect 15183 17094 15214 17128
rect 15248 17094 15282 17128
rect 15183 17038 15282 17094
rect 15183 17004 15214 17038
rect 15248 17004 15282 17038
rect 15183 16948 15282 17004
rect 15183 16914 15214 16948
rect 15248 16914 15282 16948
rect 15183 16858 15282 16914
rect 15183 16824 15214 16858
rect 15248 16824 15282 16858
rect 15183 16768 15282 16824
rect 15183 16734 15214 16768
rect 15248 16734 15282 16768
rect 15183 16678 15282 16734
rect 15183 16644 15214 16678
rect 15248 16644 15282 16678
rect 15183 16588 15282 16644
rect 15183 16554 15214 16588
rect 15248 16554 15282 16588
rect 15183 16498 15282 16554
rect 15183 16464 15214 16498
rect 15248 16464 15282 16498
rect 15183 16408 15282 16464
rect 15183 16380 15214 16408
rect 15100 16375 15214 16380
rect 14061 16374 15214 16375
rect 15248 16380 15282 16408
rect 15248 16374 15288 16380
rect 11268 16352 15288 16374
rect 11268 16318 11514 16352
rect 11548 16318 11604 16352
rect 11638 16318 11694 16352
rect 11728 16318 11784 16352
rect 11818 16318 11874 16352
rect 11908 16318 11964 16352
rect 11998 16318 12054 16352
rect 12088 16318 12144 16352
rect 12178 16318 12234 16352
rect 12268 16318 12874 16352
rect 12908 16318 12964 16352
rect 12998 16318 13054 16352
rect 13088 16318 13144 16352
rect 13178 16318 13234 16352
rect 13268 16318 13324 16352
rect 13358 16318 13414 16352
rect 13448 16318 13504 16352
rect 13538 16318 13594 16352
rect 13628 16318 14234 16352
rect 14268 16318 14324 16352
rect 14358 16318 14414 16352
rect 14448 16318 14504 16352
rect 14538 16318 14594 16352
rect 14628 16318 14684 16352
rect 14718 16318 14774 16352
rect 14808 16318 14864 16352
rect 14898 16318 14954 16352
rect 14988 16318 15288 16352
rect 11268 16284 11307 16318
rect 11341 16284 12494 16318
rect 12528 16284 12667 16318
rect 12701 16284 13854 16318
rect 13888 16284 14027 16318
rect 14061 16284 15214 16318
rect 15248 16284 15288 16318
rect 11268 16228 15288 16284
rect 11268 16194 11307 16228
rect 11341 16205 12494 16228
rect 11341 16194 11408 16205
rect 11268 16171 11408 16194
rect 11442 16171 11498 16205
rect 11532 16171 11588 16205
rect 11622 16171 11678 16205
rect 11712 16171 11768 16205
rect 11802 16171 11858 16205
rect 11892 16171 11948 16205
rect 11982 16171 12038 16205
rect 12072 16171 12128 16205
rect 12162 16171 12218 16205
rect 12252 16171 12308 16205
rect 12342 16171 12398 16205
rect 12432 16194 12494 16205
rect 12528 16194 12667 16228
rect 12701 16205 13854 16228
rect 12701 16194 12768 16205
rect 12432 16171 12768 16194
rect 12802 16171 12858 16205
rect 12892 16171 12948 16205
rect 12982 16171 13038 16205
rect 13072 16171 13128 16205
rect 13162 16171 13218 16205
rect 13252 16171 13308 16205
rect 13342 16171 13398 16205
rect 13432 16171 13488 16205
rect 13522 16171 13578 16205
rect 13612 16171 13668 16205
rect 13702 16171 13758 16205
rect 13792 16194 13854 16205
rect 13888 16194 14027 16228
rect 14061 16205 15214 16228
rect 14061 16194 14128 16205
rect 13792 16171 14128 16194
rect 14162 16171 14218 16205
rect 14252 16171 14308 16205
rect 14342 16171 14398 16205
rect 14432 16171 14488 16205
rect 14522 16171 14578 16205
rect 14612 16171 14668 16205
rect 14702 16171 14758 16205
rect 14792 16171 14848 16205
rect 14882 16171 14938 16205
rect 14972 16171 15028 16205
rect 15062 16171 15118 16205
rect 15152 16194 15214 16205
rect 15248 16194 15288 16228
rect 15152 16171 15288 16194
rect 11268 16130 15288 16171
rect 16231 18501 16265 18563
rect 15481 16181 15515 16243
rect 16594 18560 16690 18594
rect 16950 18560 17046 18594
rect 16594 18498 16628 18560
rect 16778 18550 16858 18560
rect 17012 18498 17046 18560
rect 16594 17318 16628 17380
rect 17012 17318 17046 17380
rect 16594 17284 16690 17318
rect 16950 17284 17046 17318
rect 17381 18563 17477 18597
rect 17737 18563 17833 18597
rect 17381 18501 17415 18563
rect 17568 18550 17648 18563
rect 17799 18501 17833 18563
rect 17381 17111 17415 17173
rect 17799 17111 17833 17173
rect 17381 17077 17477 17111
rect 17737 17077 17833 17111
rect 16231 16181 16265 16243
rect 15481 16147 15577 16181
rect 16169 16147 16265 16181
rect 12558 16064 12638 16130
rect 13918 16064 13998 16130
rect 11274 16032 15282 16064
rect 11274 15998 11408 16032
rect 11442 15998 11498 16032
rect 11532 15998 11588 16032
rect 11622 15998 11678 16032
rect 11712 15998 11768 16032
rect 11802 15998 11858 16032
rect 11892 15998 11948 16032
rect 11982 15998 12038 16032
rect 12072 15998 12128 16032
rect 12162 15998 12218 16032
rect 12252 15998 12308 16032
rect 12342 15998 12398 16032
rect 12432 15998 12768 16032
rect 12802 15998 12858 16032
rect 12892 15998 12948 16032
rect 12982 15998 13038 16032
rect 13072 15998 13128 16032
rect 13162 15998 13218 16032
rect 13252 15998 13308 16032
rect 13342 15998 13398 16032
rect 13432 15998 13488 16032
rect 13522 15998 13578 16032
rect 13612 15998 13668 16032
rect 13702 15998 13758 16032
rect 13792 15998 14128 16032
rect 14162 15998 14218 16032
rect 14252 15998 14308 16032
rect 14342 15998 14398 16032
rect 14432 15998 14488 16032
rect 14522 15998 14578 16032
rect 14612 15998 14668 16032
rect 14702 15998 14758 16032
rect 14792 15998 14848 16032
rect 14882 15998 14938 16032
rect 14972 15998 15028 16032
rect 15062 15998 15118 16032
rect 15152 15998 15282 16032
rect 11274 15965 15282 15998
rect 11274 15948 11373 15965
rect 11274 15914 11307 15948
rect 11341 15914 11373 15948
rect 11274 15858 11373 15914
rect 12463 15948 12733 15965
rect 12463 15914 12494 15948
rect 12528 15914 12667 15948
rect 12701 15914 12733 15948
rect 11274 15824 11307 15858
rect 11341 15824 11373 15858
rect 11274 15768 11373 15824
rect 11274 15734 11307 15768
rect 11341 15734 11373 15768
rect 11274 15678 11373 15734
rect 11274 15644 11307 15678
rect 11341 15644 11373 15678
rect 11274 15588 11373 15644
rect 11274 15554 11307 15588
rect 11341 15554 11373 15588
rect 11274 15498 11373 15554
rect 11274 15464 11307 15498
rect 11341 15464 11373 15498
rect 11274 15408 11373 15464
rect 11274 15374 11307 15408
rect 11341 15374 11373 15408
rect 11274 15318 11373 15374
rect 11274 15284 11307 15318
rect 11341 15284 11373 15318
rect 11274 15228 11373 15284
rect 11274 15194 11307 15228
rect 11341 15194 11373 15228
rect 11274 15138 11373 15194
rect 11274 15104 11307 15138
rect 11341 15104 11373 15138
rect 11274 15048 11373 15104
rect 11274 15020 11307 15048
rect 11268 15014 11307 15020
rect 11341 15020 11373 15048
rect 11437 15882 12399 15901
rect 11437 15848 11548 15882
rect 11582 15848 11638 15882
rect 11672 15848 11728 15882
rect 11762 15848 11818 15882
rect 11852 15848 11908 15882
rect 11942 15848 11998 15882
rect 12032 15848 12088 15882
rect 12122 15848 12178 15882
rect 12212 15848 12268 15882
rect 12302 15848 12399 15882
rect 11437 15829 12399 15848
rect 11437 15788 11509 15829
rect 11437 15754 11456 15788
rect 11490 15754 11509 15788
rect 12327 15769 12399 15829
rect 11437 15698 11509 15754
rect 11437 15664 11456 15698
rect 11490 15664 11509 15698
rect 11437 15608 11509 15664
rect 11437 15574 11456 15608
rect 11490 15574 11509 15608
rect 11437 15518 11509 15574
rect 11437 15484 11456 15518
rect 11490 15484 11509 15518
rect 11437 15428 11509 15484
rect 11437 15394 11456 15428
rect 11490 15394 11509 15428
rect 11437 15338 11509 15394
rect 11437 15304 11456 15338
rect 11490 15304 11509 15338
rect 11437 15248 11509 15304
rect 11437 15214 11456 15248
rect 11490 15214 11509 15248
rect 11437 15158 11509 15214
rect 11437 15124 11456 15158
rect 11490 15124 11509 15158
rect 11437 15068 11509 15124
rect 11571 15706 12265 15767
rect 11571 15672 11630 15706
rect 11664 15694 11720 15706
rect 11692 15672 11720 15694
rect 11754 15694 11810 15706
rect 11754 15672 11758 15694
rect 11571 15660 11658 15672
rect 11692 15660 11758 15672
rect 11792 15672 11810 15694
rect 11844 15694 11900 15706
rect 11844 15672 11858 15694
rect 11792 15660 11858 15672
rect 11892 15672 11900 15694
rect 11934 15694 11990 15706
rect 12024 15694 12080 15706
rect 12114 15694 12170 15706
rect 11934 15672 11958 15694
rect 12024 15672 12058 15694
rect 12114 15672 12158 15694
rect 12204 15672 12265 15706
rect 11892 15660 11958 15672
rect 11992 15660 12058 15672
rect 12092 15660 12158 15672
rect 12192 15660 12265 15672
rect 11571 15616 12265 15660
rect 11571 15582 11630 15616
rect 11664 15594 11720 15616
rect 11692 15582 11720 15594
rect 11754 15594 11810 15616
rect 11754 15582 11758 15594
rect 11571 15560 11658 15582
rect 11692 15560 11758 15582
rect 11792 15582 11810 15594
rect 11844 15594 11900 15616
rect 11844 15582 11858 15594
rect 11792 15560 11858 15582
rect 11892 15582 11900 15594
rect 11934 15594 11990 15616
rect 12024 15594 12080 15616
rect 12114 15594 12170 15616
rect 11934 15582 11958 15594
rect 12024 15582 12058 15594
rect 12114 15582 12158 15594
rect 12204 15582 12265 15616
rect 11892 15560 11958 15582
rect 11992 15560 12058 15582
rect 12092 15560 12158 15582
rect 12192 15560 12265 15582
rect 11571 15526 12265 15560
rect 11571 15492 11630 15526
rect 11664 15494 11720 15526
rect 11692 15492 11720 15494
rect 11754 15494 11810 15526
rect 11754 15492 11758 15494
rect 11571 15460 11658 15492
rect 11692 15460 11758 15492
rect 11792 15492 11810 15494
rect 11844 15494 11900 15526
rect 11844 15492 11858 15494
rect 11792 15460 11858 15492
rect 11892 15492 11900 15494
rect 11934 15494 11990 15526
rect 12024 15494 12080 15526
rect 12114 15494 12170 15526
rect 11934 15492 11958 15494
rect 12024 15492 12058 15494
rect 12114 15492 12158 15494
rect 12204 15492 12265 15526
rect 11892 15460 11958 15492
rect 11992 15460 12058 15492
rect 12092 15460 12158 15492
rect 12192 15460 12265 15492
rect 11571 15436 12265 15460
rect 11571 15402 11630 15436
rect 11664 15402 11720 15436
rect 11754 15402 11810 15436
rect 11844 15402 11900 15436
rect 11934 15402 11990 15436
rect 12024 15402 12080 15436
rect 12114 15402 12170 15436
rect 12204 15402 12265 15436
rect 11571 15394 12265 15402
rect 11571 15360 11658 15394
rect 11692 15360 11758 15394
rect 11792 15360 11858 15394
rect 11892 15360 11958 15394
rect 11992 15360 12058 15394
rect 12092 15360 12158 15394
rect 12192 15360 12265 15394
rect 11571 15346 12265 15360
rect 11571 15312 11630 15346
rect 11664 15312 11720 15346
rect 11754 15312 11810 15346
rect 11844 15312 11900 15346
rect 11934 15312 11990 15346
rect 12024 15312 12080 15346
rect 12114 15312 12170 15346
rect 12204 15312 12265 15346
rect 11571 15294 12265 15312
rect 11571 15260 11658 15294
rect 11692 15260 11758 15294
rect 11792 15260 11858 15294
rect 11892 15260 11958 15294
rect 11992 15260 12058 15294
rect 12092 15260 12158 15294
rect 12192 15260 12265 15294
rect 11571 15256 12265 15260
rect 11571 15222 11630 15256
rect 11664 15222 11720 15256
rect 11754 15222 11810 15256
rect 11844 15222 11900 15256
rect 11934 15222 11990 15256
rect 12024 15222 12080 15256
rect 12114 15222 12170 15256
rect 12204 15222 12265 15256
rect 11571 15194 12265 15222
rect 11571 15166 11658 15194
rect 11692 15166 11758 15194
rect 11571 15132 11630 15166
rect 11692 15160 11720 15166
rect 11664 15132 11720 15160
rect 11754 15160 11758 15166
rect 11792 15166 11858 15194
rect 11792 15160 11810 15166
rect 11754 15132 11810 15160
rect 11844 15160 11858 15166
rect 11892 15166 11958 15194
rect 11992 15166 12058 15194
rect 12092 15166 12158 15194
rect 12192 15166 12265 15194
rect 11892 15160 11900 15166
rect 11844 15132 11900 15160
rect 11934 15160 11958 15166
rect 12024 15160 12058 15166
rect 12114 15160 12158 15166
rect 11934 15132 11990 15160
rect 12024 15132 12080 15160
rect 12114 15132 12170 15160
rect 12204 15132 12265 15166
rect 11571 15073 12265 15132
rect 12327 15735 12346 15769
rect 12380 15735 12399 15769
rect 12327 15679 12399 15735
rect 12327 15645 12346 15679
rect 12380 15645 12399 15679
rect 12327 15589 12399 15645
rect 12327 15555 12346 15589
rect 12380 15555 12399 15589
rect 12327 15499 12399 15555
rect 12327 15465 12346 15499
rect 12380 15465 12399 15499
rect 12327 15409 12399 15465
rect 12327 15375 12346 15409
rect 12380 15375 12399 15409
rect 12327 15319 12399 15375
rect 12327 15285 12346 15319
rect 12380 15285 12399 15319
rect 12327 15229 12399 15285
rect 12327 15195 12346 15229
rect 12380 15195 12399 15229
rect 12327 15139 12399 15195
rect 12327 15105 12346 15139
rect 12380 15105 12399 15139
rect 11437 15034 11456 15068
rect 11490 15034 11509 15068
rect 11437 15020 11509 15034
rect 12327 15049 12399 15105
rect 12327 15020 12346 15049
rect 11341 15015 12346 15020
rect 12380 15020 12399 15049
rect 12463 15858 12733 15914
rect 13823 15948 14093 15965
rect 13823 15914 13854 15948
rect 13888 15914 14027 15948
rect 14061 15914 14093 15948
rect 12463 15824 12494 15858
rect 12528 15824 12667 15858
rect 12701 15824 12733 15858
rect 12463 15768 12733 15824
rect 12463 15734 12494 15768
rect 12528 15734 12667 15768
rect 12701 15734 12733 15768
rect 12463 15678 12733 15734
rect 12463 15644 12494 15678
rect 12528 15644 12667 15678
rect 12701 15644 12733 15678
rect 12463 15588 12733 15644
rect 12463 15554 12494 15588
rect 12528 15554 12667 15588
rect 12701 15554 12733 15588
rect 12463 15498 12733 15554
rect 12463 15464 12494 15498
rect 12528 15464 12667 15498
rect 12701 15464 12733 15498
rect 12463 15408 12733 15464
rect 12463 15374 12494 15408
rect 12528 15374 12667 15408
rect 12701 15374 12733 15408
rect 12463 15318 12733 15374
rect 12463 15284 12494 15318
rect 12528 15284 12667 15318
rect 12701 15284 12733 15318
rect 12463 15228 12733 15284
rect 12463 15194 12494 15228
rect 12528 15194 12667 15228
rect 12701 15194 12733 15228
rect 12463 15138 12733 15194
rect 12463 15104 12494 15138
rect 12528 15104 12667 15138
rect 12701 15104 12733 15138
rect 12463 15048 12733 15104
rect 12463 15020 12494 15048
rect 12380 15015 12494 15020
rect 11341 15014 12494 15015
rect 12528 15014 12667 15048
rect 12701 15020 12733 15048
rect 12797 15882 13759 15901
rect 12797 15848 12908 15882
rect 12942 15848 12998 15882
rect 13032 15848 13088 15882
rect 13122 15848 13178 15882
rect 13212 15848 13268 15882
rect 13302 15848 13358 15882
rect 13392 15848 13448 15882
rect 13482 15848 13538 15882
rect 13572 15848 13628 15882
rect 13662 15848 13759 15882
rect 12797 15829 13759 15848
rect 12797 15788 12869 15829
rect 12797 15754 12816 15788
rect 12850 15754 12869 15788
rect 13687 15769 13759 15829
rect 12797 15698 12869 15754
rect 12797 15664 12816 15698
rect 12850 15664 12869 15698
rect 12797 15608 12869 15664
rect 12797 15574 12816 15608
rect 12850 15574 12869 15608
rect 12797 15518 12869 15574
rect 12797 15484 12816 15518
rect 12850 15484 12869 15518
rect 12797 15428 12869 15484
rect 12797 15394 12816 15428
rect 12850 15394 12869 15428
rect 12797 15338 12869 15394
rect 12797 15304 12816 15338
rect 12850 15304 12869 15338
rect 12797 15248 12869 15304
rect 12797 15214 12816 15248
rect 12850 15214 12869 15248
rect 12797 15158 12869 15214
rect 12797 15124 12816 15158
rect 12850 15124 12869 15158
rect 12797 15068 12869 15124
rect 12931 15706 13625 15767
rect 12931 15672 12990 15706
rect 13024 15694 13080 15706
rect 13052 15672 13080 15694
rect 13114 15694 13170 15706
rect 13114 15672 13118 15694
rect 12931 15660 13018 15672
rect 13052 15660 13118 15672
rect 13152 15672 13170 15694
rect 13204 15694 13260 15706
rect 13204 15672 13218 15694
rect 13152 15660 13218 15672
rect 13252 15672 13260 15694
rect 13294 15694 13350 15706
rect 13384 15694 13440 15706
rect 13474 15694 13530 15706
rect 13294 15672 13318 15694
rect 13384 15672 13418 15694
rect 13474 15672 13518 15694
rect 13564 15672 13625 15706
rect 13252 15660 13318 15672
rect 13352 15660 13418 15672
rect 13452 15660 13518 15672
rect 13552 15660 13625 15672
rect 12931 15616 13625 15660
rect 12931 15582 12990 15616
rect 13024 15594 13080 15616
rect 13052 15582 13080 15594
rect 13114 15594 13170 15616
rect 13114 15582 13118 15594
rect 12931 15560 13018 15582
rect 13052 15560 13118 15582
rect 13152 15582 13170 15594
rect 13204 15594 13260 15616
rect 13204 15582 13218 15594
rect 13152 15560 13218 15582
rect 13252 15582 13260 15594
rect 13294 15594 13350 15616
rect 13384 15594 13440 15616
rect 13474 15594 13530 15616
rect 13294 15582 13318 15594
rect 13384 15582 13418 15594
rect 13474 15582 13518 15594
rect 13564 15582 13625 15616
rect 13252 15560 13318 15582
rect 13352 15560 13418 15582
rect 13452 15560 13518 15582
rect 13552 15560 13625 15582
rect 12931 15526 13625 15560
rect 12931 15492 12990 15526
rect 13024 15494 13080 15526
rect 13052 15492 13080 15494
rect 13114 15494 13170 15526
rect 13114 15492 13118 15494
rect 12931 15460 13018 15492
rect 13052 15460 13118 15492
rect 13152 15492 13170 15494
rect 13204 15494 13260 15526
rect 13204 15492 13218 15494
rect 13152 15460 13218 15492
rect 13252 15492 13260 15494
rect 13294 15494 13350 15526
rect 13384 15494 13440 15526
rect 13474 15494 13530 15526
rect 13294 15492 13318 15494
rect 13384 15492 13418 15494
rect 13474 15492 13518 15494
rect 13564 15492 13625 15526
rect 13252 15460 13318 15492
rect 13352 15460 13418 15492
rect 13452 15460 13518 15492
rect 13552 15460 13625 15492
rect 12931 15436 13625 15460
rect 12931 15402 12990 15436
rect 13024 15402 13080 15436
rect 13114 15402 13170 15436
rect 13204 15402 13260 15436
rect 13294 15402 13350 15436
rect 13384 15402 13440 15436
rect 13474 15402 13530 15436
rect 13564 15402 13625 15436
rect 12931 15394 13625 15402
rect 12931 15360 13018 15394
rect 13052 15360 13118 15394
rect 13152 15360 13218 15394
rect 13252 15360 13318 15394
rect 13352 15360 13418 15394
rect 13452 15360 13518 15394
rect 13552 15360 13625 15394
rect 12931 15346 13625 15360
rect 12931 15312 12990 15346
rect 13024 15312 13080 15346
rect 13114 15312 13170 15346
rect 13204 15312 13260 15346
rect 13294 15312 13350 15346
rect 13384 15312 13440 15346
rect 13474 15312 13530 15346
rect 13564 15312 13625 15346
rect 12931 15294 13625 15312
rect 12931 15260 13018 15294
rect 13052 15260 13118 15294
rect 13152 15260 13218 15294
rect 13252 15260 13318 15294
rect 13352 15260 13418 15294
rect 13452 15260 13518 15294
rect 13552 15260 13625 15294
rect 12931 15256 13625 15260
rect 12931 15222 12990 15256
rect 13024 15222 13080 15256
rect 13114 15222 13170 15256
rect 13204 15222 13260 15256
rect 13294 15222 13350 15256
rect 13384 15222 13440 15256
rect 13474 15222 13530 15256
rect 13564 15222 13625 15256
rect 12931 15194 13625 15222
rect 12931 15166 13018 15194
rect 13052 15166 13118 15194
rect 12931 15132 12990 15166
rect 13052 15160 13080 15166
rect 13024 15132 13080 15160
rect 13114 15160 13118 15166
rect 13152 15166 13218 15194
rect 13152 15160 13170 15166
rect 13114 15132 13170 15160
rect 13204 15160 13218 15166
rect 13252 15166 13318 15194
rect 13352 15166 13418 15194
rect 13452 15166 13518 15194
rect 13552 15166 13625 15194
rect 13252 15160 13260 15166
rect 13204 15132 13260 15160
rect 13294 15160 13318 15166
rect 13384 15160 13418 15166
rect 13474 15160 13518 15166
rect 13294 15132 13350 15160
rect 13384 15132 13440 15160
rect 13474 15132 13530 15160
rect 13564 15132 13625 15166
rect 12931 15073 13625 15132
rect 13687 15735 13706 15769
rect 13740 15735 13759 15769
rect 13687 15679 13759 15735
rect 13687 15645 13706 15679
rect 13740 15645 13759 15679
rect 13687 15589 13759 15645
rect 13687 15555 13706 15589
rect 13740 15555 13759 15589
rect 13687 15499 13759 15555
rect 13687 15465 13706 15499
rect 13740 15465 13759 15499
rect 13687 15409 13759 15465
rect 13687 15375 13706 15409
rect 13740 15375 13759 15409
rect 13687 15319 13759 15375
rect 13687 15285 13706 15319
rect 13740 15285 13759 15319
rect 13687 15229 13759 15285
rect 13687 15195 13706 15229
rect 13740 15195 13759 15229
rect 13687 15139 13759 15195
rect 13687 15105 13706 15139
rect 13740 15105 13759 15139
rect 12797 15034 12816 15068
rect 12850 15034 12869 15068
rect 12797 15020 12869 15034
rect 13687 15049 13759 15105
rect 13687 15020 13706 15049
rect 12701 15015 13706 15020
rect 13740 15020 13759 15049
rect 13823 15858 14093 15914
rect 15183 15948 15282 15965
rect 15183 15914 15214 15948
rect 15248 15914 15282 15948
rect 13823 15824 13854 15858
rect 13888 15824 14027 15858
rect 14061 15824 14093 15858
rect 13823 15768 14093 15824
rect 13823 15734 13854 15768
rect 13888 15734 14027 15768
rect 14061 15734 14093 15768
rect 13823 15678 14093 15734
rect 13823 15644 13854 15678
rect 13888 15644 14027 15678
rect 14061 15644 14093 15678
rect 13823 15588 14093 15644
rect 13823 15554 13854 15588
rect 13888 15554 14027 15588
rect 14061 15554 14093 15588
rect 13823 15498 14093 15554
rect 13823 15464 13854 15498
rect 13888 15464 14027 15498
rect 14061 15464 14093 15498
rect 13823 15408 14093 15464
rect 13823 15374 13854 15408
rect 13888 15374 14027 15408
rect 14061 15374 14093 15408
rect 13823 15318 14093 15374
rect 13823 15284 13854 15318
rect 13888 15284 14027 15318
rect 14061 15284 14093 15318
rect 13823 15228 14093 15284
rect 13823 15194 13854 15228
rect 13888 15194 14027 15228
rect 14061 15194 14093 15228
rect 13823 15138 14093 15194
rect 13823 15104 13854 15138
rect 13888 15104 14027 15138
rect 14061 15104 14093 15138
rect 13823 15048 14093 15104
rect 13823 15020 13854 15048
rect 13740 15015 13854 15020
rect 12701 15014 13854 15015
rect 13888 15014 14027 15048
rect 14061 15020 14093 15048
rect 14157 15882 15119 15901
rect 14157 15848 14268 15882
rect 14302 15848 14358 15882
rect 14392 15848 14448 15882
rect 14482 15848 14538 15882
rect 14572 15848 14628 15882
rect 14662 15848 14718 15882
rect 14752 15848 14808 15882
rect 14842 15848 14898 15882
rect 14932 15848 14988 15882
rect 15022 15848 15119 15882
rect 14157 15829 15119 15848
rect 14157 15788 14229 15829
rect 14157 15754 14176 15788
rect 14210 15754 14229 15788
rect 15047 15769 15119 15829
rect 14157 15698 14229 15754
rect 14157 15664 14176 15698
rect 14210 15664 14229 15698
rect 14157 15608 14229 15664
rect 14157 15574 14176 15608
rect 14210 15574 14229 15608
rect 14157 15518 14229 15574
rect 14157 15484 14176 15518
rect 14210 15484 14229 15518
rect 14157 15428 14229 15484
rect 14157 15394 14176 15428
rect 14210 15394 14229 15428
rect 14157 15338 14229 15394
rect 14157 15304 14176 15338
rect 14210 15304 14229 15338
rect 14157 15248 14229 15304
rect 14157 15214 14176 15248
rect 14210 15214 14229 15248
rect 14157 15158 14229 15214
rect 14157 15124 14176 15158
rect 14210 15124 14229 15158
rect 14157 15068 14229 15124
rect 14291 15706 14985 15767
rect 14291 15672 14350 15706
rect 14384 15694 14440 15706
rect 14412 15672 14440 15694
rect 14474 15694 14530 15706
rect 14474 15672 14478 15694
rect 14291 15660 14378 15672
rect 14412 15660 14478 15672
rect 14512 15672 14530 15694
rect 14564 15694 14620 15706
rect 14564 15672 14578 15694
rect 14512 15660 14578 15672
rect 14612 15672 14620 15694
rect 14654 15694 14710 15706
rect 14744 15694 14800 15706
rect 14834 15694 14890 15706
rect 14654 15672 14678 15694
rect 14744 15672 14778 15694
rect 14834 15672 14878 15694
rect 14924 15672 14985 15706
rect 14612 15660 14678 15672
rect 14712 15660 14778 15672
rect 14812 15660 14878 15672
rect 14912 15660 14985 15672
rect 14291 15616 14985 15660
rect 14291 15582 14350 15616
rect 14384 15594 14440 15616
rect 14412 15582 14440 15594
rect 14474 15594 14530 15616
rect 14474 15582 14478 15594
rect 14291 15560 14378 15582
rect 14412 15560 14478 15582
rect 14512 15582 14530 15594
rect 14564 15594 14620 15616
rect 14564 15582 14578 15594
rect 14512 15560 14578 15582
rect 14612 15582 14620 15594
rect 14654 15594 14710 15616
rect 14744 15594 14800 15616
rect 14834 15594 14890 15616
rect 14654 15582 14678 15594
rect 14744 15582 14778 15594
rect 14834 15582 14878 15594
rect 14924 15582 14985 15616
rect 14612 15560 14678 15582
rect 14712 15560 14778 15582
rect 14812 15560 14878 15582
rect 14912 15560 14985 15582
rect 14291 15526 14985 15560
rect 14291 15492 14350 15526
rect 14384 15494 14440 15526
rect 14412 15492 14440 15494
rect 14474 15494 14530 15526
rect 14474 15492 14478 15494
rect 14291 15460 14378 15492
rect 14412 15460 14478 15492
rect 14512 15492 14530 15494
rect 14564 15494 14620 15526
rect 14564 15492 14578 15494
rect 14512 15460 14578 15492
rect 14612 15492 14620 15494
rect 14654 15494 14710 15526
rect 14744 15494 14800 15526
rect 14834 15494 14890 15526
rect 14654 15492 14678 15494
rect 14744 15492 14778 15494
rect 14834 15492 14878 15494
rect 14924 15492 14985 15526
rect 14612 15460 14678 15492
rect 14712 15460 14778 15492
rect 14812 15460 14878 15492
rect 14912 15460 14985 15492
rect 14291 15436 14985 15460
rect 14291 15402 14350 15436
rect 14384 15402 14440 15436
rect 14474 15402 14530 15436
rect 14564 15402 14620 15436
rect 14654 15402 14710 15436
rect 14744 15402 14800 15436
rect 14834 15402 14890 15436
rect 14924 15402 14985 15436
rect 14291 15394 14985 15402
rect 14291 15360 14378 15394
rect 14412 15360 14478 15394
rect 14512 15360 14578 15394
rect 14612 15360 14678 15394
rect 14712 15360 14778 15394
rect 14812 15360 14878 15394
rect 14912 15360 14985 15394
rect 14291 15346 14985 15360
rect 14291 15312 14350 15346
rect 14384 15312 14440 15346
rect 14474 15312 14530 15346
rect 14564 15312 14620 15346
rect 14654 15312 14710 15346
rect 14744 15312 14800 15346
rect 14834 15312 14890 15346
rect 14924 15312 14985 15346
rect 14291 15294 14985 15312
rect 14291 15260 14378 15294
rect 14412 15260 14478 15294
rect 14512 15260 14578 15294
rect 14612 15260 14678 15294
rect 14712 15260 14778 15294
rect 14812 15260 14878 15294
rect 14912 15260 14985 15294
rect 14291 15256 14985 15260
rect 14291 15222 14350 15256
rect 14384 15222 14440 15256
rect 14474 15222 14530 15256
rect 14564 15222 14620 15256
rect 14654 15222 14710 15256
rect 14744 15222 14800 15256
rect 14834 15222 14890 15256
rect 14924 15222 14985 15256
rect 14291 15194 14985 15222
rect 14291 15166 14378 15194
rect 14412 15166 14478 15194
rect 14291 15132 14350 15166
rect 14412 15160 14440 15166
rect 14384 15132 14440 15160
rect 14474 15160 14478 15166
rect 14512 15166 14578 15194
rect 14512 15160 14530 15166
rect 14474 15132 14530 15160
rect 14564 15160 14578 15166
rect 14612 15166 14678 15194
rect 14712 15166 14778 15194
rect 14812 15166 14878 15194
rect 14912 15166 14985 15194
rect 14612 15160 14620 15166
rect 14564 15132 14620 15160
rect 14654 15160 14678 15166
rect 14744 15160 14778 15166
rect 14834 15160 14878 15166
rect 14654 15132 14710 15160
rect 14744 15132 14800 15160
rect 14834 15132 14890 15160
rect 14924 15132 14985 15166
rect 14291 15073 14985 15132
rect 15047 15735 15066 15769
rect 15100 15735 15119 15769
rect 15047 15679 15119 15735
rect 15047 15645 15066 15679
rect 15100 15645 15119 15679
rect 15047 15589 15119 15645
rect 15047 15555 15066 15589
rect 15100 15555 15119 15589
rect 15047 15499 15119 15555
rect 15047 15465 15066 15499
rect 15100 15465 15119 15499
rect 15047 15409 15119 15465
rect 15047 15375 15066 15409
rect 15100 15375 15119 15409
rect 15047 15319 15119 15375
rect 15047 15285 15066 15319
rect 15100 15285 15119 15319
rect 15047 15229 15119 15285
rect 15047 15195 15066 15229
rect 15100 15195 15119 15229
rect 15047 15139 15119 15195
rect 15047 15105 15066 15139
rect 15100 15105 15119 15139
rect 14157 15034 14176 15068
rect 14210 15034 14229 15068
rect 14157 15020 14229 15034
rect 15047 15049 15119 15105
rect 15047 15020 15066 15049
rect 14061 15015 15066 15020
rect 15100 15020 15119 15049
rect 15183 15858 15282 15914
rect 15183 15824 15214 15858
rect 15248 15824 15282 15858
rect 15183 15768 15282 15824
rect 15183 15734 15214 15768
rect 15248 15734 15282 15768
rect 15183 15678 15282 15734
rect 15183 15644 15214 15678
rect 15248 15644 15282 15678
rect 15183 15588 15282 15644
rect 15183 15554 15214 15588
rect 15248 15554 15282 15588
rect 15183 15498 15282 15554
rect 15183 15464 15214 15498
rect 15248 15464 15282 15498
rect 15183 15408 15282 15464
rect 15183 15374 15214 15408
rect 15248 15374 15282 15408
rect 15183 15318 15282 15374
rect 15183 15284 15214 15318
rect 15248 15284 15282 15318
rect 15183 15228 15282 15284
rect 15183 15194 15214 15228
rect 15248 15194 15282 15228
rect 15183 15138 15282 15194
rect 15183 15104 15214 15138
rect 15248 15104 15282 15138
rect 15183 15048 15282 15104
rect 15183 15020 15214 15048
rect 15100 15015 15214 15020
rect 14061 15014 15214 15015
rect 15248 15020 15282 15048
rect 15248 15014 15288 15020
rect 11268 14992 15288 15014
rect 11268 14958 11514 14992
rect 11548 14958 11604 14992
rect 11638 14958 11694 14992
rect 11728 14958 11784 14992
rect 11818 14958 11874 14992
rect 11908 14958 11964 14992
rect 11998 14958 12054 14992
rect 12088 14958 12144 14992
rect 12178 14958 12234 14992
rect 12268 14958 12874 14992
rect 12908 14958 12964 14992
rect 12998 14958 13054 14992
rect 13088 14958 13144 14992
rect 13178 14958 13234 14992
rect 13268 14958 13324 14992
rect 13358 14958 13414 14992
rect 13448 14958 13504 14992
rect 13538 14958 13594 14992
rect 13628 14958 14234 14992
rect 14268 14958 14324 14992
rect 14358 14958 14414 14992
rect 14448 14958 14504 14992
rect 14538 14958 14594 14992
rect 14628 14958 14684 14992
rect 14718 14958 14774 14992
rect 14808 14958 14864 14992
rect 14898 14958 14954 14992
rect 14988 14958 15288 14992
rect 11268 14924 11307 14958
rect 11341 14924 12494 14958
rect 12528 14924 12667 14958
rect 12701 14924 13854 14958
rect 13888 14924 14027 14958
rect 14061 14924 15214 14958
rect 15248 14924 15288 14958
rect 11268 14868 15288 14924
rect 11268 14834 11307 14868
rect 11341 14845 12494 14868
rect 11341 14834 11408 14845
rect 11268 14811 11408 14834
rect 11442 14811 11498 14845
rect 11532 14811 11588 14845
rect 11622 14811 11678 14845
rect 11712 14811 11768 14845
rect 11802 14811 11858 14845
rect 11892 14811 11948 14845
rect 11982 14811 12038 14845
rect 12072 14811 12128 14845
rect 12162 14811 12218 14845
rect 12252 14811 12308 14845
rect 12342 14811 12398 14845
rect 12432 14834 12494 14845
rect 12528 14834 12667 14868
rect 12701 14845 13854 14868
rect 12701 14834 12768 14845
rect 12432 14811 12768 14834
rect 12802 14811 12858 14845
rect 12892 14811 12948 14845
rect 12982 14811 13038 14845
rect 13072 14811 13128 14845
rect 13162 14811 13218 14845
rect 13252 14811 13308 14845
rect 13342 14811 13398 14845
rect 13432 14811 13488 14845
rect 13522 14811 13578 14845
rect 13612 14811 13668 14845
rect 13702 14811 13758 14845
rect 13792 14834 13854 14845
rect 13888 14834 14027 14868
rect 14061 14845 15214 14868
rect 14061 14834 14128 14845
rect 13792 14811 14128 14834
rect 14162 14811 14218 14845
rect 14252 14811 14308 14845
rect 14342 14811 14398 14845
rect 14432 14811 14488 14845
rect 14522 14811 14578 14845
rect 14612 14811 14668 14845
rect 14702 14811 14758 14845
rect 14792 14811 14848 14845
rect 14882 14811 14938 14845
rect 14972 14811 15028 14845
rect 15062 14811 15118 14845
rect 15152 14834 15214 14845
rect 15248 14834 15288 14868
rect 15152 14811 15288 14834
rect 11268 14770 15288 14811
rect 12540 14600 12630 14610
rect 12540 14550 12560 14600
rect 12610 14550 12630 14600
rect 12540 14540 12630 14550
rect 13938 14600 14028 14610
rect 13938 14550 13958 14600
rect 14008 14550 14028 14600
rect 13938 14540 14028 14550
rect 11168 14250 11228 14270
rect 11168 14220 11178 14250
rect 11078 14210 11178 14220
rect 11218 14210 11228 14250
rect 11078 14200 11228 14210
rect 11078 14160 11098 14200
rect 11138 14160 11228 14200
rect 11078 14150 11228 14160
rect 11078 14140 11178 14150
rect 11168 14110 11178 14140
rect 11218 14110 11228 14150
rect 11168 14090 11228 14110
rect 13248 14250 13308 14270
rect 13248 14210 13258 14250
rect 13298 14210 13308 14250
rect 13248 14150 13308 14210
rect 13248 14110 13258 14150
rect 13298 14110 13308 14150
rect 13248 14090 13308 14110
rect 15328 14260 15468 14270
rect 15328 14250 15548 14260
rect 15328 14210 15338 14250
rect 15378 14210 15418 14250
rect 15458 14240 15548 14250
rect 15458 14210 15488 14240
rect 15328 14200 15488 14210
rect 15528 14200 15548 14240
rect 15328 14160 15548 14200
rect 15328 14150 15488 14160
rect 15328 14110 15338 14150
rect 15378 14110 15418 14150
rect 15458 14120 15488 14150
rect 15528 14120 15548 14160
rect 15458 14110 15548 14120
rect 15328 14100 15548 14110
rect 15328 14090 15468 14100
rect 11178 14050 11218 14090
rect 13258 14050 13298 14090
rect 11158 14030 11238 14050
rect 11158 13990 11178 14030
rect 11218 13990 11238 14030
rect 11158 13970 11238 13990
rect 11318 14030 11398 14050
rect 11318 13990 11338 14030
rect 11378 13990 11398 14030
rect 11318 13970 11398 13990
rect 11478 14030 11558 14050
rect 11478 13990 11498 14030
rect 11538 13990 11558 14030
rect 11478 13970 11558 13990
rect 11638 14030 11718 14050
rect 11638 13990 11658 14030
rect 11698 13990 11718 14030
rect 11638 13970 11718 13990
rect 11798 14030 11878 14050
rect 11798 13990 11818 14030
rect 11858 13990 11878 14030
rect 11798 13970 11878 13990
rect 11958 14030 12038 14050
rect 11958 13990 11978 14030
rect 12018 13990 12038 14030
rect 11958 13970 12038 13990
rect 12118 14030 12198 14050
rect 12118 13990 12138 14030
rect 12178 13990 12198 14030
rect 12118 13970 12198 13990
rect 12278 14030 12358 14050
rect 12278 13990 12298 14030
rect 12338 13990 12358 14030
rect 12278 13970 12358 13990
rect 12438 14030 12518 14050
rect 12438 13990 12458 14030
rect 12498 13990 12518 14030
rect 12438 13970 12518 13990
rect 12598 14030 12678 14050
rect 12598 13990 12618 14030
rect 12658 13990 12678 14030
rect 12598 13970 12678 13990
rect 12758 14030 12838 14050
rect 12758 13990 12778 14030
rect 12818 13990 12838 14030
rect 12758 13970 12838 13990
rect 12918 14030 12998 14050
rect 12918 13990 12938 14030
rect 12978 13990 12998 14030
rect 12918 13970 12998 13990
rect 13078 14030 13158 14050
rect 13078 13990 13098 14030
rect 13138 13990 13158 14030
rect 13078 13970 13158 13990
rect 13238 14030 13318 14050
rect 13238 13990 13258 14030
rect 13298 13990 13318 14030
rect 13238 13970 13318 13990
rect 13398 14030 13478 14050
rect 13398 13990 13418 14030
rect 13458 13990 13478 14030
rect 13398 13970 13478 13990
rect 13558 14030 13638 14050
rect 13558 13990 13578 14030
rect 13618 13990 13638 14030
rect 13558 13970 13638 13990
rect 13718 14030 13798 14050
rect 13718 13990 13738 14030
rect 13778 13990 13798 14030
rect 13718 13970 13798 13990
rect 13878 14030 13958 14050
rect 13878 13990 13898 14030
rect 13938 13990 13958 14030
rect 13878 13970 13958 13990
rect 14038 14030 14118 14050
rect 14038 13990 14058 14030
rect 14098 13990 14118 14030
rect 14038 13970 14118 13990
rect 14198 14030 14278 14050
rect 14198 13990 14218 14030
rect 14258 13990 14278 14030
rect 14198 13970 14278 13990
rect 14358 14030 14438 14050
rect 14358 13990 14378 14030
rect 14418 13990 14438 14030
rect 14358 13970 14438 13990
rect 14518 14030 14598 14050
rect 14518 13990 14538 14030
rect 14578 13990 14598 14030
rect 14518 13970 14598 13990
rect 14678 14030 14758 14050
rect 14678 13990 14698 14030
rect 14738 13990 14758 14030
rect 14678 13970 14758 13990
rect 14838 14030 14918 14050
rect 14838 13990 14858 14030
rect 14898 13990 14918 14030
rect 14838 13970 14918 13990
rect 14998 14030 15078 14050
rect 14998 13990 15018 14030
rect 15058 13990 15078 14030
rect 14998 13970 15078 13990
rect 15158 14030 15238 14050
rect 15158 13990 15178 14030
rect 15218 13990 15238 14030
rect 15158 13970 15238 13990
rect 11898 13760 11978 13780
rect 11898 13720 11918 13760
rect 11958 13720 11978 13760
rect 11898 13700 11978 13720
rect 14578 13760 14658 13780
rect 14578 13720 14598 13760
rect 14638 13720 14658 13760
rect 14578 13700 14658 13720
rect 11918 13660 11958 13700
rect 14598 13660 14638 13700
rect 10748 13640 10808 13660
rect 10748 13600 10758 13640
rect 10798 13600 10808 13640
rect 10748 13540 10808 13600
rect 10748 13500 10758 13540
rect 10798 13500 10808 13540
rect 10748 13440 10808 13500
rect 10748 13400 10758 13440
rect 10798 13400 10808 13440
rect 10748 13340 10808 13400
rect 10748 13300 10758 13340
rect 10798 13300 10808 13340
rect 10748 13240 10808 13300
rect 10748 13200 10758 13240
rect 10798 13200 10808 13240
rect 10748 13180 10808 13200
rect 11828 13640 12048 13660
rect 11828 13600 11838 13640
rect 11878 13600 11918 13640
rect 11958 13600 11998 13640
rect 12038 13600 12048 13640
rect 11828 13540 12048 13600
rect 11828 13500 11838 13540
rect 11878 13500 11918 13540
rect 11958 13500 11998 13540
rect 12038 13500 12048 13540
rect 11828 13440 12048 13500
rect 11828 13400 11838 13440
rect 11878 13400 11918 13440
rect 11958 13400 11998 13440
rect 12038 13400 12048 13440
rect 11828 13340 12048 13400
rect 11828 13300 11838 13340
rect 11878 13300 11918 13340
rect 11958 13300 11998 13340
rect 12038 13300 12048 13340
rect 11828 13240 12048 13300
rect 11828 13200 11838 13240
rect 11878 13200 11918 13240
rect 11958 13200 11998 13240
rect 12038 13200 12048 13240
rect 11828 13180 12048 13200
rect 13068 13640 13128 13660
rect 13068 13600 13078 13640
rect 13118 13600 13128 13640
rect 13068 13540 13128 13600
rect 13068 13500 13078 13540
rect 13118 13500 13128 13540
rect 13068 13440 13128 13500
rect 13068 13400 13078 13440
rect 13118 13400 13128 13440
rect 13068 13340 13128 13400
rect 13068 13300 13078 13340
rect 13118 13300 13128 13340
rect 13068 13240 13128 13300
rect 13068 13200 13078 13240
rect 13118 13200 13128 13240
rect 10738 13160 10818 13180
rect 10738 13120 10758 13160
rect 10798 13120 10818 13160
rect 13068 13150 13128 13200
rect 10738 13100 10818 13120
rect 10918 13120 10998 13140
rect 10918 13080 10938 13120
rect 10978 13080 10998 13120
rect 10918 13060 10998 13080
rect 11158 13120 11238 13140
rect 11158 13080 11178 13120
rect 11218 13080 11238 13120
rect 11158 13060 11238 13080
rect 11398 13120 11478 13140
rect 11398 13080 11418 13120
rect 11458 13080 11478 13120
rect 11398 13060 11478 13080
rect 11638 13120 11718 13140
rect 11638 13080 11658 13120
rect 11698 13080 11718 13120
rect 11638 13060 11718 13080
rect 12278 13120 12358 13140
rect 12278 13080 12298 13120
rect 12338 13080 12358 13120
rect 12278 13060 12358 13080
rect 12518 13120 12598 13140
rect 12518 13080 12538 13120
rect 12578 13080 12598 13120
rect 12518 13060 12598 13080
rect 12758 13120 12838 13140
rect 12758 13080 12778 13120
rect 12818 13080 12838 13120
rect 13068 13110 13078 13150
rect 13118 13110 13128 13150
rect 13068 13090 13128 13110
rect 13428 13640 13488 13660
rect 13428 13600 13438 13640
rect 13478 13600 13488 13640
rect 13428 13540 13488 13600
rect 13428 13500 13438 13540
rect 13478 13500 13488 13540
rect 13428 13440 13488 13500
rect 13428 13400 13438 13440
rect 13478 13400 13488 13440
rect 13428 13340 13488 13400
rect 13428 13300 13438 13340
rect 13478 13300 13488 13340
rect 13428 13240 13488 13300
rect 13428 13200 13438 13240
rect 13478 13200 13488 13240
rect 13428 13150 13488 13200
rect 14508 13640 14728 13660
rect 14508 13600 14518 13640
rect 14558 13600 14598 13640
rect 14638 13600 14678 13640
rect 14718 13600 14728 13640
rect 14508 13540 14728 13600
rect 14508 13500 14518 13540
rect 14558 13500 14598 13540
rect 14638 13500 14678 13540
rect 14718 13500 14728 13540
rect 14508 13440 14728 13500
rect 14508 13400 14518 13440
rect 14558 13400 14598 13440
rect 14638 13400 14678 13440
rect 14718 13400 14728 13440
rect 14508 13340 14728 13400
rect 14508 13300 14518 13340
rect 14558 13300 14598 13340
rect 14638 13300 14678 13340
rect 14718 13300 14728 13340
rect 14508 13240 14728 13300
rect 14508 13200 14518 13240
rect 14558 13200 14598 13240
rect 14638 13200 14678 13240
rect 14718 13200 14728 13240
rect 14508 13180 14728 13200
rect 15748 13640 15808 13660
rect 15748 13600 15758 13640
rect 15798 13600 15808 13640
rect 15748 13540 15808 13600
rect 15748 13500 15758 13540
rect 15798 13500 15808 13540
rect 15748 13440 15808 13500
rect 15748 13400 15758 13440
rect 15798 13400 15808 13440
rect 23208 13510 23308 13530
rect 23208 13450 23228 13510
rect 23288 13450 23308 13510
rect 23208 13430 23308 13450
rect 15748 13340 15808 13400
rect 15748 13300 15758 13340
rect 15798 13300 15808 13340
rect 15748 13240 15808 13300
rect 15748 13200 15758 13240
rect 15798 13200 15808 13240
rect 15748 13180 15808 13200
rect 23031 13253 23127 13287
rect 23387 13253 23483 13287
rect 23031 13191 23065 13253
rect 13428 13110 13438 13150
rect 13478 13110 13488 13150
rect 23008 13170 23031 13190
rect 23449 13191 23483 13253
rect 23065 13170 23088 13190
rect 13428 13090 13488 13110
rect 13718 13120 13798 13140
rect 12758 13060 12838 13080
rect 13718 13080 13738 13120
rect 13778 13080 13798 13120
rect 13718 13060 13798 13080
rect 13958 13120 14038 13140
rect 13958 13080 13978 13120
rect 14018 13080 14038 13120
rect 13958 13060 14038 13080
rect 14198 13120 14278 13140
rect 14198 13080 14218 13120
rect 14258 13080 14278 13120
rect 14198 13060 14278 13080
rect 14838 13120 14918 13140
rect 14838 13080 14858 13120
rect 14898 13080 14918 13120
rect 14838 13060 14918 13080
rect 15078 13120 15158 13140
rect 15078 13080 15098 13120
rect 15138 13080 15158 13120
rect 15078 13060 15158 13080
rect 15318 13120 15398 13140
rect 15318 13080 15338 13120
rect 15378 13080 15398 13120
rect 15318 13060 15398 13080
rect 15558 13120 15638 13140
rect 15558 13080 15578 13120
rect 15618 13080 15638 13120
rect 23008 13130 23028 13170
rect 23068 13130 23088 13170
rect 23008 13110 23031 13130
rect 15558 13060 15638 13080
rect 20318 12780 20398 12800
rect 11429 12742 11487 12760
rect 11429 12708 11441 12742
rect 11475 12708 11487 12742
rect 11429 12690 11487 12708
rect 11789 12742 11847 12760
rect 11789 12708 11801 12742
rect 11835 12708 11847 12742
rect 11789 12690 11847 12708
rect 11909 12742 11967 12760
rect 11909 12708 11921 12742
rect 11955 12708 11967 12742
rect 11909 12690 11967 12708
rect 12269 12742 12327 12760
rect 12269 12708 12281 12742
rect 12315 12708 12327 12742
rect 12269 12690 12327 12708
rect 12389 12742 12447 12760
rect 12389 12708 12401 12742
rect 12435 12708 12447 12742
rect 14109 12742 14167 12760
rect 12389 12690 12447 12708
rect 12798 12720 12878 12740
rect 12798 12680 12818 12720
rect 12858 12680 12878 12720
rect 11368 12630 11428 12650
rect 11368 12590 11378 12630
rect 11418 12590 11428 12630
rect 11368 12570 11428 12590
rect 11488 12630 11548 12650
rect 11488 12590 11498 12630
rect 11538 12590 11548 12630
rect 11488 12570 11548 12590
rect 11608 12630 11668 12650
rect 11608 12590 11618 12630
rect 11658 12590 11668 12630
rect 11608 12570 11668 12590
rect 11728 12630 11788 12650
rect 11728 12590 11738 12630
rect 11778 12590 11788 12630
rect 11728 12570 11788 12590
rect 11848 12630 11908 12650
rect 11848 12590 11858 12630
rect 11898 12590 11908 12630
rect 11848 12570 11908 12590
rect 11968 12630 12028 12650
rect 11968 12590 11978 12630
rect 12018 12590 12028 12630
rect 11968 12570 12028 12590
rect 12088 12630 12148 12650
rect 12088 12590 12098 12630
rect 12138 12590 12148 12630
rect 12088 12570 12148 12590
rect 12208 12630 12268 12650
rect 12208 12590 12218 12630
rect 12258 12590 12268 12630
rect 12208 12570 12268 12590
rect 12328 12630 12388 12650
rect 12328 12590 12338 12630
rect 12378 12590 12388 12630
rect 12328 12570 12388 12590
rect 12448 12630 12508 12650
rect 12448 12590 12458 12630
rect 12498 12590 12508 12630
rect 12448 12570 12508 12590
rect 12568 12630 12628 12650
rect 12568 12590 12578 12630
rect 12618 12590 12628 12630
rect 12568 12570 12628 12590
rect 12798 12640 12878 12680
rect 12798 12600 12818 12640
rect 12858 12600 12878 12640
rect 12798 12560 12878 12600
rect 11530 12512 11588 12530
rect 11530 12478 11542 12512
rect 11576 12478 11588 12512
rect 11530 12460 11588 12478
rect 11688 12512 11746 12530
rect 11688 12478 11700 12512
rect 11734 12478 11746 12512
rect 11688 12460 11746 12478
rect 12012 12512 12070 12530
rect 12012 12478 12024 12512
rect 12058 12478 12070 12512
rect 12012 12460 12070 12478
rect 12166 12512 12224 12530
rect 12166 12478 12178 12512
rect 12212 12478 12224 12512
rect 12166 12460 12224 12478
rect 12490 12512 12548 12530
rect 12490 12478 12502 12512
rect 12536 12478 12548 12512
rect 12798 12520 12818 12560
rect 12858 12520 12878 12560
rect 12798 12500 12878 12520
rect 13678 12720 13758 12740
rect 13678 12680 13698 12720
rect 13738 12680 13758 12720
rect 14109 12708 14121 12742
rect 14155 12708 14167 12742
rect 14109 12690 14167 12708
rect 14229 12742 14287 12760
rect 14229 12708 14241 12742
rect 14275 12708 14287 12742
rect 14229 12690 14287 12708
rect 14589 12742 14647 12760
rect 14589 12708 14601 12742
rect 14635 12708 14647 12742
rect 14589 12690 14647 12708
rect 14709 12742 14767 12760
rect 14709 12708 14721 12742
rect 14755 12708 14767 12742
rect 14709 12690 14767 12708
rect 15069 12742 15127 12760
rect 15069 12708 15081 12742
rect 15115 12708 15127 12742
rect 20318 12740 20338 12780
rect 20378 12740 20398 12780
rect 20318 12720 20398 12740
rect 20718 12780 20798 12800
rect 20718 12740 20738 12780
rect 20778 12740 20798 12780
rect 20718 12720 20798 12740
rect 15069 12690 15127 12708
rect 13678 12640 13758 12680
rect 19418 12660 19598 12680
rect 13678 12600 13698 12640
rect 13738 12600 13758 12640
rect 13678 12560 13758 12600
rect 13928 12630 13988 12650
rect 13928 12590 13938 12630
rect 13978 12590 13988 12630
rect 13928 12570 13988 12590
rect 14048 12630 14108 12650
rect 14048 12590 14058 12630
rect 14098 12590 14108 12630
rect 14048 12570 14108 12590
rect 14168 12630 14228 12650
rect 14168 12590 14178 12630
rect 14218 12590 14228 12630
rect 14168 12570 14228 12590
rect 14288 12630 14348 12650
rect 14288 12590 14298 12630
rect 14338 12590 14348 12630
rect 14288 12570 14348 12590
rect 14408 12630 14468 12650
rect 14408 12590 14418 12630
rect 14458 12590 14468 12630
rect 14408 12570 14468 12590
rect 14528 12630 14588 12650
rect 14528 12590 14538 12630
rect 14578 12590 14588 12630
rect 14528 12570 14588 12590
rect 14648 12630 14708 12650
rect 14648 12590 14658 12630
rect 14698 12590 14708 12630
rect 14648 12570 14708 12590
rect 14768 12630 14828 12650
rect 14768 12590 14778 12630
rect 14818 12590 14828 12630
rect 14768 12570 14828 12590
rect 14888 12630 14948 12650
rect 14888 12590 14898 12630
rect 14938 12590 14948 12630
rect 14888 12570 14948 12590
rect 15008 12630 15068 12650
rect 15008 12590 15018 12630
rect 15058 12590 15068 12630
rect 15008 12570 15068 12590
rect 15128 12630 15188 12650
rect 15128 12590 15138 12630
rect 15178 12590 15188 12630
rect 15128 12570 15188 12590
rect 19418 12620 19438 12660
rect 19478 12620 19538 12660
rect 19578 12620 19598 12660
rect 13678 12520 13698 12560
rect 13738 12520 13758 12560
rect 19418 12560 19598 12620
rect 13678 12500 13758 12520
rect 14008 12512 14066 12530
rect 12490 12460 12548 12478
rect 14008 12478 14020 12512
rect 14054 12478 14066 12512
rect 14008 12460 14066 12478
rect 14332 12512 14390 12530
rect 14332 12478 14344 12512
rect 14378 12478 14390 12512
rect 14332 12460 14390 12478
rect 14486 12512 14544 12530
rect 14486 12478 14498 12512
rect 14532 12478 14544 12512
rect 14486 12460 14544 12478
rect 14810 12512 14868 12530
rect 14810 12478 14822 12512
rect 14856 12478 14868 12512
rect 14810 12460 14868 12478
rect 14968 12512 15026 12530
rect 14968 12478 14980 12512
rect 15014 12478 15026 12512
rect 14968 12460 15026 12478
rect 19418 12520 19438 12560
rect 19478 12520 19538 12560
rect 19578 12520 19598 12560
rect 19418 12460 19598 12520
rect 19418 12420 19438 12460
rect 19478 12420 19538 12460
rect 19578 12420 19598 12460
rect 19418 12360 19598 12420
rect 19418 12320 19438 12360
rect 19478 12320 19538 12360
rect 19578 12320 19598 12360
rect 19418 12260 19598 12320
rect 19418 12220 19438 12260
rect 19478 12220 19538 12260
rect 19578 12220 19598 12260
rect 19418 12200 19598 12220
rect 19718 12660 19798 12680
rect 19718 12620 19738 12660
rect 19778 12620 19798 12660
rect 19718 12560 19798 12620
rect 19718 12520 19738 12560
rect 19778 12520 19798 12560
rect 19718 12460 19798 12520
rect 19718 12420 19738 12460
rect 19778 12420 19798 12460
rect 19718 12360 19798 12420
rect 19718 12320 19738 12360
rect 19778 12320 19798 12360
rect 19718 12260 19798 12320
rect 19718 12220 19738 12260
rect 19778 12220 19798 12260
rect 19718 12200 19798 12220
rect 19918 12660 19998 12680
rect 19918 12620 19938 12660
rect 19978 12620 19998 12660
rect 19918 12560 19998 12620
rect 19918 12520 19938 12560
rect 19978 12520 19998 12560
rect 19918 12460 19998 12520
rect 19918 12420 19938 12460
rect 19978 12420 19998 12460
rect 19918 12360 19998 12420
rect 19918 12320 19938 12360
rect 19978 12320 19998 12360
rect 19918 12260 19998 12320
rect 19918 12220 19938 12260
rect 19978 12220 19998 12260
rect 19918 12200 19998 12220
rect 20118 12660 20198 12680
rect 20118 12620 20138 12660
rect 20178 12620 20198 12660
rect 20118 12560 20198 12620
rect 20118 12520 20138 12560
rect 20178 12520 20198 12560
rect 20118 12460 20198 12520
rect 20118 12420 20138 12460
rect 20178 12420 20198 12460
rect 20118 12360 20198 12420
rect 20118 12320 20138 12360
rect 20178 12320 20198 12360
rect 20118 12260 20198 12320
rect 20118 12220 20138 12260
rect 20178 12220 20198 12260
rect 20118 12200 20198 12220
rect 20318 12660 20398 12680
rect 20318 12620 20338 12660
rect 20378 12620 20398 12660
rect 20318 12560 20398 12620
rect 20318 12520 20338 12560
rect 20378 12520 20398 12560
rect 20318 12460 20398 12520
rect 20318 12420 20338 12460
rect 20378 12420 20398 12460
rect 20318 12360 20398 12420
rect 20318 12320 20338 12360
rect 20378 12320 20398 12360
rect 20318 12260 20398 12320
rect 20318 12220 20338 12260
rect 20378 12220 20398 12260
rect 20318 12200 20398 12220
rect 20518 12660 20598 12680
rect 20518 12620 20538 12660
rect 20578 12620 20598 12660
rect 20518 12560 20598 12620
rect 20518 12520 20538 12560
rect 20578 12520 20598 12560
rect 20518 12460 20598 12520
rect 20518 12420 20538 12460
rect 20578 12420 20598 12460
rect 20518 12360 20598 12420
rect 20518 12320 20538 12360
rect 20578 12320 20598 12360
rect 20518 12260 20598 12320
rect 20518 12220 20538 12260
rect 20578 12220 20598 12260
rect 20518 12200 20598 12220
rect 20718 12660 20798 12680
rect 20718 12620 20738 12660
rect 20778 12620 20798 12660
rect 20718 12560 20798 12620
rect 20718 12520 20738 12560
rect 20778 12520 20798 12560
rect 20718 12460 20798 12520
rect 20718 12420 20738 12460
rect 20778 12420 20798 12460
rect 20718 12360 20798 12420
rect 20718 12320 20738 12360
rect 20778 12320 20798 12360
rect 20718 12260 20798 12320
rect 20718 12220 20738 12260
rect 20778 12220 20798 12260
rect 20718 12200 20798 12220
rect 20918 12660 20998 12680
rect 20918 12620 20938 12660
rect 20978 12620 20998 12660
rect 20918 12560 20998 12620
rect 20918 12520 20938 12560
rect 20978 12520 20998 12560
rect 20918 12460 20998 12520
rect 20918 12420 20938 12460
rect 20978 12420 20998 12460
rect 20918 12360 20998 12420
rect 20918 12320 20938 12360
rect 20978 12320 20998 12360
rect 20918 12260 20998 12320
rect 20918 12220 20938 12260
rect 20978 12220 20998 12260
rect 20918 12200 20998 12220
rect 21118 12660 21198 12680
rect 21118 12620 21138 12660
rect 21178 12620 21198 12660
rect 21118 12560 21198 12620
rect 21118 12520 21138 12560
rect 21178 12520 21198 12560
rect 21118 12460 21198 12520
rect 21118 12420 21138 12460
rect 21178 12420 21198 12460
rect 21118 12360 21198 12420
rect 21118 12320 21138 12360
rect 21178 12320 21198 12360
rect 21118 12260 21198 12320
rect 21118 12220 21138 12260
rect 21178 12220 21198 12260
rect 21118 12200 21198 12220
rect 21318 12660 21398 12680
rect 21318 12620 21338 12660
rect 21378 12620 21398 12660
rect 21318 12560 21398 12620
rect 21318 12520 21338 12560
rect 21378 12520 21398 12560
rect 21318 12460 21398 12520
rect 21318 12420 21338 12460
rect 21378 12420 21398 12460
rect 21318 12360 21398 12420
rect 21318 12320 21338 12360
rect 21378 12320 21398 12360
rect 21318 12260 21398 12320
rect 21318 12220 21338 12260
rect 21378 12220 21398 12260
rect 21318 12200 21398 12220
rect 21518 12660 21698 12680
rect 21518 12620 21538 12660
rect 21578 12620 21638 12660
rect 21678 12620 21698 12660
rect 21518 12560 21698 12620
rect 21518 12520 21538 12560
rect 21578 12520 21638 12560
rect 21678 12520 21698 12560
rect 21518 12460 21698 12520
rect 21518 12420 21538 12460
rect 21578 12420 21638 12460
rect 21678 12420 21698 12460
rect 21518 12360 21698 12420
rect 21518 12320 21538 12360
rect 21578 12320 21638 12360
rect 21678 12320 21698 12360
rect 21518 12260 21698 12320
rect 21518 12220 21538 12260
rect 21578 12220 21638 12260
rect 21678 12220 21698 12260
rect 21518 12200 21698 12220
rect 19518 12140 19598 12200
rect 19518 12100 19538 12140
rect 19578 12100 19598 12140
rect 19518 12080 19598 12100
rect 21518 12140 21598 12160
rect 21518 12100 21538 12140
rect 21578 12100 21598 12140
rect 21518 12080 21598 12100
rect 23065 13110 23088 13130
rect 20998 11980 21078 12000
rect 20998 11940 21018 11980
rect 21058 11940 21078 11980
rect 10708 11920 10768 11940
rect 10708 11880 10718 11920
rect 10758 11880 10768 11920
rect 10708 11860 10768 11880
rect 10878 11910 10958 11930
rect 10878 11870 10898 11910
rect 10938 11870 10958 11910
rect 10878 11850 10958 11870
rect 11368 11910 11428 11930
rect 11368 11870 11378 11910
rect 11418 11870 11428 11910
rect 11368 11850 11428 11870
rect 11598 11910 11678 11930
rect 11598 11870 11618 11910
rect 11658 11870 11678 11910
rect 11598 11850 11678 11870
rect 12088 11910 12148 11930
rect 12088 11870 12098 11910
rect 12138 11870 12148 11910
rect 12088 11850 12148 11870
rect 12318 11910 12398 11930
rect 12318 11870 12338 11910
rect 12378 11870 12398 11910
rect 12318 11850 12398 11870
rect 12748 11910 12808 11930
rect 12748 11870 12758 11910
rect 12798 11870 12808 11910
rect 12748 11850 12808 11870
rect 13748 11910 13808 11930
rect 13748 11870 13758 11910
rect 13798 11870 13808 11910
rect 13748 11850 13808 11870
rect 14158 11910 14238 11930
rect 14158 11870 14178 11910
rect 14218 11870 14238 11910
rect 14158 11850 14238 11870
rect 14408 11910 14468 11930
rect 14408 11870 14418 11910
rect 14458 11870 14468 11910
rect 14408 11850 14468 11870
rect 14878 11910 14958 11930
rect 14878 11870 14898 11910
rect 14938 11870 14958 11910
rect 14878 11850 14958 11870
rect 15128 11910 15188 11930
rect 15128 11870 15138 11910
rect 15178 11870 15188 11910
rect 15128 11850 15188 11870
rect 15598 11910 15678 11930
rect 15598 11870 15618 11910
rect 15658 11870 15678 11910
rect 15598 11850 15678 11870
rect 15788 11920 15848 11940
rect 15788 11880 15798 11920
rect 15838 11880 15848 11920
rect 20998 11920 21078 11940
rect 22118 11980 22198 12000
rect 22118 11940 22138 11980
rect 22178 11940 22198 11980
rect 23031 11983 23065 12045
rect 23449 11983 23483 12045
rect 23031 11949 23127 11983
rect 23387 11949 23483 11983
rect 22118 11920 22198 11940
rect 15788 11860 15848 11880
rect 19918 11870 19998 11890
rect 19508 11830 19588 11850
rect 19508 11810 19528 11830
rect 10448 11790 10588 11810
rect 10448 11750 10458 11790
rect 10498 11750 10538 11790
rect 10578 11750 10588 11790
rect 10448 11690 10588 11750
rect 10448 11650 10458 11690
rect 10498 11650 10538 11690
rect 10578 11650 10588 11690
rect 10448 11630 10588 11650
rect 10648 11790 10708 11810
rect 10648 11750 10658 11790
rect 10698 11750 10708 11790
rect 10648 11690 10708 11750
rect 10648 11650 10658 11690
rect 10698 11650 10708 11690
rect 10648 11630 10708 11650
rect 10768 11790 10828 11810
rect 10768 11750 10778 11790
rect 10818 11750 10828 11790
rect 10768 11690 10828 11750
rect 10768 11650 10778 11690
rect 10818 11650 10828 11690
rect 10768 11630 10828 11650
rect 10888 11790 10948 11810
rect 10888 11750 10898 11790
rect 10938 11750 10948 11790
rect 10888 11690 10948 11750
rect 10888 11650 10898 11690
rect 10938 11650 10948 11690
rect 10888 11630 10948 11650
rect 11008 11790 11068 11810
rect 11008 11750 11018 11790
rect 11058 11750 11068 11790
rect 11008 11690 11068 11750
rect 11008 11650 11018 11690
rect 11058 11650 11068 11690
rect 11008 11630 11068 11650
rect 11128 11790 11188 11810
rect 11128 11750 11138 11790
rect 11178 11750 11188 11790
rect 11128 11690 11188 11750
rect 11128 11650 11138 11690
rect 11178 11650 11188 11690
rect 11128 11630 11188 11650
rect 11248 11790 11308 11810
rect 11248 11750 11258 11790
rect 11298 11750 11308 11790
rect 11248 11690 11308 11750
rect 11248 11650 11258 11690
rect 11298 11650 11308 11690
rect 11248 11630 11308 11650
rect 11368 11790 11428 11810
rect 11368 11750 11378 11790
rect 11418 11750 11428 11790
rect 11368 11690 11428 11750
rect 11368 11650 11378 11690
rect 11418 11650 11428 11690
rect 11368 11630 11428 11650
rect 11488 11790 11548 11810
rect 11488 11750 11498 11790
rect 11538 11750 11548 11790
rect 11488 11690 11548 11750
rect 11488 11650 11498 11690
rect 11538 11650 11548 11690
rect 11488 11630 11548 11650
rect 11608 11790 11668 11810
rect 11608 11750 11618 11790
rect 11658 11750 11668 11790
rect 11608 11690 11668 11750
rect 11608 11650 11618 11690
rect 11658 11650 11668 11690
rect 11608 11630 11668 11650
rect 11728 11790 11788 11810
rect 11728 11750 11738 11790
rect 11778 11750 11788 11790
rect 11728 11690 11788 11750
rect 11728 11650 11738 11690
rect 11778 11650 11788 11690
rect 11728 11630 11788 11650
rect 11848 11790 11908 11810
rect 11848 11750 11858 11790
rect 11898 11750 11908 11790
rect 11848 11690 11908 11750
rect 11848 11650 11858 11690
rect 11898 11650 11908 11690
rect 11848 11630 11908 11650
rect 11968 11790 12028 11810
rect 11968 11750 11978 11790
rect 12018 11750 12028 11790
rect 11968 11690 12028 11750
rect 11968 11650 11978 11690
rect 12018 11650 12028 11690
rect 11968 11630 12028 11650
rect 12088 11790 12148 11810
rect 12088 11750 12098 11790
rect 12138 11750 12148 11790
rect 12088 11690 12148 11750
rect 12088 11650 12098 11690
rect 12138 11650 12148 11690
rect 12088 11630 12148 11650
rect 12208 11790 12268 11810
rect 12208 11750 12218 11790
rect 12258 11750 12268 11790
rect 12208 11690 12268 11750
rect 12208 11650 12218 11690
rect 12258 11650 12268 11690
rect 12208 11630 12268 11650
rect 12328 11790 12388 11810
rect 12328 11750 12338 11790
rect 12378 11750 12388 11790
rect 12328 11690 12388 11750
rect 12328 11650 12338 11690
rect 12378 11650 12388 11690
rect 12328 11630 12388 11650
rect 12448 11790 12508 11810
rect 12448 11750 12458 11790
rect 12498 11750 12508 11790
rect 12448 11690 12508 11750
rect 12448 11650 12458 11690
rect 12498 11650 12508 11690
rect 12448 11630 12508 11650
rect 12568 11790 12628 11810
rect 12568 11750 12578 11790
rect 12618 11750 12628 11790
rect 12568 11690 12628 11750
rect 12568 11650 12578 11690
rect 12618 11650 12628 11690
rect 12568 11630 12628 11650
rect 12688 11790 12748 11810
rect 12688 11750 12698 11790
rect 12738 11750 12748 11790
rect 12688 11690 12748 11750
rect 12688 11650 12698 11690
rect 12738 11650 12748 11690
rect 12688 11630 12748 11650
rect 12808 11790 12868 11810
rect 12808 11750 12818 11790
rect 12858 11750 12868 11790
rect 12808 11690 12868 11750
rect 12808 11650 12818 11690
rect 12858 11650 12868 11690
rect 12808 11630 12868 11650
rect 12928 11790 13068 11810
rect 12928 11750 12938 11790
rect 12978 11750 13018 11790
rect 13058 11750 13068 11790
rect 12928 11690 13068 11750
rect 12928 11650 12938 11690
rect 12978 11650 13018 11690
rect 13058 11650 13068 11690
rect 12928 11630 13068 11650
rect 13488 11790 13628 11810
rect 13488 11750 13498 11790
rect 13538 11750 13578 11790
rect 13618 11750 13628 11790
rect 13488 11690 13628 11750
rect 13488 11650 13498 11690
rect 13538 11650 13578 11690
rect 13618 11650 13628 11690
rect 13488 11630 13628 11650
rect 13688 11790 13748 11810
rect 13688 11750 13698 11790
rect 13738 11750 13748 11790
rect 13688 11690 13748 11750
rect 13688 11650 13698 11690
rect 13738 11650 13748 11690
rect 13688 11630 13748 11650
rect 13808 11790 13868 11810
rect 13808 11750 13818 11790
rect 13858 11750 13868 11790
rect 13808 11690 13868 11750
rect 13808 11650 13818 11690
rect 13858 11650 13868 11690
rect 13808 11630 13868 11650
rect 13928 11790 13988 11810
rect 13928 11750 13938 11790
rect 13978 11750 13988 11790
rect 13928 11690 13988 11750
rect 13928 11650 13938 11690
rect 13978 11650 13988 11690
rect 13928 11630 13988 11650
rect 14048 11790 14108 11810
rect 14048 11750 14058 11790
rect 14098 11750 14108 11790
rect 14048 11690 14108 11750
rect 14048 11650 14058 11690
rect 14098 11650 14108 11690
rect 14048 11630 14108 11650
rect 14168 11790 14228 11810
rect 14168 11750 14178 11790
rect 14218 11750 14228 11790
rect 14168 11690 14228 11750
rect 14168 11650 14178 11690
rect 14218 11650 14228 11690
rect 14168 11630 14228 11650
rect 14288 11790 14348 11810
rect 14288 11750 14298 11790
rect 14338 11750 14348 11790
rect 14288 11690 14348 11750
rect 14288 11650 14298 11690
rect 14338 11650 14348 11690
rect 14288 11630 14348 11650
rect 14408 11790 14468 11810
rect 14408 11750 14418 11790
rect 14458 11750 14468 11790
rect 14408 11690 14468 11750
rect 14408 11650 14418 11690
rect 14458 11650 14468 11690
rect 14408 11630 14468 11650
rect 14528 11790 14588 11810
rect 14528 11750 14538 11790
rect 14578 11750 14588 11790
rect 14528 11690 14588 11750
rect 14528 11650 14538 11690
rect 14578 11650 14588 11690
rect 14528 11630 14588 11650
rect 14648 11790 14708 11810
rect 14648 11750 14658 11790
rect 14698 11750 14708 11790
rect 14648 11690 14708 11750
rect 14648 11650 14658 11690
rect 14698 11650 14708 11690
rect 14648 11630 14708 11650
rect 14768 11790 14828 11810
rect 14768 11750 14778 11790
rect 14818 11750 14828 11790
rect 14768 11690 14828 11750
rect 14768 11650 14778 11690
rect 14818 11650 14828 11690
rect 14768 11630 14828 11650
rect 14888 11790 14948 11810
rect 14888 11750 14898 11790
rect 14938 11750 14948 11790
rect 14888 11690 14948 11750
rect 14888 11650 14898 11690
rect 14938 11650 14948 11690
rect 14888 11630 14948 11650
rect 15008 11790 15068 11810
rect 15008 11750 15018 11790
rect 15058 11750 15068 11790
rect 15008 11690 15068 11750
rect 15008 11650 15018 11690
rect 15058 11650 15068 11690
rect 15008 11630 15068 11650
rect 15128 11790 15188 11810
rect 15128 11750 15138 11790
rect 15178 11750 15188 11790
rect 15128 11690 15188 11750
rect 15128 11650 15138 11690
rect 15178 11650 15188 11690
rect 15128 11630 15188 11650
rect 15248 11790 15308 11810
rect 15248 11750 15258 11790
rect 15298 11750 15308 11790
rect 15248 11690 15308 11750
rect 15248 11650 15258 11690
rect 15298 11650 15308 11690
rect 15248 11630 15308 11650
rect 15368 11790 15428 11810
rect 15368 11750 15378 11790
rect 15418 11750 15428 11790
rect 15368 11690 15428 11750
rect 15368 11650 15378 11690
rect 15418 11650 15428 11690
rect 15368 11630 15428 11650
rect 15488 11790 15548 11810
rect 15488 11750 15498 11790
rect 15538 11750 15548 11790
rect 15488 11690 15548 11750
rect 15488 11650 15498 11690
rect 15538 11650 15548 11690
rect 15488 11630 15548 11650
rect 15608 11790 15668 11810
rect 15608 11750 15618 11790
rect 15658 11750 15668 11790
rect 15608 11690 15668 11750
rect 15608 11650 15618 11690
rect 15658 11650 15668 11690
rect 15608 11630 15668 11650
rect 15728 11790 15788 11810
rect 15728 11750 15738 11790
rect 15778 11750 15788 11790
rect 15728 11690 15788 11750
rect 15728 11650 15738 11690
rect 15778 11650 15788 11690
rect 15728 11630 15788 11650
rect 15848 11790 15908 11810
rect 15848 11750 15858 11790
rect 15898 11750 15908 11790
rect 15848 11690 15908 11750
rect 15848 11650 15858 11690
rect 15898 11650 15908 11690
rect 15848 11630 15908 11650
rect 15968 11790 16108 11810
rect 15968 11750 15978 11790
rect 16018 11750 16058 11790
rect 16098 11750 16108 11790
rect 15968 11690 16108 11750
rect 19468 11790 19528 11810
rect 19568 11810 19588 11830
rect 19918 11830 19938 11870
rect 19978 11830 19998 11870
rect 19918 11810 19998 11830
rect 20168 11830 20248 11850
rect 20168 11810 20188 11830
rect 19568 11790 20188 11810
rect 20228 11810 20248 11830
rect 20648 11830 20728 11850
rect 20648 11810 20668 11830
rect 20228 11790 20288 11810
rect 19468 11770 20288 11790
rect 19468 11730 19508 11770
rect 19598 11730 19638 11770
rect 19858 11730 19898 11770
rect 20118 11730 20158 11770
rect 20248 11730 20288 11770
rect 20608 11790 20668 11810
rect 20708 11810 20728 11830
rect 20998 11810 21038 11920
rect 21308 11830 21388 11850
rect 21308 11810 21328 11830
rect 20708 11790 21328 11810
rect 21368 11810 21388 11830
rect 21788 11830 21868 11850
rect 21788 11810 21808 11830
rect 21368 11790 21428 11810
rect 20608 11770 21428 11790
rect 20608 11730 20648 11770
rect 20738 11730 20778 11770
rect 20998 11730 21038 11770
rect 21258 11730 21298 11770
rect 21388 11730 21428 11770
rect 21748 11790 21808 11810
rect 21848 11810 21868 11830
rect 22138 11810 22178 11920
rect 22448 11830 22528 11850
rect 22448 11810 22468 11830
rect 21848 11790 22468 11810
rect 22508 11810 22528 11830
rect 22508 11790 22568 11810
rect 21748 11770 22568 11790
rect 21748 11730 21788 11770
rect 21878 11730 21918 11770
rect 22138 11730 22178 11770
rect 22398 11730 22438 11770
rect 22528 11730 22568 11770
rect 15968 11650 15978 11690
rect 16018 11650 16058 11690
rect 16098 11650 16108 11690
rect 15968 11630 16108 11650
rect 19448 11710 19528 11730
rect 19448 11670 19468 11710
rect 19508 11670 19528 11710
rect 19448 11610 19528 11670
rect 10528 11570 10588 11590
rect 10528 11530 10538 11570
rect 10578 11530 10588 11570
rect 10528 11510 10588 11530
rect 12928 11570 12988 11590
rect 12928 11530 12938 11570
rect 12978 11530 12988 11570
rect 12928 11510 12988 11530
rect 13568 11570 13628 11590
rect 13568 11530 13578 11570
rect 13618 11530 13628 11570
rect 13568 11510 13628 11530
rect 15968 11570 16028 11590
rect 15968 11530 15978 11570
rect 16018 11530 16028 11570
rect 19448 11570 19468 11610
rect 19508 11570 19528 11610
rect 19448 11550 19528 11570
rect 19578 11710 19658 11730
rect 19578 11670 19598 11710
rect 19638 11670 19658 11710
rect 19578 11610 19658 11670
rect 19578 11570 19598 11610
rect 19638 11570 19658 11610
rect 19578 11550 19658 11570
rect 19708 11710 19788 11730
rect 19708 11670 19728 11710
rect 19768 11670 19788 11710
rect 19708 11610 19788 11670
rect 19708 11570 19728 11610
rect 19768 11570 19788 11610
rect 19708 11550 19788 11570
rect 19838 11710 19918 11730
rect 19838 11670 19858 11710
rect 19898 11670 19918 11710
rect 19838 11610 19918 11670
rect 19838 11570 19858 11610
rect 19898 11570 19918 11610
rect 19838 11550 19918 11570
rect 19968 11710 20048 11730
rect 19968 11670 19988 11710
rect 20028 11670 20048 11710
rect 19968 11610 20048 11670
rect 19968 11570 19988 11610
rect 20028 11570 20048 11610
rect 19968 11550 20048 11570
rect 20098 11710 20188 11730
rect 20098 11670 20118 11710
rect 20158 11670 20188 11710
rect 20098 11610 20188 11670
rect 20098 11570 20118 11610
rect 20158 11570 20188 11610
rect 20098 11550 20188 11570
rect 20228 11710 20308 11730
rect 20228 11670 20248 11710
rect 20288 11670 20308 11710
rect 20228 11610 20308 11670
rect 20228 11570 20248 11610
rect 20288 11570 20308 11610
rect 20228 11550 20308 11570
rect 20488 11710 20668 11730
rect 20488 11670 20508 11710
rect 20548 11670 20608 11710
rect 20648 11670 20668 11710
rect 20488 11610 20668 11670
rect 20488 11570 20508 11610
rect 20548 11570 20608 11610
rect 20648 11570 20668 11610
rect 20488 11550 20668 11570
rect 20718 11710 20798 11730
rect 20718 11670 20738 11710
rect 20778 11670 20798 11710
rect 20718 11610 20798 11670
rect 20718 11570 20738 11610
rect 20778 11570 20798 11610
rect 20718 11550 20798 11570
rect 20848 11710 20928 11730
rect 20848 11670 20868 11710
rect 20908 11670 20928 11710
rect 20848 11610 20928 11670
rect 20848 11570 20868 11610
rect 20908 11570 20928 11610
rect 20848 11550 20928 11570
rect 20978 11710 21058 11730
rect 20978 11670 20998 11710
rect 21038 11670 21058 11710
rect 20978 11610 21058 11670
rect 20978 11570 20998 11610
rect 21038 11570 21058 11610
rect 20978 11550 21058 11570
rect 21108 11710 21188 11730
rect 21108 11670 21128 11710
rect 21168 11670 21188 11710
rect 21108 11610 21188 11670
rect 21108 11570 21128 11610
rect 21168 11570 21188 11610
rect 21108 11550 21188 11570
rect 21238 11710 21318 11730
rect 21238 11670 21258 11710
rect 21298 11670 21318 11710
rect 21238 11610 21318 11670
rect 21238 11570 21258 11610
rect 21298 11570 21318 11610
rect 21238 11550 21318 11570
rect 21368 11710 21548 11730
rect 21368 11670 21388 11710
rect 21428 11670 21488 11710
rect 21528 11670 21548 11710
rect 21368 11610 21548 11670
rect 21368 11570 21388 11610
rect 21428 11570 21488 11610
rect 21528 11570 21548 11610
rect 21368 11550 21548 11570
rect 21628 11710 21808 11730
rect 21628 11670 21648 11710
rect 21688 11670 21748 11710
rect 21788 11670 21808 11710
rect 21628 11610 21808 11670
rect 21628 11570 21648 11610
rect 21688 11570 21748 11610
rect 21788 11570 21808 11610
rect 21628 11550 21808 11570
rect 21858 11710 21938 11730
rect 21858 11670 21878 11710
rect 21918 11670 21938 11710
rect 21858 11610 21938 11670
rect 21858 11570 21878 11610
rect 21918 11570 21938 11610
rect 21858 11550 21938 11570
rect 21988 11710 22068 11730
rect 21988 11670 22008 11710
rect 22048 11670 22068 11710
rect 21988 11610 22068 11670
rect 21988 11570 22008 11610
rect 22048 11570 22068 11610
rect 21988 11550 22068 11570
rect 22118 11710 22198 11730
rect 22118 11670 22138 11710
rect 22178 11670 22198 11710
rect 22118 11610 22198 11670
rect 22118 11570 22138 11610
rect 22178 11570 22198 11610
rect 22118 11550 22198 11570
rect 22248 11710 22328 11730
rect 22248 11670 22268 11710
rect 22308 11670 22328 11710
rect 22248 11610 22328 11670
rect 22248 11570 22268 11610
rect 22308 11570 22328 11610
rect 22248 11550 22328 11570
rect 22378 11710 22458 11730
rect 22378 11670 22398 11710
rect 22438 11670 22458 11710
rect 22378 11610 22458 11670
rect 22378 11570 22398 11610
rect 22438 11570 22458 11610
rect 22378 11550 22458 11570
rect 22508 11710 22688 11730
rect 22508 11670 22528 11710
rect 22568 11670 22628 11710
rect 22668 11670 22688 11710
rect 22508 11610 22688 11670
rect 22508 11570 22528 11610
rect 22568 11570 22628 11610
rect 22668 11570 22688 11610
rect 22508 11550 22688 11570
rect 23438 11580 23548 11600
rect 15968 11510 16028 11530
rect 19618 11490 19698 11510
rect 19618 11450 19638 11490
rect 19678 11450 19698 11490
rect 19618 11430 19698 11450
rect 20058 11490 20138 11510
rect 20058 11450 20078 11490
rect 20118 11450 20138 11490
rect 20058 11430 20138 11450
rect 20848 11480 20928 11500
rect 20848 11440 20868 11480
rect 20908 11440 20928 11480
rect 20848 11420 20928 11440
rect 21898 11490 21978 11510
rect 21898 11450 21918 11490
rect 21958 11450 21978 11490
rect 21898 11430 21978 11450
rect 22028 11390 22068 11550
rect 22248 11390 22288 11550
rect 23438 11510 23458 11580
rect 23528 11510 23548 11580
rect 22738 11490 22818 11510
rect 22738 11450 22758 11490
rect 22798 11450 22818 11490
rect 22738 11430 22818 11450
rect 23438 11490 23548 11510
rect 23438 11390 23478 11490
rect 22028 11350 23648 11390
rect 23608 11340 23648 11350
rect 23608 11320 23688 11340
rect 21898 11270 21978 11290
rect 21898 11230 21918 11270
rect 21958 11230 21978 11270
rect 23608 11280 23628 11320
rect 23668 11280 23688 11320
rect 23608 11260 23688 11280
rect 23608 11250 23648 11260
rect 21898 11210 21978 11230
rect 22028 11210 23648 11250
rect 19708 11150 19788 11170
rect 19708 11110 19728 11150
rect 19768 11110 19788 11150
rect 19708 11090 19788 11110
rect 20758 11150 20838 11170
rect 20758 11110 20778 11150
rect 20818 11110 20838 11150
rect 20758 11090 20838 11110
rect 21198 11150 21278 11170
rect 21198 11110 21218 11150
rect 21258 11110 21278 11150
rect 21198 11090 21278 11110
rect 22028 11050 22068 11210
rect 22248 11050 22288 11210
rect 22738 11150 22818 11170
rect 22738 11110 22758 11150
rect 22798 11110 22818 11150
rect 22738 11090 22818 11110
rect 23438 11090 23478 11210
rect 23438 11070 23548 11090
rect 19348 11030 19528 11050
rect 19348 10990 19368 11030
rect 19408 10990 19468 11030
rect 19508 10990 19528 11030
rect 19348 10970 19528 10990
rect 19578 11030 19658 11050
rect 19578 10990 19598 11030
rect 19638 10990 19658 11030
rect 19578 10970 19658 10990
rect 19708 11030 19788 11050
rect 19708 10990 19728 11030
rect 19768 10990 19788 11030
rect 19708 10970 19788 10990
rect 19838 11030 19918 11050
rect 19838 10990 19858 11030
rect 19898 10990 19918 11030
rect 19838 10970 19918 10990
rect 19968 11030 20048 11050
rect 19968 10990 19988 11030
rect 20028 10990 20048 11030
rect 19968 10970 20048 10990
rect 20098 11030 20178 11050
rect 20098 10990 20118 11030
rect 20158 10990 20178 11030
rect 20098 10970 20178 10990
rect 20228 11030 20408 11050
rect 20228 10990 20248 11030
rect 20288 10990 20348 11030
rect 20388 10990 20408 11030
rect 20228 10970 20408 10990
rect 20588 11030 20668 11050
rect 20588 10990 20608 11030
rect 20648 10990 20668 11030
rect 20588 10970 20668 10990
rect 20718 11030 20798 11050
rect 20718 10990 20738 11030
rect 20778 10990 20798 11030
rect 20718 10970 20798 10990
rect 20848 11030 20928 11050
rect 20848 10990 20868 11030
rect 20908 10990 20928 11030
rect 20848 10970 20928 10990
rect 20978 11030 21058 11050
rect 20978 10990 20998 11030
rect 21038 10990 21058 11030
rect 20978 10970 21058 10990
rect 21108 11030 21188 11050
rect 21108 10990 21128 11030
rect 21168 10990 21188 11030
rect 21108 10970 21188 10990
rect 21238 11030 21318 11050
rect 21238 10990 21258 11030
rect 21298 10990 21318 11030
rect 21238 10970 21318 10990
rect 21368 11030 21448 11050
rect 21368 10990 21388 11030
rect 21428 10990 21448 11030
rect 21368 10970 21448 10990
rect 21628 11030 21808 11050
rect 21628 10990 21648 11030
rect 21688 10990 21748 11030
rect 21788 10990 21808 11030
rect 21628 10970 21808 10990
rect 21858 11030 21938 11050
rect 21858 10990 21878 11030
rect 21918 10990 21938 11030
rect 21858 10970 21938 10990
rect 21988 11030 22068 11050
rect 21988 10990 22008 11030
rect 22048 10990 22068 11030
rect 21988 10970 22068 10990
rect 22118 11030 22198 11050
rect 22118 10990 22138 11030
rect 22178 10990 22198 11030
rect 22118 10970 22198 10990
rect 22248 11030 22328 11050
rect 22248 10990 22268 11030
rect 22308 10990 22328 11030
rect 22248 10970 22328 10990
rect 22378 11030 22458 11050
rect 22378 10990 22398 11030
rect 22438 10990 22458 11030
rect 22378 10970 22458 10990
rect 22508 11030 22688 11050
rect 22508 10990 22528 11030
rect 22568 10990 22628 11030
rect 22668 10990 22688 11030
rect 22508 10970 22688 10990
rect 23438 11000 23458 11070
rect 23528 11000 23548 11070
rect 23438 10980 23548 11000
rect 19468 10930 19508 10970
rect 19598 10930 19638 10970
rect 19858 10930 19898 10970
rect 20118 10930 20158 10970
rect 20248 10930 20288 10970
rect 19468 10910 20288 10930
rect 19468 10890 19528 10910
rect 19508 10860 19528 10890
rect 19578 10890 20178 10910
rect 19578 10860 19598 10890
rect 19508 10840 19598 10860
rect 19858 10780 19898 10890
rect 20158 10860 20178 10890
rect 20228 10890 20288 10910
rect 20608 10930 20648 10970
rect 20738 10930 20778 10970
rect 20998 10930 21038 10970
rect 21258 10930 21298 10970
rect 21388 10930 21428 10970
rect 20608 10910 21428 10930
rect 20608 10890 20668 10910
rect 20228 10860 20248 10890
rect 20158 10840 20248 10860
rect 20648 10870 20668 10890
rect 20708 10890 21328 10910
rect 20708 10870 20728 10890
rect 20648 10850 20728 10870
rect 20978 10870 21058 10890
rect 20978 10830 20998 10870
rect 21038 10830 21058 10870
rect 21308 10870 21328 10890
rect 21368 10890 21428 10910
rect 21748 10930 21788 10970
rect 21878 10930 21918 10970
rect 22138 10930 22178 10970
rect 22398 10930 22438 10970
rect 22528 10930 22568 10970
rect 21748 10910 22568 10930
rect 21368 10870 21388 10890
rect 21748 10880 21808 10910
rect 21308 10850 21388 10870
rect 21788 10870 21808 10880
rect 21848 10880 22468 10910
rect 21848 10870 21868 10880
rect 21788 10850 21868 10870
rect 20978 10810 21058 10830
rect 22138 10780 22178 10880
rect 22448 10870 22468 10880
rect 22508 10880 22568 10910
rect 22508 10870 22528 10880
rect 22448 10850 22528 10870
rect 11898 10750 11968 10770
rect 11898 10710 11908 10750
rect 11948 10710 11968 10750
rect 11898 10690 11968 10710
rect 12068 10750 12148 10770
rect 12068 10710 12088 10750
rect 12128 10710 12148 10750
rect 12068 10690 12148 10710
rect 12248 10750 12328 10770
rect 12248 10710 12268 10750
rect 12308 10710 12328 10750
rect 12248 10690 12328 10710
rect 12428 10750 12508 10770
rect 12428 10710 12448 10750
rect 12488 10710 12508 10750
rect 12428 10690 12508 10710
rect 12608 10750 12688 10770
rect 12608 10710 12628 10750
rect 12668 10710 12688 10750
rect 12608 10690 12688 10710
rect 12788 10750 12868 10770
rect 12788 10710 12808 10750
rect 12848 10710 12868 10750
rect 12788 10690 12868 10710
rect 12968 10750 13048 10770
rect 12968 10710 12988 10750
rect 13028 10710 13048 10750
rect 12968 10690 13048 10710
rect 13148 10750 13218 10770
rect 13148 10710 13168 10750
rect 13208 10710 13218 10750
rect 13148 10690 13218 10710
rect 13338 10750 13408 10770
rect 13338 10710 13348 10750
rect 13388 10710 13408 10750
rect 13338 10690 13408 10710
rect 13508 10750 13588 10770
rect 13508 10710 13528 10750
rect 13568 10710 13588 10750
rect 13508 10690 13588 10710
rect 13688 10750 13768 10770
rect 13688 10710 13708 10750
rect 13748 10710 13768 10750
rect 13688 10690 13768 10710
rect 13868 10750 13948 10770
rect 13868 10710 13888 10750
rect 13928 10710 13948 10750
rect 13868 10690 13948 10710
rect 14048 10750 14128 10770
rect 14048 10710 14068 10750
rect 14108 10710 14128 10750
rect 14048 10690 14128 10710
rect 14228 10750 14308 10770
rect 14228 10710 14248 10750
rect 14288 10710 14308 10750
rect 14228 10690 14308 10710
rect 14408 10750 14488 10770
rect 14408 10710 14428 10750
rect 14468 10710 14488 10750
rect 14408 10690 14488 10710
rect 14588 10750 14658 10770
rect 14588 10710 14608 10750
rect 14648 10710 14658 10750
rect 14588 10690 14658 10710
rect 19838 10760 19918 10780
rect 19838 10720 19858 10760
rect 19898 10720 19918 10760
rect 19838 10700 19918 10720
rect 22118 10760 22198 10780
rect 22118 10720 22138 10760
rect 22178 10720 22198 10760
rect 22118 10700 22198 10720
rect 23031 10733 23127 10767
rect 23387 10733 23483 10767
rect 23031 10671 23065 10733
rect 20978 10650 21058 10670
rect 11548 10630 11688 10650
rect 11548 10590 11558 10630
rect 11598 10590 11638 10630
rect 11678 10590 11688 10630
rect 11548 10530 11688 10590
rect 11548 10490 11558 10530
rect 11598 10490 11638 10530
rect 11678 10490 11688 10530
rect 11548 10430 11688 10490
rect 11548 10390 11558 10430
rect 11598 10390 11638 10430
rect 11678 10390 11688 10430
rect 11548 10330 11688 10390
rect 11548 10290 11558 10330
rect 11598 10290 11638 10330
rect 11678 10290 11688 10330
rect 11548 10230 11688 10290
rect 11548 10190 11558 10230
rect 11598 10190 11638 10230
rect 11678 10190 11688 10230
rect 11548 10130 11688 10190
rect 11548 10090 11558 10130
rect 11598 10090 11638 10130
rect 11678 10090 11688 10130
rect 11548 10070 11688 10090
rect 11808 10630 11868 10650
rect 11808 10590 11818 10630
rect 11858 10590 11868 10630
rect 11808 10530 11868 10590
rect 11808 10490 11818 10530
rect 11858 10490 11868 10530
rect 11808 10430 11868 10490
rect 11808 10390 11818 10430
rect 11858 10390 11868 10430
rect 11808 10330 11868 10390
rect 11808 10290 11818 10330
rect 11858 10290 11868 10330
rect 11808 10230 11868 10290
rect 11808 10190 11818 10230
rect 11858 10190 11868 10230
rect 11808 10130 11868 10190
rect 11808 10090 11818 10130
rect 11858 10090 11868 10130
rect 11808 10070 11868 10090
rect 11988 10630 12048 10650
rect 11988 10590 11998 10630
rect 12038 10590 12048 10630
rect 11988 10530 12048 10590
rect 11988 10490 11998 10530
rect 12038 10490 12048 10530
rect 11988 10430 12048 10490
rect 11988 10390 11998 10430
rect 12038 10390 12048 10430
rect 11988 10330 12048 10390
rect 11988 10290 11998 10330
rect 12038 10290 12048 10330
rect 11988 10230 12048 10290
rect 11988 10190 11998 10230
rect 12038 10190 12048 10230
rect 11988 10130 12048 10190
rect 11988 10090 11998 10130
rect 12038 10090 12048 10130
rect 11988 10070 12048 10090
rect 12168 10630 12228 10650
rect 12168 10590 12178 10630
rect 12218 10590 12228 10630
rect 12168 10530 12228 10590
rect 12168 10490 12178 10530
rect 12218 10490 12228 10530
rect 12168 10430 12228 10490
rect 12168 10390 12178 10430
rect 12218 10390 12228 10430
rect 12168 10330 12228 10390
rect 12168 10290 12178 10330
rect 12218 10290 12228 10330
rect 12168 10230 12228 10290
rect 12168 10190 12178 10230
rect 12218 10190 12228 10230
rect 12168 10130 12228 10190
rect 12168 10090 12178 10130
rect 12218 10090 12228 10130
rect 12168 10070 12228 10090
rect 12348 10630 12408 10650
rect 12348 10590 12358 10630
rect 12398 10590 12408 10630
rect 12348 10530 12408 10590
rect 12348 10490 12358 10530
rect 12398 10490 12408 10530
rect 12348 10430 12408 10490
rect 12348 10390 12358 10430
rect 12398 10390 12408 10430
rect 12348 10330 12408 10390
rect 12348 10290 12358 10330
rect 12398 10290 12408 10330
rect 12348 10230 12408 10290
rect 12348 10190 12358 10230
rect 12398 10190 12408 10230
rect 12348 10130 12408 10190
rect 12348 10090 12358 10130
rect 12398 10090 12408 10130
rect 12348 10070 12408 10090
rect 12528 10630 12588 10650
rect 12528 10590 12538 10630
rect 12578 10590 12588 10630
rect 12528 10530 12588 10590
rect 12528 10490 12538 10530
rect 12578 10490 12588 10530
rect 12528 10430 12588 10490
rect 12528 10390 12538 10430
rect 12578 10390 12588 10430
rect 12528 10330 12588 10390
rect 12528 10290 12538 10330
rect 12578 10290 12588 10330
rect 12528 10230 12588 10290
rect 12528 10190 12538 10230
rect 12578 10190 12588 10230
rect 12528 10130 12588 10190
rect 12528 10090 12538 10130
rect 12578 10090 12588 10130
rect 12528 10070 12588 10090
rect 12708 10630 12768 10650
rect 12708 10590 12718 10630
rect 12758 10590 12768 10630
rect 12708 10530 12768 10590
rect 12708 10490 12718 10530
rect 12758 10490 12768 10530
rect 12708 10430 12768 10490
rect 12708 10390 12718 10430
rect 12758 10390 12768 10430
rect 12708 10330 12768 10390
rect 12708 10290 12718 10330
rect 12758 10290 12768 10330
rect 12708 10230 12768 10290
rect 12708 10190 12718 10230
rect 12758 10190 12768 10230
rect 12708 10130 12768 10190
rect 12708 10090 12718 10130
rect 12758 10090 12768 10130
rect 12708 10070 12768 10090
rect 12888 10630 12948 10650
rect 12888 10590 12898 10630
rect 12938 10590 12948 10630
rect 12888 10530 12948 10590
rect 12888 10490 12898 10530
rect 12938 10490 12948 10530
rect 12888 10430 12948 10490
rect 12888 10390 12898 10430
rect 12938 10390 12948 10430
rect 12888 10330 12948 10390
rect 12888 10290 12898 10330
rect 12938 10290 12948 10330
rect 12888 10230 12948 10290
rect 12888 10190 12898 10230
rect 12938 10190 12948 10230
rect 12888 10130 12948 10190
rect 12888 10090 12898 10130
rect 12938 10090 12948 10130
rect 12888 10070 12948 10090
rect 13068 10630 13128 10650
rect 13068 10590 13078 10630
rect 13118 10590 13128 10630
rect 13068 10530 13128 10590
rect 13068 10490 13078 10530
rect 13118 10490 13128 10530
rect 13068 10430 13128 10490
rect 13068 10390 13078 10430
rect 13118 10390 13128 10430
rect 13068 10330 13128 10390
rect 13068 10290 13078 10330
rect 13118 10290 13128 10330
rect 13068 10230 13128 10290
rect 13068 10190 13078 10230
rect 13118 10190 13128 10230
rect 13068 10130 13128 10190
rect 13068 10090 13078 10130
rect 13118 10090 13128 10130
rect 13068 10070 13128 10090
rect 13248 10630 13308 10650
rect 13248 10590 13258 10630
rect 13298 10590 13308 10630
rect 13248 10530 13308 10590
rect 13248 10490 13258 10530
rect 13298 10490 13308 10530
rect 13248 10430 13308 10490
rect 13248 10390 13258 10430
rect 13298 10390 13308 10430
rect 13248 10330 13308 10390
rect 13248 10290 13258 10330
rect 13298 10290 13308 10330
rect 13248 10230 13308 10290
rect 13248 10190 13258 10230
rect 13298 10190 13308 10230
rect 13248 10130 13308 10190
rect 13248 10090 13258 10130
rect 13298 10090 13308 10130
rect 13248 10070 13308 10090
rect 13428 10630 13488 10650
rect 13428 10590 13438 10630
rect 13478 10590 13488 10630
rect 13428 10530 13488 10590
rect 13428 10490 13438 10530
rect 13478 10490 13488 10530
rect 13428 10430 13488 10490
rect 13428 10390 13438 10430
rect 13478 10390 13488 10430
rect 13428 10330 13488 10390
rect 13428 10290 13438 10330
rect 13478 10290 13488 10330
rect 13428 10230 13488 10290
rect 13428 10190 13438 10230
rect 13478 10190 13488 10230
rect 13428 10130 13488 10190
rect 13428 10090 13438 10130
rect 13478 10090 13488 10130
rect 13428 10070 13488 10090
rect 13608 10630 13668 10650
rect 13608 10590 13618 10630
rect 13658 10590 13668 10630
rect 13608 10530 13668 10590
rect 13608 10490 13618 10530
rect 13658 10490 13668 10530
rect 13608 10430 13668 10490
rect 13608 10390 13618 10430
rect 13658 10390 13668 10430
rect 13608 10330 13668 10390
rect 13608 10290 13618 10330
rect 13658 10290 13668 10330
rect 13608 10230 13668 10290
rect 13608 10190 13618 10230
rect 13658 10190 13668 10230
rect 13608 10130 13668 10190
rect 13608 10090 13618 10130
rect 13658 10090 13668 10130
rect 13608 10070 13668 10090
rect 13788 10630 13848 10650
rect 13788 10590 13798 10630
rect 13838 10590 13848 10630
rect 13788 10530 13848 10590
rect 13788 10490 13798 10530
rect 13838 10490 13848 10530
rect 13788 10430 13848 10490
rect 13788 10390 13798 10430
rect 13838 10390 13848 10430
rect 13788 10330 13848 10390
rect 13788 10290 13798 10330
rect 13838 10290 13848 10330
rect 13788 10230 13848 10290
rect 13788 10190 13798 10230
rect 13838 10190 13848 10230
rect 13788 10130 13848 10190
rect 13788 10090 13798 10130
rect 13838 10090 13848 10130
rect 13788 10070 13848 10090
rect 13968 10630 14028 10650
rect 13968 10590 13978 10630
rect 14018 10590 14028 10630
rect 13968 10530 14028 10590
rect 13968 10490 13978 10530
rect 14018 10490 14028 10530
rect 13968 10430 14028 10490
rect 13968 10390 13978 10430
rect 14018 10390 14028 10430
rect 13968 10330 14028 10390
rect 13968 10290 13978 10330
rect 14018 10290 14028 10330
rect 13968 10230 14028 10290
rect 13968 10190 13978 10230
rect 14018 10190 14028 10230
rect 13968 10130 14028 10190
rect 13968 10090 13978 10130
rect 14018 10090 14028 10130
rect 13968 10070 14028 10090
rect 14148 10630 14208 10650
rect 14148 10590 14158 10630
rect 14198 10590 14208 10630
rect 14148 10530 14208 10590
rect 14148 10490 14158 10530
rect 14198 10490 14208 10530
rect 14148 10430 14208 10490
rect 14148 10390 14158 10430
rect 14198 10390 14208 10430
rect 14148 10330 14208 10390
rect 14148 10290 14158 10330
rect 14198 10290 14208 10330
rect 14148 10230 14208 10290
rect 14148 10190 14158 10230
rect 14198 10190 14208 10230
rect 14148 10130 14208 10190
rect 14148 10090 14158 10130
rect 14198 10090 14208 10130
rect 14148 10070 14208 10090
rect 14328 10630 14388 10650
rect 14328 10590 14338 10630
rect 14378 10590 14388 10630
rect 14328 10530 14388 10590
rect 14328 10490 14338 10530
rect 14378 10490 14388 10530
rect 14328 10430 14388 10490
rect 14328 10390 14338 10430
rect 14378 10390 14388 10430
rect 14328 10330 14388 10390
rect 14328 10290 14338 10330
rect 14378 10290 14388 10330
rect 14328 10230 14388 10290
rect 14328 10190 14338 10230
rect 14378 10190 14388 10230
rect 14328 10130 14388 10190
rect 14328 10090 14338 10130
rect 14378 10090 14388 10130
rect 14328 10070 14388 10090
rect 14508 10630 14568 10650
rect 14508 10590 14518 10630
rect 14558 10590 14568 10630
rect 14508 10530 14568 10590
rect 14508 10490 14518 10530
rect 14558 10490 14568 10530
rect 14508 10430 14568 10490
rect 14508 10390 14518 10430
rect 14558 10390 14568 10430
rect 14508 10330 14568 10390
rect 14508 10290 14518 10330
rect 14558 10290 14568 10330
rect 14508 10230 14568 10290
rect 14508 10190 14518 10230
rect 14558 10190 14568 10230
rect 14508 10130 14568 10190
rect 14508 10090 14518 10130
rect 14558 10090 14568 10130
rect 14508 10070 14568 10090
rect 14688 10630 14748 10650
rect 14688 10590 14698 10630
rect 14738 10590 14748 10630
rect 14688 10530 14748 10590
rect 14688 10490 14698 10530
rect 14738 10490 14748 10530
rect 14688 10430 14748 10490
rect 14688 10390 14698 10430
rect 14738 10390 14748 10430
rect 14688 10330 14748 10390
rect 14688 10290 14698 10330
rect 14738 10290 14748 10330
rect 14688 10230 14748 10290
rect 14688 10190 14698 10230
rect 14738 10190 14748 10230
rect 14688 10130 14748 10190
rect 14688 10090 14698 10130
rect 14738 10090 14748 10130
rect 14688 10070 14748 10090
rect 14868 10630 15008 10650
rect 14868 10590 14878 10630
rect 14918 10590 14958 10630
rect 14998 10590 15008 10630
rect 14868 10530 15008 10590
rect 19398 10610 19478 10630
rect 19398 10570 19418 10610
rect 19458 10570 19478 10610
rect 20978 10610 20998 10650
rect 21038 10610 21058 10650
rect 20978 10590 21058 10610
rect 14868 10490 14878 10530
rect 14918 10490 14958 10530
rect 14998 10490 15008 10530
rect 15588 10550 15668 10570
rect 15588 10510 15608 10550
rect 15648 10510 15668 10550
rect 15588 10490 15668 10510
rect 15708 10550 15788 10570
rect 15708 10510 15728 10550
rect 15768 10510 15788 10550
rect 15708 10490 15788 10510
rect 15828 10550 15908 10570
rect 19398 10550 19478 10570
rect 19818 10550 21058 10590
rect 21398 10610 21478 10630
rect 21398 10570 21418 10610
rect 21458 10570 21478 10610
rect 21398 10550 21478 10570
rect 15828 10510 15848 10550
rect 15888 10510 15908 10550
rect 19418 10510 19458 10550
rect 19818 10510 19858 10550
rect 21018 10510 21058 10550
rect 21418 10510 21458 10550
rect 15828 10490 15908 10510
rect 19298 10490 19478 10510
rect 14868 10430 15008 10490
rect 14868 10390 14878 10430
rect 14918 10390 14958 10430
rect 14998 10390 15008 10430
rect 14868 10330 15008 10390
rect 14868 10290 14878 10330
rect 14918 10290 14958 10330
rect 14998 10290 15008 10330
rect 14868 10230 15008 10290
rect 15408 10430 15558 10450
rect 15408 10390 15418 10430
rect 15458 10390 15508 10430
rect 15548 10390 15558 10430
rect 15408 10330 15558 10390
rect 15408 10290 15418 10330
rect 15458 10290 15508 10330
rect 15548 10290 15558 10330
rect 15408 10270 15558 10290
rect 15608 10430 15668 10450
rect 15608 10390 15618 10430
rect 15658 10390 15668 10430
rect 15608 10330 15668 10390
rect 15608 10290 15618 10330
rect 15658 10290 15668 10330
rect 15608 10270 15668 10290
rect 15718 10430 15778 10450
rect 15718 10390 15728 10430
rect 15768 10390 15778 10430
rect 15718 10330 15778 10390
rect 15718 10290 15728 10330
rect 15768 10290 15778 10330
rect 15718 10270 15778 10290
rect 15828 10430 15888 10450
rect 15828 10390 15838 10430
rect 15878 10390 15888 10430
rect 15828 10330 15888 10390
rect 15828 10290 15838 10330
rect 15878 10290 15888 10330
rect 15828 10270 15888 10290
rect 15938 10430 16078 10450
rect 15938 10390 15948 10430
rect 15988 10390 16028 10430
rect 16068 10390 16078 10430
rect 15938 10330 16078 10390
rect 15938 10290 15948 10330
rect 15988 10290 16028 10330
rect 16068 10290 16078 10330
rect 15938 10270 16078 10290
rect 19298 10440 19318 10490
rect 19358 10440 19418 10490
rect 19458 10440 19478 10490
rect 19298 10350 19478 10440
rect 19298 10300 19318 10350
rect 19358 10300 19418 10350
rect 19458 10300 19478 10350
rect 19298 10280 19478 10300
rect 19598 10490 19678 10510
rect 19598 10440 19618 10490
rect 19658 10440 19678 10490
rect 19598 10350 19678 10440
rect 19598 10300 19618 10350
rect 19658 10300 19678 10350
rect 19598 10280 19678 10300
rect 19798 10490 19878 10510
rect 19798 10440 19818 10490
rect 19858 10440 19878 10490
rect 19798 10350 19878 10440
rect 19798 10300 19818 10350
rect 19858 10300 19878 10350
rect 19798 10280 19878 10300
rect 19998 10490 20078 10510
rect 19998 10440 20018 10490
rect 20058 10440 20078 10490
rect 19998 10350 20078 10440
rect 19998 10300 20018 10350
rect 20058 10300 20078 10350
rect 19998 10280 20078 10300
rect 20198 10490 20278 10510
rect 20198 10440 20218 10490
rect 20258 10440 20278 10490
rect 20198 10350 20278 10440
rect 20198 10300 20218 10350
rect 20258 10300 20278 10350
rect 20198 10280 20278 10300
rect 20398 10490 20478 10510
rect 20398 10440 20418 10490
rect 20458 10440 20478 10490
rect 20398 10350 20478 10440
rect 20398 10300 20418 10350
rect 20458 10300 20478 10350
rect 20398 10280 20478 10300
rect 20598 10490 20678 10510
rect 20598 10440 20618 10490
rect 20658 10440 20678 10490
rect 20598 10350 20678 10440
rect 20598 10300 20618 10350
rect 20658 10300 20678 10350
rect 20598 10280 20678 10300
rect 20798 10490 20878 10510
rect 20798 10440 20818 10490
rect 20858 10440 20878 10490
rect 20798 10350 20878 10440
rect 20798 10300 20818 10350
rect 20858 10300 20878 10350
rect 20798 10280 20878 10300
rect 20998 10490 21078 10510
rect 20998 10440 21018 10490
rect 21058 10440 21078 10490
rect 20998 10350 21078 10440
rect 20998 10300 21018 10350
rect 21058 10300 21078 10350
rect 20998 10280 21078 10300
rect 21198 10490 21278 10510
rect 21198 10440 21218 10490
rect 21258 10440 21278 10490
rect 21198 10350 21278 10440
rect 21198 10300 21218 10350
rect 21258 10300 21278 10350
rect 21198 10280 21278 10300
rect 21398 10490 21578 10510
rect 21398 10440 21418 10490
rect 21458 10440 21518 10490
rect 21558 10440 21578 10490
rect 21398 10350 21578 10440
rect 21398 10300 21418 10350
rect 21458 10300 21518 10350
rect 21558 10300 21578 10350
rect 21398 10280 21578 10300
rect 20218 10240 20258 10280
rect 20618 10240 20658 10280
rect 14868 10190 14878 10230
rect 14918 10190 14958 10230
rect 14998 10190 15008 10230
rect 14868 10130 15008 10190
rect 15488 10210 15568 10230
rect 15488 10170 15508 10210
rect 15548 10170 15568 10210
rect 15488 10150 15568 10170
rect 15708 10210 15788 10230
rect 15708 10170 15728 10210
rect 15768 10170 15788 10210
rect 15708 10150 15788 10170
rect 15938 10210 15998 10230
rect 15938 10170 15948 10210
rect 15988 10170 15998 10210
rect 15938 10150 15998 10170
rect 20198 10220 20678 10240
rect 20198 10180 20218 10220
rect 20258 10180 20618 10220
rect 20658 10180 20678 10220
rect 20198 10160 20678 10180
rect 14868 10090 14878 10130
rect 14918 10090 14958 10130
rect 14998 10090 15008 10130
rect 14868 10070 15008 10090
rect 11638 10030 11678 10070
rect 11998 10030 12038 10070
rect 12358 10030 12398 10070
rect 12718 10030 12758 10070
rect 13078 10030 13118 10070
rect 13438 10030 13478 10070
rect 13798 10030 13838 10070
rect 14158 10030 14198 10070
rect 14518 10030 14558 10070
rect 14878 10030 14918 10070
rect 19138 10040 19258 10050
rect 20588 10040 20678 10160
rect 19138 10030 19292 10040
rect 11618 10010 11698 10030
rect 11618 9970 11638 10010
rect 11678 9970 11698 10010
rect 11618 9950 11698 9970
rect 11978 10010 12058 10030
rect 11978 9970 11998 10010
rect 12038 9970 12058 10010
rect 11978 9950 12058 9970
rect 12338 10010 12418 10030
rect 12338 9970 12358 10010
rect 12398 9970 12418 10010
rect 12338 9950 12418 9970
rect 12698 10010 12778 10030
rect 12698 9970 12718 10010
rect 12758 9970 12778 10010
rect 12698 9950 12778 9970
rect 13058 10010 13138 10030
rect 13058 9970 13078 10010
rect 13118 9970 13138 10010
rect 13058 9950 13138 9970
rect 13418 10010 13498 10030
rect 13418 9970 13438 10010
rect 13478 9970 13498 10010
rect 13418 9950 13498 9970
rect 13778 10010 13858 10030
rect 13778 9970 13798 10010
rect 13838 9970 13858 10010
rect 13778 9950 13858 9970
rect 14138 10010 14218 10030
rect 14138 9970 14158 10010
rect 14198 9970 14218 10010
rect 14138 9950 14218 9970
rect 14498 10010 14578 10030
rect 14498 9970 14518 10010
rect 14558 9970 14578 10010
rect 14498 9950 14578 9970
rect 14858 10010 14938 10030
rect 14858 9970 14878 10010
rect 14918 9970 14938 10010
rect 19138 9990 19158 10030
rect 19198 10024 19292 10030
rect 19198 9990 19258 10024
rect 19138 9974 19292 9990
rect 20532 10024 20678 10040
rect 20566 9990 20678 10024
rect 20532 9974 20678 9990
rect 19138 9970 19258 9974
rect 20558 9970 20678 9974
rect 14858 9950 14938 9970
rect 11804 9742 11862 9760
rect 11804 9708 11816 9742
rect 11850 9708 11862 9742
rect 11804 9690 11862 9708
rect 11914 9742 11972 9760
rect 11914 9708 11926 9742
rect 11960 9708 11972 9742
rect 11914 9690 11972 9708
rect 12024 9742 12082 9760
rect 12024 9708 12036 9742
rect 12070 9708 12082 9742
rect 12024 9690 12082 9708
rect 12134 9742 12192 9760
rect 12134 9708 12146 9742
rect 12180 9708 12192 9742
rect 12134 9690 12192 9708
rect 12244 9742 12302 9760
rect 12244 9708 12256 9742
rect 12290 9708 12302 9742
rect 12244 9690 12302 9708
rect 12354 9742 12412 9760
rect 12354 9708 12366 9742
rect 12400 9708 12412 9742
rect 12354 9690 12412 9708
rect 12464 9742 12522 9760
rect 12464 9708 12476 9742
rect 12510 9708 12522 9742
rect 12464 9690 12522 9708
rect 12574 9742 12632 9760
rect 12574 9708 12586 9742
rect 12620 9708 12632 9742
rect 12574 9690 12632 9708
rect 12684 9742 12742 9760
rect 12684 9708 12696 9742
rect 12730 9708 12742 9742
rect 12684 9690 12742 9708
rect 12794 9742 12852 9760
rect 12794 9708 12806 9742
rect 12840 9708 12852 9742
rect 12794 9690 12852 9708
rect 13704 9742 13762 9760
rect 13704 9708 13716 9742
rect 13750 9708 13762 9742
rect 13704 9690 13762 9708
rect 13814 9742 13872 9760
rect 13814 9708 13826 9742
rect 13860 9708 13872 9742
rect 13814 9690 13872 9708
rect 13924 9742 13982 9760
rect 13924 9708 13936 9742
rect 13970 9708 13982 9742
rect 13924 9690 13982 9708
rect 14034 9742 14092 9760
rect 14034 9708 14046 9742
rect 14080 9708 14092 9742
rect 14034 9690 14092 9708
rect 14144 9742 14202 9760
rect 14144 9708 14156 9742
rect 14190 9708 14202 9742
rect 14144 9690 14202 9708
rect 14254 9742 14312 9760
rect 14254 9708 14266 9742
rect 14300 9708 14312 9742
rect 14254 9690 14312 9708
rect 14364 9742 14422 9760
rect 14364 9708 14376 9742
rect 14410 9708 14422 9742
rect 14364 9690 14422 9708
rect 14474 9742 14532 9760
rect 14474 9708 14486 9742
rect 14520 9708 14532 9742
rect 14474 9690 14532 9708
rect 14584 9742 14642 9760
rect 14584 9708 14596 9742
rect 14630 9708 14642 9742
rect 14584 9690 14642 9708
rect 14694 9742 14752 9760
rect 14694 9708 14706 9742
rect 14740 9708 14752 9742
rect 14694 9690 14752 9708
rect 11558 9630 11698 9650
rect 11558 9590 11568 9630
rect 11608 9590 11648 9630
rect 11688 9590 11698 9630
rect 11558 9530 11698 9590
rect 11558 9490 11568 9530
rect 11608 9490 11648 9530
rect 11688 9490 11698 9530
rect 11558 9470 11698 9490
rect 11748 9630 11808 9650
rect 11748 9590 11758 9630
rect 11798 9590 11808 9630
rect 11748 9530 11808 9590
rect 11748 9490 11758 9530
rect 11798 9490 11808 9530
rect 11748 9470 11808 9490
rect 11858 9630 11918 9650
rect 11858 9590 11868 9630
rect 11908 9590 11918 9630
rect 11858 9530 11918 9590
rect 11858 9490 11868 9530
rect 11908 9490 11918 9530
rect 11858 9470 11918 9490
rect 11968 9630 12028 9650
rect 11968 9590 11978 9630
rect 12018 9590 12028 9630
rect 11968 9530 12028 9590
rect 11968 9490 11978 9530
rect 12018 9490 12028 9530
rect 11968 9470 12028 9490
rect 12078 9630 12138 9650
rect 12078 9590 12088 9630
rect 12128 9590 12138 9630
rect 12078 9530 12138 9590
rect 12078 9490 12088 9530
rect 12128 9490 12138 9530
rect 12078 9470 12138 9490
rect 12188 9630 12248 9650
rect 12188 9590 12198 9630
rect 12238 9590 12248 9630
rect 12188 9530 12248 9590
rect 12188 9490 12198 9530
rect 12238 9490 12248 9530
rect 12188 9470 12248 9490
rect 12298 9630 12358 9650
rect 12298 9590 12308 9630
rect 12348 9590 12358 9630
rect 12298 9530 12358 9590
rect 12298 9490 12308 9530
rect 12348 9490 12358 9530
rect 12298 9470 12358 9490
rect 12408 9630 12468 9650
rect 12408 9590 12418 9630
rect 12458 9590 12468 9630
rect 12408 9530 12468 9590
rect 12408 9490 12418 9530
rect 12458 9490 12468 9530
rect 12408 9470 12468 9490
rect 12518 9630 12578 9650
rect 12518 9590 12528 9630
rect 12568 9590 12578 9630
rect 12518 9530 12578 9590
rect 12518 9490 12528 9530
rect 12568 9490 12578 9530
rect 12518 9470 12578 9490
rect 12628 9630 12688 9650
rect 12628 9590 12638 9630
rect 12678 9590 12688 9630
rect 12628 9530 12688 9590
rect 12628 9490 12638 9530
rect 12678 9490 12688 9530
rect 12628 9470 12688 9490
rect 12738 9630 12798 9650
rect 12738 9590 12748 9630
rect 12788 9590 12798 9630
rect 12738 9530 12798 9590
rect 12738 9490 12748 9530
rect 12788 9490 12798 9530
rect 12738 9470 12798 9490
rect 12848 9630 12908 9650
rect 12848 9590 12858 9630
rect 12898 9590 12908 9630
rect 12848 9530 12908 9590
rect 12848 9490 12858 9530
rect 12898 9490 12908 9530
rect 12848 9470 12908 9490
rect 12958 9630 13098 9650
rect 12958 9590 12968 9630
rect 13008 9590 13048 9630
rect 13088 9590 13098 9630
rect 12958 9530 13098 9590
rect 12958 9490 12968 9530
rect 13008 9490 13048 9530
rect 13088 9490 13098 9530
rect 12958 9470 13098 9490
rect 13458 9630 13598 9650
rect 13458 9590 13468 9630
rect 13508 9590 13548 9630
rect 13588 9590 13598 9630
rect 13458 9530 13598 9590
rect 13458 9490 13468 9530
rect 13508 9490 13548 9530
rect 13588 9490 13598 9530
rect 13458 9470 13598 9490
rect 13648 9630 13708 9650
rect 13648 9590 13658 9630
rect 13698 9590 13708 9630
rect 13648 9530 13708 9590
rect 13648 9490 13658 9530
rect 13698 9490 13708 9530
rect 13648 9470 13708 9490
rect 13758 9630 13818 9650
rect 13758 9590 13768 9630
rect 13808 9590 13818 9630
rect 13758 9530 13818 9590
rect 13758 9490 13768 9530
rect 13808 9490 13818 9530
rect 13758 9470 13818 9490
rect 13868 9630 13928 9650
rect 13868 9590 13878 9630
rect 13918 9590 13928 9630
rect 13868 9530 13928 9590
rect 13868 9490 13878 9530
rect 13918 9490 13928 9530
rect 13868 9470 13928 9490
rect 13978 9630 14038 9650
rect 13978 9590 13988 9630
rect 14028 9590 14038 9630
rect 13978 9530 14038 9590
rect 13978 9490 13988 9530
rect 14028 9490 14038 9530
rect 13978 9470 14038 9490
rect 14088 9630 14148 9650
rect 14088 9590 14098 9630
rect 14138 9590 14148 9630
rect 14088 9530 14148 9590
rect 14088 9490 14098 9530
rect 14138 9490 14148 9530
rect 14088 9470 14148 9490
rect 14198 9630 14258 9650
rect 14198 9590 14208 9630
rect 14248 9590 14258 9630
rect 14198 9530 14258 9590
rect 14198 9490 14208 9530
rect 14248 9490 14258 9530
rect 14198 9470 14258 9490
rect 14308 9630 14368 9650
rect 14308 9590 14318 9630
rect 14358 9590 14368 9630
rect 14308 9530 14368 9590
rect 14308 9490 14318 9530
rect 14358 9490 14368 9530
rect 14308 9470 14368 9490
rect 14418 9630 14478 9650
rect 14418 9590 14428 9630
rect 14468 9590 14478 9630
rect 14418 9530 14478 9590
rect 14418 9490 14428 9530
rect 14468 9490 14478 9530
rect 14418 9470 14478 9490
rect 14528 9630 14588 9650
rect 14528 9590 14538 9630
rect 14578 9590 14588 9630
rect 14528 9530 14588 9590
rect 14528 9490 14538 9530
rect 14578 9490 14588 9530
rect 14528 9470 14588 9490
rect 14638 9630 14698 9650
rect 14638 9590 14648 9630
rect 14688 9590 14698 9630
rect 14638 9530 14698 9590
rect 14638 9490 14648 9530
rect 14688 9490 14698 9530
rect 14638 9470 14698 9490
rect 14748 9630 14808 9650
rect 14748 9590 14758 9630
rect 14798 9590 14808 9630
rect 14748 9530 14808 9590
rect 14748 9490 14758 9530
rect 14798 9490 14808 9530
rect 14748 9470 14808 9490
rect 14858 9630 14998 9650
rect 14858 9590 14868 9630
rect 14908 9590 14948 9630
rect 14988 9590 14998 9630
rect 14858 9530 14998 9590
rect 23008 9640 23031 9660
rect 23449 10671 23483 10733
rect 23065 9640 23088 9660
rect 23008 9600 23028 9640
rect 23068 9600 23088 9640
rect 23008 9581 23031 9600
rect 23065 9581 23088 9600
rect 23008 9580 23088 9581
rect 14858 9490 14868 9530
rect 14908 9490 14948 9530
rect 14988 9490 14998 9530
rect 14858 9470 14998 9490
rect 23031 9519 23065 9580
rect 23449 9519 23483 9581
rect 23031 9485 23127 9519
rect 23387 9485 23483 9519
rect 11628 9410 11708 9430
rect 11628 9370 11648 9410
rect 11688 9370 11708 9410
rect 11628 9350 11708 9370
rect 12948 9410 13028 9430
rect 12948 9370 12968 9410
rect 13008 9370 13028 9410
rect 12948 9350 13028 9370
rect 13528 9410 13608 9430
rect 13528 9370 13548 9410
rect 13588 9370 13608 9410
rect 13528 9350 13608 9370
rect 14848 9410 14928 9430
rect 14848 9370 14868 9410
rect 14908 9370 14928 9410
rect 14848 9350 14928 9370
rect 23208 9130 23308 9150
rect 23208 9070 23228 9130
rect 23288 9070 23308 9130
rect 23208 9050 23308 9070
rect 23088 8380 23198 8400
rect 23088 8310 23108 8380
rect 23178 8310 23198 8380
rect 13248 8290 13328 8310
rect 13248 8250 13268 8290
rect 13308 8250 13328 8290
rect 13248 8230 13328 8250
rect 13468 8290 13548 8310
rect 13468 8250 13488 8290
rect 13528 8250 13548 8290
rect 13468 8230 13548 8250
rect 13768 8290 13848 8310
rect 13768 8250 13788 8290
rect 13828 8250 13848 8290
rect 13768 8230 13848 8250
rect 13998 8290 14078 8310
rect 13998 8250 14018 8290
rect 14058 8250 14078 8290
rect 13998 8230 14078 8250
rect 14148 8290 14228 8310
rect 14148 8250 14168 8290
rect 14208 8250 14228 8290
rect 14148 8230 14228 8250
rect 14368 8290 14448 8310
rect 14368 8250 14388 8290
rect 14428 8250 14448 8290
rect 14368 8230 14448 8250
rect 14668 8290 14748 8310
rect 14668 8250 14688 8290
rect 14728 8250 14748 8290
rect 14668 8230 14748 8250
rect 14888 8290 14968 8310
rect 14888 8250 14908 8290
rect 14948 8250 14968 8290
rect 14888 8230 14968 8250
rect 15288 8290 15368 8310
rect 15288 8250 15308 8290
rect 15348 8250 15368 8290
rect 15288 8230 15368 8250
rect 15618 8290 15698 8310
rect 15618 8250 15638 8290
rect 15678 8250 15698 8290
rect 15618 8230 15698 8250
rect 15948 8290 16028 8310
rect 15948 8250 15968 8290
rect 16008 8250 16028 8290
rect 15948 8230 16028 8250
rect 16388 8290 16468 8310
rect 16388 8250 16408 8290
rect 16448 8250 16468 8290
rect 16388 8230 16468 8250
rect 17168 8290 17248 8310
rect 17168 8250 17188 8290
rect 17228 8250 17248 8290
rect 17168 8230 17248 8250
rect 17848 8290 17928 8310
rect 23088 8290 23198 8310
rect 17848 8250 17868 8290
rect 17908 8250 17928 8290
rect 17848 8230 17928 8250
rect 13268 8080 13308 8230
rect 13488 8080 13528 8230
rect 13788 8080 13828 8230
rect 14018 8080 14058 8230
rect 14168 8080 14208 8230
rect 14388 8080 14428 8230
rect 14688 8080 14728 8230
rect 14908 8080 14948 8230
rect 15308 8080 15348 8230
rect 15638 8080 15678 8230
rect 15968 8080 16008 8230
rect 16408 8080 16448 8230
rect 16898 8180 16978 8200
rect 16898 8140 16918 8180
rect 16958 8140 16978 8180
rect 16898 8120 16978 8140
rect 17188 8080 17228 8230
rect 17528 8180 17608 8200
rect 17528 8140 17548 8180
rect 17588 8140 17608 8180
rect 17528 8120 17608 8140
rect 17868 8080 17908 8230
rect 19338 8130 19418 8150
rect 19338 8090 19358 8130
rect 19398 8090 19418 8130
rect 13178 8060 13318 8080
rect 13178 8020 13188 8060
rect 13228 8020 13268 8060
rect 13308 8020 13318 8060
rect 13178 7960 13318 8020
rect 13178 7920 13188 7960
rect 13228 7920 13268 7960
rect 13308 7920 13318 7960
rect 13178 7900 13318 7920
rect 13368 8060 13428 8080
rect 13368 8020 13378 8060
rect 13418 8020 13428 8060
rect 13368 7960 13428 8020
rect 13368 7920 13378 7960
rect 13418 7920 13428 7960
rect 13368 7900 13428 7920
rect 13478 8060 13538 8080
rect 13478 8020 13488 8060
rect 13528 8020 13538 8060
rect 13478 7960 13538 8020
rect 13478 7920 13488 7960
rect 13528 7920 13538 7960
rect 13478 7900 13538 7920
rect 13778 8060 13838 8080
rect 13778 8020 13788 8060
rect 13828 8020 13838 8060
rect 13778 7960 13838 8020
rect 13778 7920 13788 7960
rect 13828 7920 13838 7960
rect 13778 7900 13838 7920
rect 13888 8060 13948 8080
rect 13888 8020 13898 8060
rect 13938 8020 13948 8060
rect 13888 7960 13948 8020
rect 13888 7920 13898 7960
rect 13938 7920 13948 7960
rect 13888 7900 13948 7920
rect 13998 8060 14218 8080
rect 13998 8020 14008 8060
rect 14048 8020 14088 8060
rect 14128 8020 14168 8060
rect 14208 8020 14218 8060
rect 13998 7960 14218 8020
rect 13998 7920 14008 7960
rect 14048 7920 14088 7960
rect 14128 7920 14168 7960
rect 14208 7920 14218 7960
rect 13998 7900 14218 7920
rect 14268 8060 14328 8080
rect 14268 8020 14278 8060
rect 14318 8020 14328 8060
rect 14268 7960 14328 8020
rect 14268 7920 14278 7960
rect 14318 7920 14328 7960
rect 14268 7900 14328 7920
rect 14378 8060 14438 8080
rect 14378 8020 14388 8060
rect 14428 8020 14438 8060
rect 14378 7960 14438 8020
rect 14378 7920 14388 7960
rect 14428 7920 14438 7960
rect 14378 7900 14438 7920
rect 14678 8060 14738 8080
rect 14678 8020 14688 8060
rect 14728 8020 14738 8060
rect 14678 7960 14738 8020
rect 14678 7920 14688 7960
rect 14728 7920 14738 7960
rect 14678 7900 14738 7920
rect 14788 8060 14848 8080
rect 14788 8020 14798 8060
rect 14838 8020 14848 8060
rect 14788 7960 14848 8020
rect 14788 7920 14798 7960
rect 14838 7920 14848 7960
rect 14788 7900 14848 7920
rect 14898 8060 15038 8080
rect 14898 8020 14908 8060
rect 14948 8020 14988 8060
rect 15028 8020 15038 8060
rect 14898 7960 15038 8020
rect 14898 7920 14908 7960
rect 14948 7920 14988 7960
rect 15028 7920 15038 7960
rect 14898 7900 15038 7920
rect 15188 8060 15248 8080
rect 15188 8020 15198 8060
rect 15238 8020 15248 8060
rect 15188 7960 15248 8020
rect 15188 7920 15198 7960
rect 15238 7920 15248 7960
rect 15188 7900 15248 7920
rect 15298 8060 15438 8080
rect 15298 8020 15308 8060
rect 15348 8020 15388 8060
rect 15428 8020 15438 8060
rect 15298 7960 15438 8020
rect 15298 7920 15308 7960
rect 15348 7920 15388 7960
rect 15428 7920 15438 7960
rect 15298 7900 15438 7920
rect 15518 8060 15578 8080
rect 15518 8020 15528 8060
rect 15568 8020 15578 8060
rect 15518 7960 15578 8020
rect 15518 7920 15528 7960
rect 15568 7920 15578 7960
rect 15518 7900 15578 7920
rect 15628 8060 15768 8080
rect 15628 8020 15638 8060
rect 15678 8020 15718 8060
rect 15758 8020 15768 8060
rect 15628 7960 15768 8020
rect 15628 7920 15638 7960
rect 15678 7920 15718 7960
rect 15758 7920 15768 7960
rect 15628 7900 15768 7920
rect 15848 8060 15908 8080
rect 15848 8020 15858 8060
rect 15898 8020 15908 8060
rect 15848 7960 15908 8020
rect 15848 7920 15858 7960
rect 15898 7920 15908 7960
rect 15848 7900 15908 7920
rect 15958 8060 16098 8080
rect 15958 8020 15968 8060
rect 16008 8020 16048 8060
rect 16088 8020 16098 8060
rect 15958 7960 16098 8020
rect 15958 7920 15968 7960
rect 16008 7920 16048 7960
rect 16088 7920 16098 7960
rect 15958 7900 16098 7920
rect 16288 8060 16468 8080
rect 16288 8020 16308 8060
rect 16348 8020 16408 8060
rect 16448 8020 16468 8060
rect 16288 7960 16468 8020
rect 16288 7920 16308 7960
rect 16348 7920 16408 7960
rect 16448 7920 16468 7960
rect 16288 7900 16468 7920
rect 16518 8060 16598 8080
rect 16518 8020 16538 8060
rect 16578 8020 16598 8060
rect 16518 7960 16598 8020
rect 16518 7920 16538 7960
rect 16578 7920 16598 7960
rect 16518 7900 16598 7920
rect 16778 8060 16858 8080
rect 16778 8020 16798 8060
rect 16838 8020 16858 8060
rect 16778 7960 16858 8020
rect 16778 7920 16798 7960
rect 16838 7920 16858 7960
rect 16778 7900 16858 7920
rect 16908 8060 16988 8080
rect 16908 8020 16928 8060
rect 16968 8020 16988 8060
rect 16908 7960 16988 8020
rect 16908 7920 16928 7960
rect 16968 7920 16988 7960
rect 16908 7900 16988 7920
rect 17068 8060 17248 8080
rect 17068 8020 17088 8060
rect 17128 8020 17188 8060
rect 17228 8020 17248 8060
rect 17068 7960 17248 8020
rect 17068 7920 17088 7960
rect 17128 7920 17188 7960
rect 17228 7920 17248 7960
rect 17068 7900 17248 7920
rect 17298 8060 17378 8080
rect 17298 8020 17318 8060
rect 17358 8020 17378 8060
rect 17298 7960 17378 8020
rect 17298 7920 17318 7960
rect 17358 7920 17378 7960
rect 17298 7900 17378 7920
rect 17458 8060 17538 8080
rect 17458 8020 17478 8060
rect 17518 8020 17538 8060
rect 17458 7960 17538 8020
rect 17458 7920 17478 7960
rect 17518 7920 17538 7960
rect 17458 7900 17538 7920
rect 17588 8060 17668 8080
rect 17588 8020 17608 8060
rect 17648 8020 17668 8060
rect 17588 7960 17668 8020
rect 17588 7920 17608 7960
rect 17648 7920 17668 7960
rect 17588 7900 17668 7920
rect 17748 8060 17928 8080
rect 17748 8020 17768 8060
rect 17808 8020 17868 8060
rect 17908 8020 17928 8060
rect 17748 7960 17928 8020
rect 17748 7920 17768 7960
rect 17808 7920 17868 7960
rect 17908 7920 17928 7960
rect 17748 7900 17928 7920
rect 17978 8060 18058 8080
rect 19338 8070 19418 8090
rect 22378 8130 22458 8150
rect 22378 8090 22398 8130
rect 22438 8090 22458 8130
rect 22378 8070 22458 8090
rect 17978 8020 17998 8060
rect 18038 8020 18058 8060
rect 17978 7960 18058 8020
rect 17978 7920 17998 7960
rect 18038 7920 18058 7960
rect 17978 7900 18058 7920
rect 19238 8010 19418 8030
rect 19238 7970 19258 8010
rect 19298 7970 19358 8010
rect 19398 7970 19418 8010
rect 19238 7910 19418 7970
rect 13128 7800 13208 7820
rect 13128 7760 13148 7800
rect 13188 7760 13208 7800
rect 13128 7740 13208 7760
rect 13368 7740 13408 7900
rect 13458 7840 13538 7860
rect 13458 7800 13478 7840
rect 13518 7820 13538 7840
rect 13518 7800 13738 7820
rect 13458 7780 13738 7800
rect 13368 7700 13528 7740
rect 13488 7660 13528 7700
rect 13178 7640 13318 7660
rect 13178 7600 13188 7640
rect 13228 7600 13268 7640
rect 13308 7600 13318 7640
rect 13178 7540 13318 7600
rect 13178 7500 13188 7540
rect 13228 7500 13268 7540
rect 13308 7500 13318 7540
rect 13178 7440 13318 7500
rect 13178 7400 13188 7440
rect 13228 7400 13268 7440
rect 13308 7400 13318 7440
rect 13178 7340 13318 7400
rect 13178 7300 13188 7340
rect 13228 7300 13268 7340
rect 13308 7300 13318 7340
rect 13178 7280 13318 7300
rect 13368 7640 13428 7660
rect 13368 7600 13378 7640
rect 13418 7600 13428 7640
rect 13368 7540 13428 7600
rect 13368 7500 13378 7540
rect 13418 7500 13428 7540
rect 13368 7440 13428 7500
rect 13368 7400 13378 7440
rect 13418 7400 13428 7440
rect 13368 7340 13428 7400
rect 13368 7300 13378 7340
rect 13418 7300 13428 7340
rect 13368 7280 13428 7300
rect 13478 7640 13538 7660
rect 13478 7600 13488 7640
rect 13528 7600 13538 7640
rect 13478 7540 13538 7600
rect 13478 7500 13488 7540
rect 13528 7500 13538 7540
rect 13478 7440 13538 7500
rect 13478 7400 13488 7440
rect 13528 7400 13538 7440
rect 13478 7340 13538 7400
rect 13478 7300 13488 7340
rect 13528 7330 13538 7340
rect 13578 7340 13658 7360
rect 13578 7330 13598 7340
rect 13528 7300 13598 7330
rect 13638 7300 13658 7340
rect 13478 7280 13658 7300
rect 13698 7320 13738 7780
rect 13898 7740 13938 7900
rect 13788 7700 13938 7740
rect 13978 7760 14058 7780
rect 13978 7720 13998 7760
rect 14038 7740 14058 7760
rect 14268 7740 14308 7900
rect 14358 7840 14438 7860
rect 14358 7800 14378 7840
rect 14418 7820 14438 7840
rect 14418 7800 14638 7820
rect 14358 7780 14638 7800
rect 14038 7720 14428 7740
rect 13978 7700 14428 7720
rect 13788 7660 13828 7700
rect 14388 7660 14428 7700
rect 13778 7640 13838 7660
rect 13778 7600 13788 7640
rect 13828 7600 13838 7640
rect 13778 7540 13838 7600
rect 13778 7500 13788 7540
rect 13828 7500 13838 7540
rect 13778 7440 13838 7500
rect 13778 7400 13788 7440
rect 13828 7400 13838 7440
rect 13778 7340 13838 7400
rect 13778 7320 13788 7340
rect 13698 7300 13788 7320
rect 13828 7300 13838 7340
rect 13698 7280 13838 7300
rect 13888 7640 13948 7660
rect 13888 7600 13898 7640
rect 13938 7600 13948 7640
rect 13888 7540 13948 7600
rect 13888 7500 13898 7540
rect 13938 7500 13948 7540
rect 13888 7440 13948 7500
rect 13888 7400 13898 7440
rect 13938 7400 13948 7440
rect 13888 7340 13948 7400
rect 13888 7300 13898 7340
rect 13938 7300 13948 7340
rect 13888 7280 13948 7300
rect 13998 7640 14218 7660
rect 13998 7600 14008 7640
rect 14048 7600 14088 7640
rect 14128 7600 14168 7640
rect 14208 7600 14218 7640
rect 13998 7540 14218 7600
rect 13998 7500 14008 7540
rect 14048 7500 14088 7540
rect 14128 7500 14168 7540
rect 14208 7500 14218 7540
rect 13998 7440 14218 7500
rect 13998 7400 14008 7440
rect 14048 7400 14088 7440
rect 14128 7400 14168 7440
rect 14208 7400 14218 7440
rect 13998 7340 14218 7400
rect 13998 7300 14008 7340
rect 14048 7300 14088 7340
rect 14128 7300 14168 7340
rect 14208 7300 14218 7340
rect 13998 7280 14218 7300
rect 14268 7640 14328 7660
rect 14268 7600 14278 7640
rect 14318 7600 14328 7640
rect 14268 7540 14328 7600
rect 14268 7500 14278 7540
rect 14318 7500 14328 7540
rect 14268 7440 14328 7500
rect 14268 7400 14278 7440
rect 14318 7400 14328 7440
rect 14268 7340 14328 7400
rect 14268 7300 14278 7340
rect 14318 7300 14328 7340
rect 14268 7280 14328 7300
rect 14378 7640 14438 7660
rect 14378 7600 14388 7640
rect 14428 7600 14438 7640
rect 14378 7540 14438 7600
rect 14378 7500 14388 7540
rect 14428 7500 14438 7540
rect 14378 7440 14438 7500
rect 14378 7400 14388 7440
rect 14428 7400 14438 7440
rect 14378 7340 14438 7400
rect 14378 7300 14388 7340
rect 14428 7330 14438 7340
rect 14478 7340 14558 7360
rect 14478 7330 14498 7340
rect 14428 7300 14498 7330
rect 14538 7300 14558 7340
rect 14378 7280 14558 7300
rect 14598 7320 14638 7780
rect 14798 7740 14838 7900
rect 15188 7810 15228 7900
rect 15518 7810 15558 7900
rect 15848 7810 15888 7900
rect 14688 7700 14838 7740
rect 15048 7790 15228 7810
rect 15048 7750 15068 7790
rect 15108 7750 15148 7790
rect 15188 7750 15228 7790
rect 15048 7730 15228 7750
rect 15458 7790 15558 7810
rect 15458 7750 15478 7790
rect 15518 7750 15558 7790
rect 15458 7730 15558 7750
rect 15788 7790 15888 7810
rect 15788 7750 15808 7790
rect 15848 7750 15888 7790
rect 15788 7730 15888 7750
rect 16078 7790 16158 7810
rect 16078 7750 16098 7790
rect 16138 7750 16158 7790
rect 16078 7730 16158 7750
rect 16228 7800 16308 7820
rect 16228 7760 16248 7800
rect 16288 7760 16308 7800
rect 16228 7740 16308 7760
rect 16538 7740 16578 7900
rect 16798 7740 16838 7900
rect 14688 7660 14728 7700
rect 15188 7660 15228 7730
rect 15518 7660 15558 7730
rect 15848 7660 15888 7730
rect 16538 7700 16838 7740
rect 16538 7660 16578 7700
rect 16798 7660 16838 7700
rect 16928 7790 16968 7900
rect 17338 7870 17378 7900
rect 17338 7850 17418 7870
rect 17338 7810 17358 7850
rect 17398 7810 17418 7850
rect 17338 7800 17418 7810
rect 16928 7770 17028 7790
rect 16928 7730 16968 7770
rect 17008 7730 17028 7770
rect 16928 7710 17028 7730
rect 16928 7660 16968 7710
rect 17338 7660 17378 7800
rect 17478 7660 17518 7900
rect 17608 7820 17648 7900
rect 17998 7860 18038 7900
rect 19238 7870 19258 7910
rect 19298 7870 19358 7910
rect 19398 7870 19418 7910
rect 17998 7840 18078 7860
rect 17998 7820 18018 7840
rect 17608 7800 18018 7820
rect 18058 7800 18078 7840
rect 17608 7780 18078 7800
rect 19238 7810 19418 7870
rect 17608 7660 17648 7780
rect 19238 7770 19258 7810
rect 19298 7770 19358 7810
rect 19398 7770 19418 7810
rect 19238 7710 19418 7770
rect 19238 7670 19258 7710
rect 19298 7670 19358 7710
rect 19398 7670 19418 7710
rect 14678 7640 14738 7660
rect 14678 7600 14688 7640
rect 14728 7600 14738 7640
rect 14678 7540 14738 7600
rect 14678 7500 14688 7540
rect 14728 7500 14738 7540
rect 14678 7440 14738 7500
rect 14678 7400 14688 7440
rect 14728 7400 14738 7440
rect 14678 7340 14738 7400
rect 14678 7320 14688 7340
rect 14598 7300 14688 7320
rect 14728 7300 14738 7340
rect 14598 7280 14738 7300
rect 14788 7640 14848 7660
rect 14788 7600 14798 7640
rect 14838 7600 14848 7640
rect 14788 7540 14848 7600
rect 14788 7500 14798 7540
rect 14838 7500 14848 7540
rect 14788 7440 14848 7500
rect 14788 7400 14798 7440
rect 14838 7400 14848 7440
rect 14788 7340 14848 7400
rect 14788 7300 14798 7340
rect 14838 7300 14848 7340
rect 14788 7280 14848 7300
rect 14898 7640 15038 7660
rect 14898 7600 14908 7640
rect 14948 7600 14988 7640
rect 15028 7600 15038 7640
rect 14898 7540 15038 7600
rect 14898 7500 14908 7540
rect 14948 7500 14988 7540
rect 15028 7500 15038 7540
rect 14898 7440 15038 7500
rect 14898 7400 14908 7440
rect 14948 7400 14988 7440
rect 15028 7400 15038 7440
rect 14898 7340 15038 7400
rect 14898 7300 14908 7340
rect 14948 7300 14988 7340
rect 15028 7300 15038 7340
rect 14898 7280 15038 7300
rect 15188 7640 15248 7660
rect 15188 7600 15198 7640
rect 15238 7600 15248 7640
rect 15188 7540 15248 7600
rect 15188 7500 15198 7540
rect 15238 7500 15248 7540
rect 15188 7440 15248 7500
rect 15188 7400 15198 7440
rect 15238 7400 15248 7440
rect 15188 7340 15248 7400
rect 15188 7300 15198 7340
rect 15238 7300 15248 7340
rect 15188 7280 15248 7300
rect 15298 7640 15438 7660
rect 15298 7600 15308 7640
rect 15348 7600 15388 7640
rect 15428 7600 15438 7640
rect 15298 7540 15438 7600
rect 15298 7500 15308 7540
rect 15348 7500 15388 7540
rect 15428 7500 15438 7540
rect 15298 7440 15438 7500
rect 15298 7400 15308 7440
rect 15348 7400 15388 7440
rect 15428 7400 15438 7440
rect 15298 7340 15438 7400
rect 15298 7300 15308 7340
rect 15348 7300 15388 7340
rect 15428 7300 15438 7340
rect 15298 7280 15438 7300
rect 15518 7640 15578 7660
rect 15518 7600 15528 7640
rect 15568 7600 15578 7640
rect 15518 7540 15578 7600
rect 15518 7500 15528 7540
rect 15568 7500 15578 7540
rect 15518 7440 15578 7500
rect 15518 7400 15528 7440
rect 15568 7400 15578 7440
rect 15518 7340 15578 7400
rect 15518 7300 15528 7340
rect 15568 7300 15578 7340
rect 15518 7280 15578 7300
rect 15628 7640 15768 7660
rect 15628 7600 15638 7640
rect 15678 7600 15718 7640
rect 15758 7600 15768 7640
rect 15628 7540 15768 7600
rect 15628 7500 15638 7540
rect 15678 7500 15718 7540
rect 15758 7500 15768 7540
rect 15628 7440 15768 7500
rect 15628 7400 15638 7440
rect 15678 7400 15718 7440
rect 15758 7400 15768 7440
rect 15628 7340 15768 7400
rect 15628 7300 15638 7340
rect 15678 7300 15718 7340
rect 15758 7300 15768 7340
rect 15628 7280 15768 7300
rect 15848 7640 15908 7660
rect 15848 7600 15858 7640
rect 15898 7600 15908 7640
rect 15848 7540 15908 7600
rect 15848 7500 15858 7540
rect 15898 7500 15908 7540
rect 15848 7440 15908 7500
rect 15848 7400 15858 7440
rect 15898 7400 15908 7440
rect 15848 7340 15908 7400
rect 15848 7300 15858 7340
rect 15898 7300 15908 7340
rect 15848 7280 15908 7300
rect 15958 7640 16098 7660
rect 15958 7600 15968 7640
rect 16008 7600 16048 7640
rect 16088 7600 16098 7640
rect 15958 7540 16098 7600
rect 15958 7500 15968 7540
rect 16008 7500 16048 7540
rect 16088 7500 16098 7540
rect 15958 7440 16098 7500
rect 15958 7400 15968 7440
rect 16008 7400 16048 7440
rect 16088 7400 16098 7440
rect 15958 7340 16098 7400
rect 15958 7300 15968 7340
rect 16008 7300 16048 7340
rect 16088 7300 16098 7340
rect 15958 7280 16098 7300
rect 16288 7640 16468 7660
rect 16288 7600 16308 7640
rect 16348 7600 16408 7640
rect 16448 7600 16468 7640
rect 16288 7540 16468 7600
rect 16288 7500 16308 7540
rect 16348 7500 16408 7540
rect 16448 7500 16468 7540
rect 16288 7440 16468 7500
rect 16288 7400 16308 7440
rect 16348 7400 16408 7440
rect 16448 7400 16468 7440
rect 16288 7340 16468 7400
rect 16288 7300 16308 7340
rect 16348 7300 16408 7340
rect 16448 7300 16468 7340
rect 16288 7280 16468 7300
rect 16518 7640 16598 7660
rect 16518 7600 16538 7640
rect 16578 7600 16598 7640
rect 16518 7540 16598 7600
rect 16518 7500 16538 7540
rect 16578 7500 16598 7540
rect 16518 7440 16598 7500
rect 16518 7400 16538 7440
rect 16578 7400 16598 7440
rect 16518 7340 16598 7400
rect 16518 7300 16538 7340
rect 16578 7300 16598 7340
rect 16518 7280 16598 7300
rect 16778 7640 16858 7660
rect 16778 7600 16798 7640
rect 16838 7600 16858 7640
rect 16778 7540 16858 7600
rect 16778 7500 16798 7540
rect 16838 7500 16858 7540
rect 16778 7440 16858 7500
rect 16778 7400 16798 7440
rect 16838 7400 16858 7440
rect 16778 7340 16858 7400
rect 16778 7300 16798 7340
rect 16838 7300 16858 7340
rect 16778 7280 16858 7300
rect 16908 7640 16988 7660
rect 16908 7600 16928 7640
rect 16968 7600 16988 7640
rect 16908 7540 16988 7600
rect 16908 7500 16928 7540
rect 16968 7500 16988 7540
rect 16908 7440 16988 7500
rect 16908 7400 16928 7440
rect 16968 7400 16988 7440
rect 16908 7340 16988 7400
rect 16908 7300 16928 7340
rect 16968 7300 16988 7340
rect 16908 7280 16988 7300
rect 17068 7640 17248 7660
rect 17068 7600 17088 7640
rect 17128 7600 17188 7640
rect 17228 7600 17248 7640
rect 17068 7540 17248 7600
rect 17068 7500 17088 7540
rect 17128 7500 17188 7540
rect 17228 7500 17248 7540
rect 17068 7440 17248 7500
rect 17068 7400 17088 7440
rect 17128 7400 17188 7440
rect 17228 7400 17248 7440
rect 17068 7340 17248 7400
rect 17068 7300 17088 7340
rect 17128 7300 17188 7340
rect 17228 7300 17248 7340
rect 17068 7280 17248 7300
rect 17298 7640 17378 7660
rect 17298 7600 17318 7640
rect 17358 7600 17378 7640
rect 17298 7540 17378 7600
rect 17298 7500 17318 7540
rect 17358 7500 17378 7540
rect 17298 7440 17378 7500
rect 17298 7400 17318 7440
rect 17358 7400 17378 7440
rect 17298 7340 17378 7400
rect 17298 7300 17318 7340
rect 17358 7300 17378 7340
rect 17298 7280 17378 7300
rect 17458 7640 17538 7660
rect 17458 7600 17478 7640
rect 17518 7600 17538 7640
rect 17458 7540 17538 7600
rect 17458 7500 17478 7540
rect 17518 7500 17538 7540
rect 17458 7440 17538 7500
rect 17458 7400 17478 7440
rect 17518 7400 17538 7440
rect 17458 7340 17538 7400
rect 17458 7300 17478 7340
rect 17518 7300 17538 7340
rect 17458 7280 17538 7300
rect 17588 7640 17668 7660
rect 19238 7650 19418 7670
rect 19558 8010 19638 8030
rect 19558 7970 19578 8010
rect 19618 7970 19638 8010
rect 19558 7910 19638 7970
rect 19558 7870 19578 7910
rect 19618 7870 19638 7910
rect 19558 7810 19638 7870
rect 19558 7770 19578 7810
rect 19618 7770 19638 7810
rect 19558 7710 19638 7770
rect 19558 7670 19578 7710
rect 19618 7670 19638 7710
rect 19558 7650 19638 7670
rect 19778 8010 19858 8030
rect 19778 7970 19798 8010
rect 19838 7970 19858 8010
rect 19778 7910 19858 7970
rect 19778 7870 19798 7910
rect 19838 7870 19858 7910
rect 19778 7810 19858 7870
rect 19778 7770 19798 7810
rect 19838 7770 19858 7810
rect 19778 7710 19858 7770
rect 19778 7670 19798 7710
rect 19838 7670 19858 7710
rect 17588 7600 17608 7640
rect 17648 7600 17668 7640
rect 17588 7540 17668 7600
rect 19778 7600 19858 7670
rect 19998 8010 20078 8030
rect 19998 7970 20018 8010
rect 20058 7970 20078 8010
rect 19998 7910 20078 7970
rect 19998 7870 20018 7910
rect 20058 7870 20078 7910
rect 19998 7810 20078 7870
rect 19998 7770 20018 7810
rect 20058 7770 20078 7810
rect 19998 7710 20078 7770
rect 19998 7670 20018 7710
rect 20058 7670 20078 7710
rect 19998 7650 20078 7670
rect 20218 8010 20498 8030
rect 20218 7970 20238 8010
rect 20278 7970 20338 8010
rect 20378 7970 20438 8010
rect 20478 7970 20498 8010
rect 20218 7910 20498 7970
rect 20218 7870 20238 7910
rect 20278 7870 20338 7910
rect 20378 7870 20438 7910
rect 20478 7870 20498 7910
rect 20218 7810 20498 7870
rect 20218 7770 20238 7810
rect 20278 7770 20338 7810
rect 20378 7770 20438 7810
rect 20478 7770 20498 7810
rect 20218 7710 20498 7770
rect 20218 7670 20238 7710
rect 20278 7670 20338 7710
rect 20378 7670 20438 7710
rect 20478 7670 20498 7710
rect 20218 7650 20498 7670
rect 20638 8010 20718 8030
rect 20638 7970 20658 8010
rect 20698 7970 20718 8010
rect 20638 7910 20718 7970
rect 20638 7870 20658 7910
rect 20698 7870 20718 7910
rect 20638 7810 20718 7870
rect 20638 7770 20658 7810
rect 20698 7770 20718 7810
rect 20638 7710 20718 7770
rect 20638 7670 20658 7710
rect 20698 7670 20718 7710
rect 20638 7650 20718 7670
rect 20858 8010 20938 8030
rect 20858 7970 20878 8010
rect 20918 7970 20938 8010
rect 20858 7910 20938 7970
rect 20858 7870 20878 7910
rect 20918 7870 20938 7910
rect 20858 7810 20938 7870
rect 20858 7770 20878 7810
rect 20918 7770 20938 7810
rect 20858 7710 20938 7770
rect 20858 7670 20878 7710
rect 20918 7670 20938 7710
rect 20858 7650 20938 7670
rect 21078 8010 21158 8030
rect 21078 7970 21098 8010
rect 21138 7970 21158 8010
rect 21078 7910 21158 7970
rect 21078 7870 21098 7910
rect 21138 7870 21158 7910
rect 21078 7810 21158 7870
rect 21078 7770 21098 7810
rect 21138 7770 21158 7810
rect 21078 7710 21158 7770
rect 21078 7670 21098 7710
rect 21138 7670 21158 7710
rect 21078 7650 21158 7670
rect 21298 8010 21578 8030
rect 21298 7970 21318 8010
rect 21358 7970 21418 8010
rect 21458 7970 21518 8010
rect 21558 7970 21578 8010
rect 21298 7910 21578 7970
rect 21298 7870 21318 7910
rect 21358 7870 21418 7910
rect 21458 7870 21518 7910
rect 21558 7870 21578 7910
rect 21298 7810 21578 7870
rect 21298 7770 21318 7810
rect 21358 7770 21418 7810
rect 21458 7770 21518 7810
rect 21558 7770 21578 7810
rect 21298 7710 21578 7770
rect 21298 7670 21318 7710
rect 21358 7670 21418 7710
rect 21458 7670 21518 7710
rect 21558 7670 21578 7710
rect 21298 7650 21578 7670
rect 21718 8010 21798 8030
rect 21718 7970 21738 8010
rect 21778 7970 21798 8010
rect 21718 7910 21798 7970
rect 21718 7870 21738 7910
rect 21778 7870 21798 7910
rect 21718 7810 21798 7870
rect 21718 7770 21738 7810
rect 21778 7770 21798 7810
rect 21718 7710 21798 7770
rect 21718 7670 21738 7710
rect 21778 7670 21798 7710
rect 21718 7650 21798 7670
rect 21938 8010 22018 8030
rect 21938 7970 21958 8010
rect 21998 7970 22018 8010
rect 21938 7910 22018 7970
rect 21938 7870 21958 7910
rect 21998 7870 22018 7910
rect 21938 7810 22018 7870
rect 21938 7770 21958 7810
rect 21998 7770 22018 7810
rect 21938 7710 22018 7770
rect 21938 7670 21958 7710
rect 21998 7670 22018 7710
rect 21938 7650 22018 7670
rect 22158 8010 22238 8030
rect 22158 7970 22178 8010
rect 22218 7970 22238 8010
rect 22158 7910 22238 7970
rect 22158 7870 22178 7910
rect 22218 7870 22238 7910
rect 22158 7810 22238 7870
rect 22158 7770 22178 7810
rect 22218 7770 22238 7810
rect 22158 7710 22238 7770
rect 22158 7670 22178 7710
rect 22218 7670 22238 7710
rect 22158 7650 22238 7670
rect 22378 8010 22558 8030
rect 22378 7970 22398 8010
rect 22438 7970 22498 8010
rect 22538 7970 22558 8010
rect 22378 7910 22558 7970
rect 22378 7870 22398 7910
rect 22438 7870 22498 7910
rect 22538 7870 22558 7910
rect 22378 7810 22558 7870
rect 22378 7770 22398 7810
rect 22438 7770 22498 7810
rect 22538 7770 22558 7810
rect 22378 7710 22558 7770
rect 22378 7670 22398 7710
rect 22438 7670 22498 7710
rect 22538 7670 22558 7710
rect 22378 7650 22558 7670
rect 19778 7560 19798 7600
rect 19838 7560 19858 7600
rect 19778 7540 19858 7560
rect 20318 7590 20398 7650
rect 20318 7550 20338 7590
rect 20378 7550 20398 7590
rect 17588 7500 17608 7540
rect 17648 7500 17668 7540
rect 20318 7530 20398 7550
rect 21398 7590 21478 7650
rect 21398 7550 21418 7590
rect 21458 7550 21478 7590
rect 22738 7590 22848 7610
rect 21398 7530 21478 7550
rect 21808 7560 21888 7580
rect 21808 7520 21828 7560
rect 21868 7520 21888 7560
rect 21808 7500 21888 7520
rect 22068 7560 22148 7580
rect 22068 7520 22088 7560
rect 22128 7520 22148 7560
rect 22068 7500 22148 7520
rect 22738 7520 22758 7590
rect 22828 7520 22848 7590
rect 22738 7500 22848 7520
rect 17588 7440 17668 7500
rect 17588 7400 17608 7440
rect 17648 7400 17668 7440
rect 17588 7340 17668 7400
rect 17588 7300 17608 7340
rect 17648 7300 17668 7340
rect 17588 7280 17668 7300
rect 13268 7130 13308 7280
rect 13698 7240 13738 7280
rect 13698 7220 13778 7240
rect 13698 7180 13718 7220
rect 13758 7180 13778 7220
rect 13698 7160 13778 7180
rect 14008 7130 14048 7280
rect 14168 7130 14208 7280
rect 14908 7130 14948 7280
rect 15328 7130 15368 7280
rect 15638 7130 15678 7280
rect 15968 7130 16008 7280
rect 16408 7130 16448 7280
rect 16818 7220 16898 7240
rect 16818 7180 16838 7220
rect 16878 7180 16898 7220
rect 16818 7170 16898 7180
rect 17188 7130 17228 7280
rect 17478 7240 17518 7280
rect 17458 7220 17538 7240
rect 17458 7180 17478 7220
rect 17518 7180 17538 7220
rect 17458 7160 17538 7180
rect 13248 7110 13328 7130
rect 13248 7070 13268 7110
rect 13308 7070 13328 7110
rect 13248 7050 13328 7070
rect 13988 7110 14068 7130
rect 13988 7070 14008 7110
rect 14048 7070 14068 7110
rect 13988 7050 14068 7070
rect 14148 7110 14228 7130
rect 14148 7070 14168 7110
rect 14208 7070 14228 7110
rect 14148 7050 14228 7070
rect 14888 7110 14968 7130
rect 14888 7070 14908 7110
rect 14948 7070 14968 7110
rect 14888 7050 14968 7070
rect 15138 7110 15218 7130
rect 15138 7070 15158 7110
rect 15198 7070 15218 7110
rect 15138 7050 15218 7070
rect 15328 7110 15488 7130
rect 15328 7070 15348 7110
rect 15388 7070 15428 7110
rect 15468 7070 15488 7110
rect 15328 7050 15488 7070
rect 15618 7110 15698 7130
rect 15618 7070 15638 7110
rect 15678 7070 15698 7110
rect 15618 7050 15698 7070
rect 15948 7110 16028 7130
rect 15948 7070 15968 7110
rect 16008 7070 16028 7110
rect 15948 7050 16028 7070
rect 16388 7110 16468 7130
rect 16388 7070 16408 7110
rect 16448 7070 16468 7110
rect 16388 7050 16468 7070
rect 16778 7110 16858 7130
rect 16778 7070 16798 7110
rect 16838 7070 16858 7110
rect 16778 7050 16858 7070
rect 17168 7110 17248 7130
rect 17168 7070 17188 7110
rect 17228 7070 17248 7110
rect 17168 7050 17248 7070
rect 17848 7110 17928 7130
rect 17848 7070 17868 7110
rect 17908 7070 17928 7110
rect 17848 7050 17928 7070
rect 21368 7060 21448 7080
rect 13268 6900 13308 7050
rect 14008 6900 14048 7050
rect 14168 6900 14208 7050
rect 14908 6900 14948 7050
rect 15168 6900 15208 7050
rect 15248 7000 15328 7010
rect 15248 6960 15268 7000
rect 15308 6960 15328 7000
rect 15248 6940 15328 6960
rect 15428 6900 15468 7050
rect 15648 6900 15688 7050
rect 15978 6900 16018 7050
rect 16408 6900 16448 7050
rect 16798 6900 16838 7050
rect 17188 6900 17228 7050
rect 17868 6900 17908 7050
rect 20198 7030 20278 7050
rect 20198 6990 20218 7030
rect 20258 6990 20278 7030
rect 20198 6970 20278 6990
rect 20958 7030 21038 7050
rect 20958 6990 20978 7030
rect 21018 6990 21038 7030
rect 21368 7020 21388 7060
rect 21428 7020 21448 7060
rect 21368 7000 21448 7020
rect 22068 7060 22148 7080
rect 22068 7020 22088 7060
rect 22128 7020 22148 7060
rect 22068 7000 22148 7020
rect 22738 7060 22848 7080
rect 20958 6930 21038 6990
rect 22738 6990 22758 7060
rect 22828 6990 22848 7060
rect 22738 6970 22848 6990
rect 19438 6910 19618 6930
rect 13178 6880 13318 6900
rect 13178 6840 13188 6880
rect 13228 6840 13268 6880
rect 13308 6840 13318 6880
rect 13178 6780 13318 6840
rect 13178 6740 13188 6780
rect 13228 6740 13268 6780
rect 13308 6740 13318 6780
rect 13178 6680 13318 6740
rect 13178 6640 13188 6680
rect 13228 6640 13268 6680
rect 13308 6640 13318 6680
rect 13178 6580 13318 6640
rect 13178 6540 13188 6580
rect 13228 6540 13268 6580
rect 13308 6540 13318 6580
rect 13178 6520 13318 6540
rect 13368 6880 13428 6900
rect 13368 6840 13378 6880
rect 13418 6840 13428 6880
rect 13368 6780 13428 6840
rect 13368 6740 13378 6780
rect 13418 6740 13428 6780
rect 13368 6680 13428 6740
rect 13368 6640 13378 6680
rect 13418 6640 13428 6680
rect 13368 6580 13428 6640
rect 13368 6540 13378 6580
rect 13418 6540 13428 6580
rect 13368 6520 13428 6540
rect 13478 6880 13658 6900
rect 13478 6840 13488 6880
rect 13528 6850 13598 6880
rect 13528 6840 13538 6850
rect 13478 6780 13538 6840
rect 13578 6840 13598 6850
rect 13638 6840 13658 6880
rect 13578 6820 13658 6840
rect 13698 6880 13838 6900
rect 13698 6860 13788 6880
rect 13478 6740 13488 6780
rect 13528 6740 13538 6780
rect 13478 6680 13538 6740
rect 13478 6640 13488 6680
rect 13528 6640 13538 6680
rect 13478 6580 13538 6640
rect 13478 6540 13488 6580
rect 13528 6540 13538 6580
rect 13478 6520 13538 6540
rect 13488 6480 13528 6520
rect 13368 6440 13528 6480
rect 13128 6420 13208 6440
rect 13128 6380 13148 6420
rect 13188 6380 13208 6420
rect 13128 6360 13208 6380
rect 13368 6280 13408 6440
rect 13698 6400 13738 6860
rect 13778 6840 13788 6860
rect 13828 6840 13838 6880
rect 13778 6780 13838 6840
rect 13778 6740 13788 6780
rect 13828 6740 13838 6780
rect 13778 6680 13838 6740
rect 13778 6640 13788 6680
rect 13828 6640 13838 6680
rect 13778 6580 13838 6640
rect 13778 6540 13788 6580
rect 13828 6540 13838 6580
rect 13778 6520 13838 6540
rect 13888 6880 13948 6900
rect 13888 6840 13898 6880
rect 13938 6840 13948 6880
rect 13888 6780 13948 6840
rect 13888 6740 13898 6780
rect 13938 6740 13948 6780
rect 13888 6680 13948 6740
rect 13888 6640 13898 6680
rect 13938 6640 13948 6680
rect 13888 6580 13948 6640
rect 13888 6540 13898 6580
rect 13938 6540 13948 6580
rect 13888 6520 13948 6540
rect 13998 6880 14218 6900
rect 13998 6840 14008 6880
rect 14048 6840 14088 6880
rect 14128 6840 14168 6880
rect 14208 6840 14218 6880
rect 13998 6780 14218 6840
rect 13998 6740 14008 6780
rect 14048 6740 14088 6780
rect 14128 6740 14168 6780
rect 14208 6740 14218 6780
rect 13998 6680 14218 6740
rect 13998 6640 14008 6680
rect 14048 6640 14088 6680
rect 14128 6640 14168 6680
rect 14208 6640 14218 6680
rect 13998 6580 14218 6640
rect 13998 6540 14008 6580
rect 14048 6540 14088 6580
rect 14128 6540 14168 6580
rect 14208 6540 14218 6580
rect 13998 6520 14218 6540
rect 14268 6880 14328 6900
rect 14268 6840 14278 6880
rect 14318 6840 14328 6880
rect 14268 6780 14328 6840
rect 14268 6740 14278 6780
rect 14318 6740 14328 6780
rect 14268 6680 14328 6740
rect 14268 6640 14278 6680
rect 14318 6640 14328 6680
rect 14268 6580 14328 6640
rect 14268 6540 14278 6580
rect 14318 6540 14328 6580
rect 14268 6520 14328 6540
rect 14378 6880 14558 6900
rect 14378 6840 14388 6880
rect 14428 6850 14498 6880
rect 14428 6840 14438 6850
rect 14378 6780 14438 6840
rect 14478 6840 14498 6850
rect 14538 6840 14558 6880
rect 14478 6820 14558 6840
rect 14598 6880 14738 6900
rect 14598 6860 14688 6880
rect 14378 6740 14388 6780
rect 14428 6740 14438 6780
rect 14378 6680 14438 6740
rect 14378 6640 14388 6680
rect 14428 6640 14438 6680
rect 14378 6580 14438 6640
rect 14378 6540 14388 6580
rect 14428 6540 14438 6580
rect 14378 6520 14438 6540
rect 13788 6480 13828 6520
rect 14388 6480 14428 6520
rect 13788 6440 13938 6480
rect 13458 6380 13738 6400
rect 13458 6340 13478 6380
rect 13518 6360 13738 6380
rect 13518 6340 13538 6360
rect 13458 6320 13538 6340
rect 13178 6260 13318 6280
rect 13178 6220 13188 6260
rect 13228 6220 13268 6260
rect 13308 6220 13318 6260
rect 13178 6160 13318 6220
rect 13178 6120 13188 6160
rect 13228 6120 13268 6160
rect 13308 6120 13318 6160
rect 13178 6100 13318 6120
rect 13368 6260 13428 6280
rect 13368 6220 13378 6260
rect 13418 6220 13428 6260
rect 13368 6160 13428 6220
rect 13368 6120 13378 6160
rect 13418 6120 13428 6160
rect 13368 6100 13428 6120
rect 13478 6260 13538 6280
rect 13478 6220 13488 6260
rect 13528 6220 13538 6260
rect 13478 6160 13538 6220
rect 13478 6120 13488 6160
rect 13528 6120 13538 6160
rect 13478 6100 13538 6120
rect 13268 5950 13308 6100
rect 13488 5950 13528 6100
rect 13698 6060 13738 6360
rect 13898 6280 13938 6440
rect 13978 6460 14428 6480
rect 13978 6420 13998 6460
rect 14038 6440 14428 6460
rect 14038 6420 14058 6440
rect 13978 6400 14058 6420
rect 14268 6280 14308 6440
rect 14598 6400 14638 6860
rect 14678 6840 14688 6860
rect 14728 6840 14738 6880
rect 14678 6780 14738 6840
rect 14678 6740 14688 6780
rect 14728 6740 14738 6780
rect 14678 6680 14738 6740
rect 14678 6640 14688 6680
rect 14728 6640 14738 6680
rect 14678 6580 14738 6640
rect 14678 6540 14688 6580
rect 14728 6540 14738 6580
rect 14678 6520 14738 6540
rect 14788 6880 14848 6900
rect 14788 6840 14798 6880
rect 14838 6840 14848 6880
rect 14788 6780 14848 6840
rect 14788 6740 14798 6780
rect 14838 6740 14848 6780
rect 14788 6680 14848 6740
rect 14788 6640 14798 6680
rect 14838 6640 14848 6680
rect 14788 6580 14848 6640
rect 14788 6540 14798 6580
rect 14838 6540 14848 6580
rect 14788 6520 14848 6540
rect 14898 6880 15038 6900
rect 14898 6840 14908 6880
rect 14948 6840 14988 6880
rect 15028 6840 15038 6880
rect 14898 6780 15038 6840
rect 14898 6740 14908 6780
rect 14948 6740 14988 6780
rect 15028 6740 15038 6780
rect 14898 6680 15038 6740
rect 14898 6640 14908 6680
rect 14948 6640 14988 6680
rect 15028 6640 15038 6680
rect 14898 6580 15038 6640
rect 14898 6540 14908 6580
rect 14948 6540 14988 6580
rect 15028 6540 15038 6580
rect 14898 6520 15038 6540
rect 15118 6880 15258 6900
rect 15118 6840 15128 6880
rect 15168 6840 15208 6880
rect 15248 6840 15258 6880
rect 15118 6780 15258 6840
rect 15118 6740 15128 6780
rect 15168 6740 15208 6780
rect 15248 6740 15258 6780
rect 15118 6680 15258 6740
rect 15118 6640 15128 6680
rect 15168 6640 15208 6680
rect 15248 6640 15258 6680
rect 15118 6580 15258 6640
rect 15118 6540 15128 6580
rect 15168 6540 15208 6580
rect 15248 6540 15258 6580
rect 15118 6520 15258 6540
rect 15308 6880 15368 6900
rect 15308 6840 15318 6880
rect 15358 6840 15368 6880
rect 15308 6780 15368 6840
rect 15308 6740 15318 6780
rect 15358 6740 15368 6780
rect 15308 6680 15368 6740
rect 15308 6640 15318 6680
rect 15358 6640 15368 6680
rect 15308 6580 15368 6640
rect 15308 6540 15318 6580
rect 15358 6540 15368 6580
rect 15308 6520 15368 6540
rect 15418 6880 15478 6900
rect 15418 6840 15428 6880
rect 15468 6840 15478 6880
rect 15418 6780 15478 6840
rect 15418 6740 15428 6780
rect 15468 6740 15478 6780
rect 15418 6680 15478 6740
rect 15418 6640 15428 6680
rect 15468 6640 15478 6680
rect 15418 6580 15478 6640
rect 15418 6540 15428 6580
rect 15468 6540 15478 6580
rect 15418 6520 15478 6540
rect 15558 6880 15698 6900
rect 15558 6840 15568 6880
rect 15608 6840 15648 6880
rect 15688 6840 15698 6880
rect 15558 6780 15698 6840
rect 15558 6740 15568 6780
rect 15608 6740 15648 6780
rect 15688 6740 15698 6780
rect 15558 6680 15698 6740
rect 15558 6640 15568 6680
rect 15608 6640 15648 6680
rect 15688 6640 15698 6680
rect 15558 6580 15698 6640
rect 15558 6540 15568 6580
rect 15608 6540 15648 6580
rect 15688 6540 15698 6580
rect 15558 6520 15698 6540
rect 15748 6880 15808 6900
rect 15748 6840 15758 6880
rect 15798 6840 15808 6880
rect 15748 6780 15808 6840
rect 15748 6740 15758 6780
rect 15798 6740 15808 6780
rect 15748 6680 15808 6740
rect 15748 6640 15758 6680
rect 15798 6640 15808 6680
rect 15748 6580 15808 6640
rect 15748 6540 15758 6580
rect 15798 6540 15808 6580
rect 15748 6520 15808 6540
rect 15888 6880 16028 6900
rect 15888 6840 15898 6880
rect 15938 6840 15978 6880
rect 16018 6840 16028 6880
rect 15888 6780 16028 6840
rect 15888 6740 15898 6780
rect 15938 6740 15978 6780
rect 16018 6740 16028 6780
rect 15888 6680 16028 6740
rect 15888 6640 15898 6680
rect 15938 6640 15978 6680
rect 16018 6640 16028 6680
rect 15888 6580 16028 6640
rect 15888 6540 15898 6580
rect 15938 6540 15978 6580
rect 16018 6540 16028 6580
rect 15888 6520 16028 6540
rect 16078 6880 16138 6900
rect 16078 6840 16088 6880
rect 16128 6840 16138 6880
rect 16078 6780 16138 6840
rect 16078 6740 16088 6780
rect 16128 6740 16138 6780
rect 16078 6680 16138 6740
rect 16078 6640 16088 6680
rect 16128 6640 16138 6680
rect 16078 6580 16138 6640
rect 16078 6540 16088 6580
rect 16128 6540 16138 6580
rect 16078 6520 16138 6540
rect 16288 6880 16468 6900
rect 16288 6840 16308 6880
rect 16348 6840 16408 6880
rect 16448 6840 16468 6880
rect 16288 6780 16468 6840
rect 16288 6740 16308 6780
rect 16348 6740 16408 6780
rect 16448 6740 16468 6780
rect 16288 6680 16468 6740
rect 16288 6640 16308 6680
rect 16348 6640 16408 6680
rect 16448 6640 16468 6680
rect 16288 6580 16468 6640
rect 16288 6540 16308 6580
rect 16348 6540 16408 6580
rect 16448 6540 16468 6580
rect 16288 6520 16468 6540
rect 16518 6880 16598 6900
rect 16518 6840 16538 6880
rect 16578 6840 16598 6880
rect 16518 6780 16598 6840
rect 16518 6740 16538 6780
rect 16578 6740 16598 6780
rect 16518 6680 16598 6740
rect 16518 6640 16538 6680
rect 16578 6640 16598 6680
rect 16518 6580 16598 6640
rect 16518 6540 16538 6580
rect 16578 6540 16598 6580
rect 16518 6520 16598 6540
rect 16678 6880 16858 6900
rect 16678 6840 16698 6880
rect 16738 6840 16798 6880
rect 16838 6840 16858 6880
rect 16678 6780 16858 6840
rect 16678 6740 16698 6780
rect 16738 6740 16798 6780
rect 16838 6740 16858 6780
rect 16678 6680 16858 6740
rect 16678 6640 16698 6680
rect 16738 6640 16798 6680
rect 16838 6640 16858 6680
rect 16678 6580 16858 6640
rect 16678 6540 16698 6580
rect 16738 6540 16798 6580
rect 16838 6540 16858 6580
rect 16678 6520 16858 6540
rect 16908 6880 16988 6900
rect 16908 6840 16928 6880
rect 16968 6840 16988 6880
rect 16908 6780 16988 6840
rect 16908 6740 16928 6780
rect 16968 6740 16988 6780
rect 16908 6680 16988 6740
rect 16908 6640 16928 6680
rect 16968 6640 16988 6680
rect 16908 6580 16988 6640
rect 16908 6540 16928 6580
rect 16968 6540 16988 6580
rect 16908 6520 16988 6540
rect 17068 6880 17248 6900
rect 17068 6840 17088 6880
rect 17128 6840 17188 6880
rect 17228 6840 17248 6880
rect 17068 6780 17248 6840
rect 17068 6740 17088 6780
rect 17128 6740 17188 6780
rect 17228 6740 17248 6780
rect 17068 6680 17248 6740
rect 17068 6640 17088 6680
rect 17128 6640 17188 6680
rect 17228 6640 17248 6680
rect 17068 6580 17248 6640
rect 17068 6540 17088 6580
rect 17128 6540 17188 6580
rect 17228 6540 17248 6580
rect 17068 6520 17248 6540
rect 17298 6880 17378 6900
rect 17298 6840 17318 6880
rect 17358 6840 17378 6880
rect 17298 6780 17378 6840
rect 17298 6740 17318 6780
rect 17358 6740 17378 6780
rect 17298 6680 17378 6740
rect 17298 6640 17318 6680
rect 17358 6640 17378 6680
rect 17298 6580 17378 6640
rect 17298 6540 17318 6580
rect 17358 6540 17378 6580
rect 17298 6520 17378 6540
rect 17458 6880 17538 6900
rect 17458 6840 17478 6880
rect 17518 6840 17538 6880
rect 17458 6780 17538 6840
rect 17458 6740 17478 6780
rect 17518 6740 17538 6780
rect 17458 6680 17538 6740
rect 17458 6640 17478 6680
rect 17518 6640 17538 6680
rect 17458 6580 17538 6640
rect 17458 6540 17478 6580
rect 17518 6540 17538 6580
rect 17458 6520 17538 6540
rect 17588 6880 17668 6900
rect 17588 6840 17608 6880
rect 17648 6840 17668 6880
rect 17588 6780 17668 6840
rect 17588 6740 17608 6780
rect 17648 6740 17668 6780
rect 17588 6680 17668 6740
rect 17588 6640 17608 6680
rect 17648 6640 17668 6680
rect 17588 6580 17668 6640
rect 17588 6540 17608 6580
rect 17648 6540 17668 6580
rect 17588 6520 17668 6540
rect 17748 6880 17928 6900
rect 17748 6840 17768 6880
rect 17808 6840 17868 6880
rect 17908 6840 17928 6880
rect 17748 6780 17928 6840
rect 17748 6740 17768 6780
rect 17808 6740 17868 6780
rect 17908 6740 17928 6780
rect 17748 6680 17928 6740
rect 17748 6640 17768 6680
rect 17808 6640 17868 6680
rect 17908 6640 17928 6680
rect 17748 6580 17928 6640
rect 17748 6540 17768 6580
rect 17808 6540 17868 6580
rect 17908 6540 17928 6580
rect 17748 6520 17928 6540
rect 17978 6880 18058 6900
rect 17978 6840 17998 6880
rect 18038 6840 18058 6880
rect 17978 6780 18058 6840
rect 17978 6740 17998 6780
rect 18038 6740 18058 6780
rect 17978 6680 18058 6740
rect 17978 6640 17998 6680
rect 18038 6640 18058 6680
rect 17978 6580 18058 6640
rect 17978 6540 17998 6580
rect 18038 6540 18058 6580
rect 19438 6870 19458 6910
rect 19498 6870 19558 6910
rect 19598 6870 19618 6910
rect 19438 6810 19618 6870
rect 19438 6770 19458 6810
rect 19498 6770 19558 6810
rect 19598 6770 19618 6810
rect 19438 6710 19618 6770
rect 19438 6670 19458 6710
rect 19498 6670 19558 6710
rect 19598 6670 19618 6710
rect 19438 6610 19618 6670
rect 19438 6570 19458 6610
rect 19498 6570 19558 6610
rect 19598 6570 19618 6610
rect 19438 6550 19618 6570
rect 19758 6910 19838 6930
rect 19758 6870 19778 6910
rect 19818 6870 19838 6910
rect 19758 6810 19838 6870
rect 19758 6770 19778 6810
rect 19818 6770 19838 6810
rect 19758 6710 19838 6770
rect 19758 6670 19778 6710
rect 19818 6670 19838 6710
rect 19758 6610 19838 6670
rect 19758 6570 19778 6610
rect 19818 6570 19838 6610
rect 19758 6550 19838 6570
rect 19978 6910 20058 6930
rect 19978 6870 19998 6910
rect 20038 6870 20058 6910
rect 19978 6810 20058 6870
rect 19978 6770 19998 6810
rect 20038 6770 20058 6810
rect 19978 6710 20058 6770
rect 19978 6670 19998 6710
rect 20038 6670 20058 6710
rect 19978 6610 20058 6670
rect 19978 6570 19998 6610
rect 20038 6570 20058 6610
rect 19978 6550 20058 6570
rect 20198 6910 20278 6930
rect 20198 6870 20218 6910
rect 20258 6870 20278 6910
rect 20198 6810 20278 6870
rect 20198 6770 20218 6810
rect 20258 6770 20278 6810
rect 20198 6710 20278 6770
rect 20198 6670 20218 6710
rect 20258 6670 20278 6710
rect 20198 6610 20278 6670
rect 20198 6570 20218 6610
rect 20258 6570 20278 6610
rect 20198 6550 20278 6570
rect 20418 6910 20498 6930
rect 20418 6870 20438 6910
rect 20478 6870 20498 6910
rect 20418 6810 20498 6870
rect 20418 6770 20438 6810
rect 20478 6770 20498 6810
rect 20418 6710 20498 6770
rect 20418 6670 20438 6710
rect 20478 6670 20498 6710
rect 20418 6610 20498 6670
rect 20418 6570 20438 6610
rect 20478 6570 20498 6610
rect 20418 6550 20498 6570
rect 20638 6910 20718 6930
rect 20638 6870 20658 6910
rect 20698 6870 20718 6910
rect 20638 6810 20718 6870
rect 20638 6770 20658 6810
rect 20698 6770 20718 6810
rect 20638 6710 20718 6770
rect 20638 6670 20658 6710
rect 20698 6670 20718 6710
rect 20638 6610 20718 6670
rect 20638 6570 20658 6610
rect 20698 6570 20718 6610
rect 20638 6550 20718 6570
rect 20858 6910 21138 6930
rect 20858 6870 20878 6910
rect 20918 6870 20978 6910
rect 21018 6870 21078 6910
rect 21118 6870 21138 6910
rect 20858 6810 21138 6870
rect 20858 6770 20878 6810
rect 20918 6770 20978 6810
rect 21018 6770 21078 6810
rect 21118 6770 21138 6810
rect 20858 6710 21138 6770
rect 20858 6670 20878 6710
rect 20918 6670 20978 6710
rect 21018 6670 21078 6710
rect 21118 6670 21138 6710
rect 20858 6610 21138 6670
rect 20858 6570 20878 6610
rect 20918 6570 20978 6610
rect 21018 6570 21078 6610
rect 21118 6570 21138 6610
rect 20858 6550 21138 6570
rect 21278 6910 21358 6930
rect 21278 6870 21298 6910
rect 21338 6870 21358 6910
rect 21278 6810 21358 6870
rect 21278 6770 21298 6810
rect 21338 6770 21358 6810
rect 21278 6710 21358 6770
rect 21278 6670 21298 6710
rect 21338 6670 21358 6710
rect 21278 6610 21358 6670
rect 21278 6570 21298 6610
rect 21338 6570 21358 6610
rect 21278 6550 21358 6570
rect 21498 6910 21578 6930
rect 21498 6870 21518 6910
rect 21558 6870 21578 6910
rect 21498 6810 21578 6870
rect 21498 6770 21518 6810
rect 21558 6770 21578 6810
rect 21498 6710 21578 6770
rect 21498 6670 21518 6710
rect 21558 6670 21578 6710
rect 21498 6610 21578 6670
rect 21498 6570 21518 6610
rect 21558 6570 21578 6610
rect 21498 6550 21578 6570
rect 21718 6910 21798 6930
rect 21718 6870 21738 6910
rect 21778 6870 21798 6910
rect 21718 6810 21798 6870
rect 21718 6770 21738 6810
rect 21778 6770 21798 6810
rect 21718 6710 21798 6770
rect 21718 6670 21738 6710
rect 21778 6670 21798 6710
rect 21718 6610 21798 6670
rect 21718 6570 21738 6610
rect 21778 6570 21798 6610
rect 21718 6550 21798 6570
rect 21938 6910 22018 6930
rect 21938 6870 21958 6910
rect 21998 6870 22018 6910
rect 21938 6810 22018 6870
rect 21938 6770 21958 6810
rect 21998 6770 22018 6810
rect 21938 6710 22018 6770
rect 21938 6670 21958 6710
rect 21998 6670 22018 6710
rect 21938 6610 22018 6670
rect 21938 6570 21958 6610
rect 21998 6570 22018 6610
rect 21938 6550 22018 6570
rect 22158 6910 22238 6930
rect 22158 6870 22178 6910
rect 22218 6870 22238 6910
rect 22158 6810 22238 6870
rect 22158 6770 22178 6810
rect 22218 6770 22238 6810
rect 22158 6710 22238 6770
rect 22158 6670 22178 6710
rect 22218 6670 22238 6710
rect 22158 6610 22238 6670
rect 22158 6570 22178 6610
rect 22218 6570 22238 6610
rect 22158 6550 22238 6570
rect 22378 6910 22558 6930
rect 22378 6870 22398 6910
rect 22438 6870 22498 6910
rect 22538 6870 22558 6910
rect 22378 6810 22558 6870
rect 22378 6770 22398 6810
rect 22438 6770 22498 6810
rect 22538 6770 22558 6810
rect 22378 6710 22558 6770
rect 22378 6670 22398 6710
rect 22438 6670 22498 6710
rect 22538 6670 22558 6710
rect 22378 6610 22558 6670
rect 22378 6570 22398 6610
rect 22438 6570 22498 6610
rect 22538 6570 22558 6610
rect 22378 6550 22558 6570
rect 17978 6520 18058 6540
rect 14688 6480 14728 6520
rect 14688 6440 14838 6480
rect 14358 6380 14638 6400
rect 14358 6340 14378 6380
rect 14418 6360 14638 6380
rect 14418 6340 14438 6360
rect 14358 6320 14438 6340
rect 14798 6280 14838 6440
rect 15318 6450 15358 6520
rect 15768 6450 15808 6520
rect 16098 6450 16138 6520
rect 15318 6430 15538 6450
rect 15318 6410 15478 6430
rect 15028 6390 15108 6410
rect 15028 6350 15048 6390
rect 15088 6350 15108 6390
rect 15028 6330 15108 6350
rect 15428 6390 15478 6410
rect 15518 6390 15538 6430
rect 15428 6370 15538 6390
rect 15768 6430 15868 6450
rect 15768 6390 15808 6430
rect 15848 6390 15868 6430
rect 15768 6370 15868 6390
rect 16098 6430 16198 6450
rect 16098 6390 16138 6430
rect 16178 6390 16198 6430
rect 16558 6430 16598 6520
rect 16818 6430 16898 6450
rect 16098 6370 16198 6390
rect 16248 6400 16328 6420
rect 15428 6280 15468 6370
rect 15768 6280 15808 6370
rect 16098 6280 16138 6370
rect 16248 6360 16268 6400
rect 16308 6360 16328 6400
rect 16248 6340 16328 6360
rect 16558 6390 16838 6430
rect 16878 6390 16898 6430
rect 16558 6280 16598 6390
rect 16818 6370 16898 6390
rect 16948 6400 16988 6520
rect 17338 6480 17378 6520
rect 17338 6460 17418 6480
rect 17338 6420 17358 6460
rect 17398 6420 17418 6460
rect 17338 6400 17418 6420
rect 16948 6380 17288 6400
rect 16948 6360 17228 6380
rect 16948 6280 16988 6360
rect 17208 6340 17228 6360
rect 17268 6340 17288 6380
rect 17208 6320 17288 6340
rect 17338 6280 17378 6400
rect 17478 6280 17518 6520
rect 17608 6360 17648 6520
rect 17688 6460 17768 6480
rect 17688 6420 17708 6460
rect 17748 6420 17768 6460
rect 17688 6400 17768 6420
rect 17998 6400 18038 6520
rect 19538 6490 19618 6510
rect 19538 6450 19558 6490
rect 19598 6450 19618 6490
rect 19538 6430 19618 6450
rect 22378 6490 22458 6510
rect 22378 6450 22398 6490
rect 22438 6450 22458 6490
rect 22378 6430 22458 6450
rect 17998 6380 18078 6400
rect 17998 6360 18018 6380
rect 17608 6340 18018 6360
rect 18058 6340 18078 6380
rect 17608 6320 18078 6340
rect 17608 6280 17648 6320
rect 13778 6260 13838 6280
rect 13778 6220 13788 6260
rect 13828 6220 13838 6260
rect 13778 6160 13838 6220
rect 13778 6120 13788 6160
rect 13828 6120 13838 6160
rect 13778 6100 13838 6120
rect 13888 6260 13948 6280
rect 13888 6220 13898 6260
rect 13938 6220 13948 6260
rect 13888 6160 13948 6220
rect 13888 6120 13898 6160
rect 13938 6120 13948 6160
rect 13888 6100 13948 6120
rect 13998 6260 14218 6280
rect 13998 6220 14008 6260
rect 14048 6220 14088 6260
rect 14128 6220 14168 6260
rect 14208 6220 14218 6260
rect 13998 6160 14218 6220
rect 13998 6120 14008 6160
rect 14048 6120 14088 6160
rect 14128 6120 14168 6160
rect 14208 6120 14218 6160
rect 13998 6100 14218 6120
rect 14268 6260 14328 6280
rect 14268 6220 14278 6260
rect 14318 6220 14328 6260
rect 14268 6160 14328 6220
rect 14268 6120 14278 6160
rect 14318 6120 14328 6160
rect 14268 6100 14328 6120
rect 14378 6260 14438 6280
rect 14378 6220 14388 6260
rect 14428 6220 14438 6260
rect 14378 6160 14438 6220
rect 14378 6120 14388 6160
rect 14428 6120 14438 6160
rect 14378 6100 14438 6120
rect 14678 6260 14738 6280
rect 14678 6220 14688 6260
rect 14728 6220 14738 6260
rect 14678 6160 14738 6220
rect 14678 6120 14688 6160
rect 14728 6120 14738 6160
rect 14678 6100 14738 6120
rect 14788 6260 14848 6280
rect 14788 6220 14798 6260
rect 14838 6220 14848 6260
rect 14788 6160 14848 6220
rect 14788 6120 14798 6160
rect 14838 6120 14848 6160
rect 14788 6100 14848 6120
rect 14898 6260 15038 6280
rect 14898 6220 14908 6260
rect 14948 6220 14988 6260
rect 15028 6220 15038 6260
rect 14898 6160 15038 6220
rect 14898 6120 14908 6160
rect 14948 6120 14988 6160
rect 15028 6120 15038 6160
rect 14898 6100 15038 6120
rect 15118 6260 15258 6280
rect 15118 6220 15128 6260
rect 15168 6220 15208 6260
rect 15248 6220 15258 6260
rect 15118 6160 15258 6220
rect 15118 6120 15128 6160
rect 15168 6120 15208 6160
rect 15248 6120 15258 6160
rect 15118 6100 15258 6120
rect 15308 6260 15368 6280
rect 15308 6220 15318 6260
rect 15358 6220 15368 6260
rect 15308 6160 15368 6220
rect 15308 6120 15318 6160
rect 15358 6120 15368 6160
rect 15308 6100 15368 6120
rect 15418 6260 15478 6280
rect 15418 6220 15428 6260
rect 15468 6220 15478 6260
rect 15418 6160 15478 6220
rect 15418 6120 15428 6160
rect 15468 6120 15478 6160
rect 15418 6100 15478 6120
rect 15558 6260 15698 6280
rect 15558 6220 15568 6260
rect 15608 6220 15648 6260
rect 15688 6220 15698 6260
rect 15558 6160 15698 6220
rect 15558 6120 15568 6160
rect 15608 6120 15648 6160
rect 15688 6120 15698 6160
rect 15558 6100 15698 6120
rect 15748 6260 15808 6280
rect 15748 6220 15758 6260
rect 15798 6220 15808 6260
rect 15748 6160 15808 6220
rect 15748 6120 15758 6160
rect 15798 6120 15808 6160
rect 15748 6100 15808 6120
rect 15888 6260 16028 6280
rect 15888 6220 15898 6260
rect 15938 6220 15978 6260
rect 16018 6220 16028 6260
rect 15888 6160 16028 6220
rect 15888 6120 15898 6160
rect 15938 6120 15978 6160
rect 16018 6120 16028 6160
rect 15888 6100 16028 6120
rect 16078 6260 16138 6280
rect 16078 6220 16088 6260
rect 16128 6220 16138 6260
rect 16078 6160 16138 6220
rect 16078 6120 16088 6160
rect 16128 6120 16138 6160
rect 16078 6100 16138 6120
rect 16308 6260 16468 6280
rect 16308 6220 16318 6260
rect 16358 6220 16408 6260
rect 16448 6220 16468 6260
rect 16308 6160 16468 6220
rect 16308 6120 16318 6160
rect 16358 6120 16408 6160
rect 16448 6120 16468 6160
rect 16308 6100 16468 6120
rect 16518 6260 16598 6280
rect 16518 6220 16538 6260
rect 16578 6220 16598 6260
rect 16518 6160 16598 6220
rect 16518 6120 16538 6160
rect 16578 6120 16598 6160
rect 16518 6100 16598 6120
rect 16698 6260 16858 6280
rect 16698 6220 16708 6260
rect 16748 6220 16798 6260
rect 16838 6220 16858 6260
rect 16698 6160 16858 6220
rect 16698 6120 16708 6160
rect 16748 6120 16798 6160
rect 16838 6120 16858 6160
rect 16698 6100 16858 6120
rect 16908 6260 16988 6280
rect 16908 6220 16928 6260
rect 16968 6220 16988 6260
rect 16908 6160 16988 6220
rect 16908 6120 16928 6160
rect 16968 6120 16988 6160
rect 16908 6100 16988 6120
rect 17088 6260 17248 6280
rect 17088 6220 17098 6260
rect 17138 6220 17188 6260
rect 17228 6220 17248 6260
rect 17088 6160 17248 6220
rect 17088 6120 17098 6160
rect 17138 6120 17188 6160
rect 17228 6120 17248 6160
rect 17088 6100 17248 6120
rect 17298 6260 17378 6280
rect 17298 6220 17318 6260
rect 17358 6220 17378 6260
rect 17298 6160 17378 6220
rect 17298 6120 17318 6160
rect 17358 6120 17378 6160
rect 17298 6100 17378 6120
rect 17458 6260 17538 6280
rect 17458 6220 17478 6260
rect 17518 6220 17538 6260
rect 17458 6160 17538 6220
rect 17458 6120 17478 6160
rect 17518 6120 17538 6160
rect 17458 6100 17538 6120
rect 17588 6260 17668 6280
rect 17588 6220 17608 6260
rect 17648 6220 17668 6260
rect 17588 6160 17668 6220
rect 17588 6120 17608 6160
rect 17648 6120 17668 6160
rect 17588 6100 17668 6120
rect 13658 6040 13738 6060
rect 13658 6000 13678 6040
rect 13718 6000 13738 6040
rect 13658 5980 13738 6000
rect 13788 5950 13828 6100
rect 14008 5950 14048 6100
rect 14168 5950 14208 6100
rect 14388 5950 14428 6100
rect 14688 5950 14728 6100
rect 14908 5950 14948 6100
rect 15208 5950 15248 6100
rect 15378 6040 15458 6060
rect 15378 6000 15398 6040
rect 15438 6000 15458 6040
rect 15378 5980 15458 6000
rect 15648 5950 15688 6100
rect 15978 5950 16018 6100
rect 16408 5950 16448 6100
rect 16798 5950 16838 6100
rect 17188 5950 17228 6100
rect 17478 6060 17518 6100
rect 17458 6040 17538 6060
rect 17458 6000 17478 6040
rect 17518 6000 17538 6040
rect 17458 5980 17538 6000
rect 13248 5930 13328 5950
rect 13248 5890 13268 5930
rect 13308 5890 13328 5930
rect 13248 5870 13328 5890
rect 13468 5930 13548 5950
rect 13468 5890 13488 5930
rect 13528 5890 13548 5930
rect 13468 5870 13548 5890
rect 13768 5930 13848 5950
rect 13768 5890 13788 5930
rect 13828 5890 13848 5930
rect 13768 5870 13848 5890
rect 13988 5930 14068 5950
rect 13988 5890 14008 5930
rect 14048 5890 14068 5930
rect 13988 5870 14068 5890
rect 14148 5930 14228 5950
rect 14148 5890 14168 5930
rect 14208 5890 14228 5930
rect 14148 5870 14228 5890
rect 14368 5930 14448 5950
rect 14368 5890 14388 5930
rect 14428 5890 14448 5930
rect 14368 5870 14448 5890
rect 14668 5930 14748 5950
rect 14668 5890 14688 5930
rect 14728 5890 14748 5930
rect 14668 5870 14748 5890
rect 14888 5930 14968 5950
rect 14888 5890 14908 5930
rect 14948 5890 14968 5930
rect 14888 5870 14968 5890
rect 15188 5930 15268 5950
rect 15188 5890 15208 5930
rect 15248 5890 15268 5930
rect 15188 5870 15268 5890
rect 15628 5930 15708 5950
rect 15628 5890 15648 5930
rect 15688 5890 15708 5930
rect 15628 5870 15708 5890
rect 15958 5930 16038 5950
rect 15958 5890 15978 5930
rect 16018 5890 16038 5930
rect 15958 5870 16038 5890
rect 16388 5930 16468 5950
rect 16388 5890 16408 5930
rect 16448 5890 16468 5930
rect 16388 5870 16468 5890
rect 16778 5930 16858 5950
rect 16778 5890 16798 5930
rect 16838 5890 16858 5930
rect 16778 5870 16858 5890
rect 17168 5930 17248 5950
rect 17168 5890 17188 5930
rect 17228 5890 17248 5930
rect 17168 5870 17248 5890
rect 22978 5880 23088 5900
rect 22978 5810 22998 5880
rect 23068 5810 23088 5880
rect 22978 5790 23088 5810
rect 23578 5530 23658 5550
rect 24098 5530 24178 5550
rect 24618 5530 24698 5550
rect 25138 5530 25218 5550
rect 23088 5490 23598 5530
rect 23638 5490 24108 5530
rect 24268 5490 24638 5530
rect 24678 5490 25148 5530
rect 25218 5490 25318 5530
rect 23088 5060 23128 5490
rect 23578 5470 23658 5490
rect 24098 5470 24178 5490
rect 24618 5470 24698 5490
rect 25138 5470 25218 5490
rect 23208 5400 23268 5420
rect 23208 5360 23218 5400
rect 23258 5360 23268 5400
rect 23208 5300 23268 5360
rect 23208 5260 23218 5300
rect 23258 5260 23268 5300
rect 23208 5200 23268 5260
rect 23208 5160 23218 5200
rect 23258 5160 23268 5200
rect 23208 5100 23268 5160
rect 23208 5060 23218 5100
rect 23258 5060 23268 5100
rect 23208 5040 23268 5060
rect 23588 5400 23648 5420
rect 23588 5360 23598 5400
rect 23638 5360 23648 5400
rect 23588 5300 23648 5360
rect 23588 5260 23598 5300
rect 23638 5260 23648 5300
rect 23588 5200 23648 5260
rect 23588 5160 23598 5200
rect 23638 5160 23648 5200
rect 23588 5100 23648 5160
rect 23588 5060 23598 5100
rect 23638 5060 23648 5100
rect 23588 5040 23648 5060
rect 23728 5400 23788 5420
rect 23728 5360 23738 5400
rect 23778 5360 23788 5400
rect 23728 5300 23788 5360
rect 23728 5260 23738 5300
rect 23778 5260 23788 5300
rect 23728 5200 23788 5260
rect 23728 5160 23738 5200
rect 23778 5160 23788 5200
rect 23728 5100 23788 5160
rect 23728 5060 23738 5100
rect 23778 5060 23788 5100
rect 23728 5040 23788 5060
rect 24108 5400 24168 5420
rect 24108 5360 24118 5400
rect 24158 5360 24168 5400
rect 24108 5300 24168 5360
rect 24108 5260 24118 5300
rect 24158 5260 24168 5300
rect 24108 5200 24168 5260
rect 24108 5160 24118 5200
rect 24158 5160 24168 5200
rect 24108 5100 24168 5160
rect 24108 5060 24118 5100
rect 24158 5060 24168 5100
rect 24108 5040 24168 5060
rect 24248 5400 24308 5420
rect 24248 5360 24258 5400
rect 24298 5360 24308 5400
rect 24248 5300 24308 5360
rect 24248 5260 24258 5300
rect 24298 5260 24308 5300
rect 24248 5200 24308 5260
rect 24248 5160 24258 5200
rect 24298 5160 24308 5200
rect 24248 5100 24308 5160
rect 24248 5060 24258 5100
rect 24298 5060 24308 5100
rect 24248 5040 24308 5060
rect 24628 5400 24688 5420
rect 24628 5360 24638 5400
rect 24678 5360 24688 5400
rect 24628 5300 24688 5360
rect 24628 5260 24638 5300
rect 24678 5260 24688 5300
rect 24628 5200 24688 5260
rect 24628 5160 24638 5200
rect 24678 5160 24688 5200
rect 24628 5100 24688 5160
rect 24628 5060 24638 5100
rect 24678 5060 24688 5100
rect 24628 5040 24688 5060
rect 24768 5400 24828 5420
rect 24768 5360 24778 5400
rect 24818 5360 24828 5400
rect 24768 5300 24828 5360
rect 24768 5260 24778 5300
rect 24818 5260 24828 5300
rect 24768 5200 24828 5260
rect 24768 5160 24778 5200
rect 24818 5160 24828 5200
rect 24768 5100 24828 5160
rect 24768 5060 24778 5100
rect 24818 5060 24828 5100
rect 24768 5040 24828 5060
rect 25148 5400 25208 5420
rect 25148 5360 25158 5400
rect 25198 5360 25208 5400
rect 25148 5300 25208 5360
rect 25148 5260 25158 5300
rect 25198 5260 25208 5300
rect 25148 5200 25208 5260
rect 25148 5160 25158 5200
rect 25198 5160 25208 5200
rect 25148 5100 25208 5160
rect 25148 5060 25158 5100
rect 25198 5060 25208 5100
rect 25148 5040 25208 5060
rect 25278 5060 25318 5490
rect 23388 4980 23468 5000
rect 23388 4940 23408 4980
rect 23448 4940 23468 4980
rect 23388 4920 23468 4940
rect 23908 4980 23988 5000
rect 23908 4940 23928 4980
rect 23968 4940 23988 4980
rect 23908 4920 23988 4940
rect 24428 4980 24508 5000
rect 24428 4940 24448 4980
rect 24488 4940 24508 4980
rect 24428 4920 24508 4940
rect 24958 4980 25018 5000
rect 24958 4940 24968 4980
rect 25008 4940 25018 4980
rect 24958 4920 25018 4940
rect 12698 3730 12778 3750
rect 12698 3690 12718 3730
rect 12758 3690 12778 3730
rect 12698 3670 12778 3690
rect 13118 3730 13198 3750
rect 13118 3690 13138 3730
rect 13178 3690 13198 3730
rect 13118 3670 13198 3690
rect 13788 3730 13868 3750
rect 13788 3690 13808 3730
rect 13848 3690 13868 3730
rect 13788 3670 13868 3690
rect 14358 3730 14438 3750
rect 14358 3690 14378 3730
rect 14418 3690 14438 3730
rect 14358 3670 14438 3690
rect 15068 3730 15148 3750
rect 15068 3690 15088 3730
rect 15128 3690 15148 3730
rect 15068 3670 15148 3690
rect 15498 3730 15578 3750
rect 15498 3690 15518 3730
rect 15558 3690 15578 3730
rect 15498 3670 15578 3690
rect 15938 3730 16018 3750
rect 15938 3690 15958 3730
rect 15998 3690 16018 3730
rect 15938 3670 16018 3690
rect 16188 3730 16268 3750
rect 16188 3690 16208 3730
rect 16248 3690 16268 3730
rect 16188 3670 16268 3690
rect 16408 3730 16488 3750
rect 16408 3690 16428 3730
rect 16468 3690 16488 3730
rect 16408 3670 16488 3690
rect 16878 3730 16958 3750
rect 16878 3690 16898 3730
rect 16938 3690 16958 3730
rect 16878 3670 16958 3690
rect 17318 3730 17398 3750
rect 17318 3690 17338 3730
rect 17378 3690 17398 3730
rect 17318 3670 17398 3690
rect 17938 3730 18018 3750
rect 17938 3690 17958 3730
rect 17998 3690 18018 3730
rect 17938 3670 18018 3690
rect 18278 3730 18358 3750
rect 18278 3690 18298 3730
rect 18338 3690 18358 3730
rect 18278 3670 18358 3690
rect 18638 3730 18718 3750
rect 18638 3690 18658 3730
rect 18698 3690 18718 3730
rect 18638 3670 18718 3690
rect 19238 3730 19318 3750
rect 19238 3690 19258 3730
rect 19298 3690 19318 3730
rect 19238 3670 19318 3690
rect 19578 3730 19658 3750
rect 19578 3690 19598 3730
rect 19638 3690 19658 3730
rect 19578 3670 19658 3690
rect 19938 3730 20018 3750
rect 19938 3690 19958 3730
rect 19998 3690 20018 3730
rect 19938 3670 20018 3690
rect 20538 3730 20618 3750
rect 20538 3690 20558 3730
rect 20598 3690 20618 3730
rect 20538 3670 20618 3690
rect 20878 3730 20958 3750
rect 20878 3690 20898 3730
rect 20938 3690 20958 3730
rect 20878 3670 20958 3690
rect 21238 3730 21318 3750
rect 21238 3690 21258 3730
rect 21298 3690 21318 3730
rect 21238 3670 21318 3690
rect 21838 3730 21918 3750
rect 21838 3690 21858 3730
rect 21898 3690 21918 3730
rect 21838 3670 21918 3690
rect 22178 3730 22258 3750
rect 22178 3690 22198 3730
rect 22238 3690 22258 3730
rect 22178 3670 22258 3690
rect 22538 3730 22618 3750
rect 22538 3690 22558 3730
rect 22598 3690 22618 3730
rect 22538 3670 22618 3690
rect 12718 3520 12758 3670
rect 13018 3620 13098 3640
rect 13018 3580 13038 3620
rect 13078 3580 13098 3620
rect 13018 3560 13098 3580
rect 13138 3520 13178 3670
rect 13218 3620 13288 3640
rect 13218 3580 13228 3620
rect 13268 3580 13288 3620
rect 13218 3560 13288 3580
rect 13248 3520 13288 3560
rect 13328 3600 13408 3620
rect 13328 3560 13348 3600
rect 13388 3560 13408 3600
rect 13328 3540 13408 3560
rect 13808 3520 13848 3670
rect 14138 3620 14218 3640
rect 14138 3580 14158 3620
rect 14198 3580 14218 3620
rect 14138 3560 14218 3580
rect 14278 3620 14338 3640
rect 14278 3580 14288 3620
rect 14328 3580 14338 3620
rect 14278 3560 14338 3580
rect 14378 3520 14418 3670
rect 15088 3520 15128 3670
rect 15398 3620 15478 3640
rect 15398 3580 15418 3620
rect 15458 3580 15478 3620
rect 15398 3560 15478 3580
rect 15518 3520 15558 3670
rect 15618 3620 15698 3640
rect 15618 3580 15638 3620
rect 15678 3580 15698 3620
rect 15618 3560 15698 3580
rect 15618 3520 15658 3560
rect 15958 3520 15998 3670
rect 16208 3520 16248 3670
rect 16428 3520 16468 3670
rect 16748 3630 16828 3640
rect 16748 3590 16768 3630
rect 16808 3590 16828 3630
rect 16748 3570 16828 3590
rect 16788 3520 16828 3570
rect 16898 3520 16938 3670
rect 17158 3630 17238 3640
rect 17158 3590 17178 3630
rect 17218 3590 17238 3630
rect 17158 3570 17238 3590
rect 17338 3520 17378 3670
rect 17958 3520 17998 3670
rect 18298 3520 18338 3670
rect 18658 3520 18698 3670
rect 19108 3620 19188 3640
rect 19108 3580 19128 3620
rect 19168 3580 19188 3620
rect 19108 3560 19188 3580
rect 19148 3520 19188 3560
rect 19258 3520 19298 3670
rect 19598 3520 19638 3670
rect 19688 3620 19768 3640
rect 19688 3580 19708 3620
rect 19748 3580 19768 3620
rect 19688 3560 19768 3580
rect 19958 3520 19998 3670
rect 20408 3620 20488 3640
rect 20408 3580 20428 3620
rect 20468 3580 20488 3620
rect 20408 3560 20488 3580
rect 20448 3520 20488 3560
rect 20558 3520 20598 3670
rect 20898 3520 20938 3670
rect 20988 3620 21068 3640
rect 20988 3580 21008 3620
rect 21048 3580 21068 3620
rect 20988 3560 21068 3580
rect 21258 3520 21298 3670
rect 21708 3620 21788 3640
rect 21708 3580 21728 3620
rect 21768 3580 21788 3620
rect 21708 3560 21788 3580
rect 21748 3520 21788 3560
rect 21858 3520 21898 3670
rect 22198 3520 22238 3670
rect 22288 3620 22368 3640
rect 22288 3580 22308 3620
rect 22348 3580 22368 3620
rect 22288 3560 22368 3580
rect 22558 3520 22598 3670
rect 12358 3500 12438 3520
rect 12598 3500 12658 3520
rect 12358 3460 12378 3500
rect 12418 3460 12608 3500
rect 12648 3460 12658 3500
rect 12358 3440 12438 3460
rect 12598 3440 12658 3460
rect 12708 3500 12848 3520
rect 13018 3500 13078 3520
rect 12708 3460 12718 3500
rect 12758 3460 12798 3500
rect 12838 3460 12848 3500
rect 12708 3440 12848 3460
rect 12888 3460 13028 3500
rect 13068 3460 13078 3500
rect 12398 3350 12438 3440
rect 12318 3330 12438 3350
rect 12318 3290 12338 3330
rect 12378 3290 12438 3330
rect 12318 3270 12438 3290
rect 12398 3200 12438 3270
rect 12488 3300 12568 3320
rect 12488 3260 12508 3300
rect 12548 3280 12568 3300
rect 12888 3280 12928 3460
rect 13018 3440 13078 3460
rect 13128 3500 13188 3520
rect 13128 3460 13138 3500
rect 13178 3460 13188 3500
rect 13128 3440 13188 3460
rect 13238 3500 13298 3520
rect 13688 3500 13748 3520
rect 13238 3460 13248 3500
rect 13288 3460 13298 3500
rect 13238 3440 13298 3460
rect 13468 3460 13698 3500
rect 13738 3460 13748 3500
rect 13248 3400 13288 3440
rect 12548 3260 12928 3280
rect 12488 3240 12928 3260
rect 12668 3200 12708 3240
rect 12888 3200 12928 3240
rect 12978 3360 13288 3400
rect 12978 3200 13018 3360
rect 13468 3320 13508 3460
rect 13688 3440 13748 3460
rect 13798 3500 13858 3520
rect 13798 3460 13808 3500
rect 13848 3460 13858 3500
rect 13798 3440 13858 3460
rect 13908 3500 13968 3520
rect 13908 3460 13918 3500
rect 13958 3460 13968 3500
rect 13908 3440 13968 3460
rect 14128 3500 14188 3520
rect 14128 3460 14138 3500
rect 14178 3460 14188 3500
rect 14128 3440 14188 3460
rect 14238 3500 14298 3520
rect 14238 3460 14248 3500
rect 14288 3460 14298 3500
rect 14238 3440 14298 3460
rect 14348 3500 14418 3520
rect 14348 3460 14358 3500
rect 14398 3460 14418 3500
rect 14348 3440 14418 3460
rect 14458 3500 14518 3520
rect 14458 3460 14468 3500
rect 14508 3460 14518 3500
rect 14458 3440 14518 3460
rect 14728 3500 14808 3520
rect 14968 3500 15028 3520
rect 14728 3460 14748 3500
rect 14788 3460 14978 3500
rect 15018 3460 15028 3500
rect 14728 3440 14808 3460
rect 14968 3440 15028 3460
rect 15078 3500 15218 3520
rect 15388 3500 15448 3520
rect 15078 3460 15088 3500
rect 15128 3460 15168 3500
rect 15208 3460 15218 3500
rect 15078 3440 15218 3460
rect 15258 3460 15398 3500
rect 15438 3460 15448 3500
rect 13608 3380 13688 3400
rect 13608 3340 13628 3380
rect 13668 3340 13688 3380
rect 13608 3320 13688 3340
rect 13068 3300 13148 3320
rect 13408 3300 13508 3320
rect 13068 3260 13088 3300
rect 13128 3260 13428 3300
rect 13468 3260 13508 3300
rect 13068 3240 13148 3260
rect 13408 3240 13508 3260
rect 13648 3280 13688 3320
rect 13908 3280 13948 3440
rect 14008 3420 14088 3440
rect 14008 3380 14028 3420
rect 14068 3400 14088 3420
rect 14138 3400 14178 3440
rect 14468 3400 14508 3440
rect 14068 3380 14668 3400
rect 14008 3360 14668 3380
rect 13648 3240 13948 3280
rect 13988 3300 14068 3310
rect 13988 3260 14008 3300
rect 14048 3260 14068 3300
rect 14508 3300 14588 3310
rect 13988 3240 14068 3260
rect 14138 3240 14398 3280
rect 14508 3260 14528 3300
rect 14568 3260 14588 3300
rect 14508 3240 14588 3260
rect 13468 3200 13508 3240
rect 13688 3200 13728 3240
rect 13908 3200 13948 3240
rect 14138 3200 14178 3240
rect 14358 3200 14398 3240
rect 14628 3200 14668 3360
rect 12398 3180 12498 3200
rect 12398 3140 12448 3180
rect 12488 3140 12498 3180
rect 12398 3120 12498 3140
rect 12548 3180 12608 3200
rect 12548 3140 12558 3180
rect 12598 3140 12608 3180
rect 12548 3120 12608 3140
rect 12658 3180 12718 3200
rect 12658 3140 12668 3180
rect 12708 3140 12718 3180
rect 12658 3120 12718 3140
rect 12768 3180 12828 3200
rect 12768 3140 12778 3180
rect 12818 3140 12828 3180
rect 12768 3120 12828 3140
rect 12878 3180 12938 3200
rect 12878 3140 12888 3180
rect 12928 3140 12938 3180
rect 12978 3180 13078 3200
rect 12978 3140 13028 3180
rect 13068 3140 13078 3180
rect 12878 3120 12938 3140
rect 13018 3120 13078 3140
rect 13128 3180 13188 3200
rect 13128 3140 13138 3180
rect 13178 3140 13188 3180
rect 13128 3120 13188 3140
rect 13238 3180 13298 3200
rect 13238 3140 13248 3180
rect 13288 3140 13298 3180
rect 13238 3120 13298 3140
rect 13468 3180 13528 3200
rect 13468 3140 13478 3180
rect 13518 3140 13528 3180
rect 13468 3120 13528 3140
rect 13578 3180 13638 3200
rect 13578 3140 13588 3180
rect 13628 3140 13638 3180
rect 13578 3120 13638 3140
rect 13688 3180 13748 3200
rect 13688 3140 13698 3180
rect 13738 3140 13748 3180
rect 13688 3120 13748 3140
rect 13798 3180 13858 3200
rect 13798 3140 13808 3180
rect 13848 3140 13858 3180
rect 13798 3120 13858 3140
rect 13908 3180 13968 3200
rect 13908 3140 13918 3180
rect 13958 3140 13968 3180
rect 13908 3120 13968 3140
rect 14128 3180 14188 3200
rect 14128 3140 14138 3180
rect 14178 3140 14188 3180
rect 14128 3120 14188 3140
rect 14238 3180 14298 3200
rect 14238 3140 14248 3180
rect 14288 3140 14298 3180
rect 14238 3120 14298 3140
rect 14348 3180 14408 3200
rect 14348 3140 14358 3180
rect 14398 3140 14408 3180
rect 14348 3120 14408 3140
rect 14458 3180 14518 3200
rect 14458 3140 14468 3180
rect 14508 3140 14518 3180
rect 14458 3120 14518 3140
rect 14568 3180 14668 3200
rect 14568 3140 14578 3180
rect 14618 3140 14668 3180
rect 14768 3200 14808 3440
rect 14858 3300 14938 3310
rect 14858 3260 14878 3300
rect 14918 3280 14938 3300
rect 15258 3280 15298 3460
rect 15388 3440 15448 3460
rect 15498 3500 15558 3520
rect 15498 3460 15508 3500
rect 15548 3460 15558 3500
rect 15498 3440 15558 3460
rect 15608 3500 15668 3520
rect 15608 3460 15618 3500
rect 15658 3460 15668 3500
rect 15608 3440 15668 3460
rect 15838 3500 15898 3520
rect 15838 3460 15848 3500
rect 15888 3460 15898 3500
rect 15838 3440 15898 3460
rect 15948 3500 16008 3520
rect 15948 3460 15958 3500
rect 15998 3460 16008 3500
rect 15948 3440 16008 3460
rect 16058 3500 16118 3520
rect 16058 3460 16068 3500
rect 16108 3460 16118 3500
rect 16058 3440 16118 3460
rect 16198 3500 16258 3520
rect 16198 3460 16208 3500
rect 16248 3460 16258 3500
rect 16198 3440 16258 3460
rect 16308 3500 16368 3520
rect 16308 3460 16318 3500
rect 16358 3460 16368 3500
rect 16308 3440 16368 3460
rect 16418 3500 16478 3520
rect 16778 3500 16838 3520
rect 16418 3460 16428 3500
rect 16468 3460 16478 3500
rect 16418 3440 16478 3460
rect 16558 3460 16788 3500
rect 16828 3460 16838 3500
rect 15618 3400 15658 3440
rect 14918 3260 15298 3280
rect 14858 3240 15298 3260
rect 15038 3200 15078 3240
rect 15258 3200 15298 3240
rect 15348 3360 15658 3400
rect 15708 3420 15788 3440
rect 15708 3380 15728 3420
rect 15768 3400 15788 3420
rect 15848 3400 15888 3440
rect 16068 3400 16108 3440
rect 15768 3380 16108 3400
rect 15708 3360 16108 3380
rect 15348 3200 15388 3360
rect 15438 3300 15518 3320
rect 15648 3300 15728 3310
rect 15438 3260 15458 3300
rect 15498 3260 15668 3300
rect 15708 3260 15728 3300
rect 15438 3240 15518 3260
rect 15648 3240 15728 3260
rect 14768 3180 14868 3200
rect 14768 3140 14818 3180
rect 14858 3140 14868 3180
rect 14568 3120 14628 3140
rect 14808 3120 14868 3140
rect 14918 3180 14978 3200
rect 14918 3140 14928 3180
rect 14968 3140 14978 3180
rect 14918 3120 14978 3140
rect 15028 3180 15088 3200
rect 15028 3140 15038 3180
rect 15078 3140 15088 3180
rect 15028 3120 15088 3140
rect 15138 3180 15198 3200
rect 15138 3140 15148 3180
rect 15188 3140 15198 3180
rect 15138 3120 15198 3140
rect 15248 3180 15308 3200
rect 15248 3140 15258 3180
rect 15298 3140 15308 3180
rect 15348 3180 15448 3200
rect 15348 3140 15398 3180
rect 15438 3140 15448 3180
rect 15248 3120 15308 3140
rect 15388 3120 15448 3140
rect 15498 3180 15558 3200
rect 15498 3140 15508 3180
rect 15548 3140 15558 3180
rect 15498 3120 15558 3140
rect 15608 3180 15748 3200
rect 15608 3140 15618 3180
rect 15658 3140 15698 3180
rect 15738 3140 15748 3180
rect 15788 3180 15828 3360
rect 16318 3330 16358 3440
rect 16558 3370 16598 3460
rect 16778 3440 16838 3460
rect 16888 3500 16948 3520
rect 16888 3460 16898 3500
rect 16938 3460 16948 3500
rect 16888 3440 16948 3460
rect 16998 3500 17058 3520
rect 16998 3460 17008 3500
rect 17048 3460 17058 3500
rect 16998 3440 17058 3460
rect 17218 3500 17278 3520
rect 17218 3460 17228 3500
rect 17268 3460 17278 3500
rect 17218 3440 17278 3460
rect 17328 3500 17388 3520
rect 17328 3460 17338 3500
rect 17378 3460 17388 3500
rect 17328 3440 17388 3460
rect 17438 3500 17498 3520
rect 17688 3500 17768 3520
rect 17838 3500 17898 3520
rect 17438 3460 17448 3500
rect 17488 3460 17648 3500
rect 17438 3440 17498 3460
rect 16228 3320 16358 3330
rect 15888 3310 16358 3320
rect 15888 3300 16248 3310
rect 15888 3260 15908 3300
rect 15948 3280 16248 3300
rect 15948 3260 15968 3280
rect 15888 3240 15968 3260
rect 16228 3270 16248 3280
rect 16288 3270 16358 3310
rect 16498 3350 16598 3370
rect 16498 3310 16518 3350
rect 16558 3310 16598 3350
rect 16698 3380 16778 3400
rect 16698 3340 16718 3380
rect 16758 3340 16778 3380
rect 16698 3320 16778 3340
rect 16498 3290 16598 3310
rect 16228 3250 16358 3270
rect 16318 3200 16358 3250
rect 16558 3200 16598 3290
rect 16738 3280 16778 3320
rect 16998 3280 17038 3440
rect 17098 3420 17178 3440
rect 17098 3380 17118 3420
rect 17158 3400 17178 3420
rect 17228 3400 17268 3440
rect 17448 3400 17488 3440
rect 17158 3380 17488 3400
rect 17098 3360 17488 3380
rect 16738 3240 17038 3280
rect 17128 3300 17208 3310
rect 17488 3300 17568 3310
rect 17128 3260 17148 3300
rect 17188 3260 17508 3300
rect 17548 3260 17568 3300
rect 17128 3240 17208 3260
rect 17488 3240 17568 3260
rect 16778 3200 16818 3240
rect 16998 3200 17038 3240
rect 17608 3200 17648 3460
rect 17688 3460 17708 3500
rect 17748 3460 17848 3500
rect 17888 3460 17898 3500
rect 17688 3440 17768 3460
rect 17838 3440 17898 3460
rect 17948 3500 18088 3520
rect 17948 3460 17958 3500
rect 17998 3460 18038 3500
rect 18078 3460 18088 3500
rect 17948 3440 18088 3460
rect 18148 3500 18238 3520
rect 18148 3460 18188 3500
rect 18228 3460 18238 3500
rect 18148 3440 18238 3460
rect 18288 3500 18348 3520
rect 18288 3460 18298 3500
rect 18338 3460 18348 3500
rect 18288 3440 18348 3460
rect 18398 3500 18458 3520
rect 18398 3460 18408 3500
rect 18448 3460 18458 3500
rect 18398 3440 18458 3460
rect 18538 3500 18598 3520
rect 18538 3460 18548 3500
rect 18588 3460 18598 3500
rect 18538 3440 18598 3460
rect 18648 3500 18708 3520
rect 18648 3460 18658 3500
rect 18698 3460 18708 3500
rect 18648 3440 18708 3460
rect 18758 3500 18818 3520
rect 19138 3500 19198 3520
rect 18758 3460 18768 3500
rect 18808 3460 18818 3500
rect 18758 3440 18818 3460
rect 19028 3460 19148 3500
rect 19188 3460 19198 3500
rect 15948 3180 16008 3200
rect 15788 3140 15958 3180
rect 15998 3140 16008 3180
rect 15608 3120 15748 3140
rect 15948 3120 16008 3140
rect 16058 3180 16118 3200
rect 16058 3140 16068 3180
rect 16108 3140 16118 3180
rect 16058 3120 16118 3140
rect 16308 3180 16368 3200
rect 16308 3140 16318 3180
rect 16358 3140 16368 3180
rect 16308 3120 16368 3140
rect 16418 3180 16478 3200
rect 16418 3140 16428 3180
rect 16468 3140 16478 3180
rect 16418 3120 16478 3140
rect 16558 3180 16618 3200
rect 16558 3140 16568 3180
rect 16608 3140 16618 3180
rect 16558 3120 16618 3140
rect 16668 3180 16728 3200
rect 16668 3140 16678 3180
rect 16718 3140 16728 3180
rect 16668 3120 16728 3140
rect 16778 3180 16838 3200
rect 16778 3140 16788 3180
rect 16828 3140 16838 3180
rect 16778 3120 16838 3140
rect 16888 3180 16948 3200
rect 16888 3140 16898 3180
rect 16938 3140 16948 3180
rect 16888 3120 16948 3140
rect 16998 3180 17058 3200
rect 16998 3140 17008 3180
rect 17048 3140 17058 3180
rect 16998 3120 17058 3140
rect 17138 3180 17278 3200
rect 17138 3140 17148 3180
rect 17188 3140 17228 3180
rect 17268 3140 17278 3180
rect 17138 3120 17278 3140
rect 17328 3180 17388 3200
rect 17328 3140 17338 3180
rect 17378 3140 17388 3180
rect 17328 3120 17388 3140
rect 17438 3180 17498 3200
rect 17438 3140 17448 3180
rect 17488 3140 17498 3180
rect 17438 3120 17498 3140
rect 17548 3180 17648 3200
rect 17548 3140 17558 3180
rect 17598 3140 17648 3180
rect 17728 3200 17768 3440
rect 17818 3300 17898 3310
rect 17818 3260 17838 3300
rect 17878 3280 17898 3300
rect 18148 3280 18188 3440
rect 18408 3400 18448 3440
rect 18228 3380 18448 3400
rect 18228 3340 18248 3380
rect 18288 3360 18448 3380
rect 18288 3340 18348 3360
rect 18228 3320 18348 3340
rect 17878 3260 18258 3280
rect 17818 3240 18258 3260
rect 17998 3200 18038 3240
rect 18218 3200 18258 3240
rect 18308 3200 18348 3320
rect 18398 3300 18478 3320
rect 18398 3260 18418 3300
rect 18458 3280 18478 3300
rect 18548 3280 18588 3440
rect 18768 3280 18808 3440
rect 19028 3340 19068 3460
rect 19138 3440 19198 3460
rect 19248 3500 19388 3520
rect 19248 3460 19258 3500
rect 19298 3460 19338 3500
rect 19378 3460 19388 3500
rect 19248 3440 19388 3460
rect 19448 3500 19538 3520
rect 19448 3460 19488 3500
rect 19528 3460 19538 3500
rect 19448 3440 19538 3460
rect 19588 3500 19648 3520
rect 19588 3460 19598 3500
rect 19638 3460 19648 3500
rect 19588 3440 19648 3460
rect 19698 3500 19758 3520
rect 19698 3460 19708 3500
rect 19748 3460 19758 3500
rect 19698 3440 19758 3460
rect 19838 3500 19898 3520
rect 19838 3460 19848 3500
rect 19888 3460 19898 3500
rect 19838 3440 19898 3460
rect 19948 3500 20008 3520
rect 19948 3460 19958 3500
rect 19998 3460 20008 3500
rect 19948 3440 20008 3460
rect 20058 3500 20118 3520
rect 20438 3500 20498 3520
rect 20058 3460 20068 3500
rect 20108 3460 20118 3500
rect 20058 3440 20118 3460
rect 20328 3460 20448 3500
rect 20488 3460 20498 3500
rect 18458 3260 18808 3280
rect 18868 3320 19068 3340
rect 18868 3280 18888 3320
rect 18928 3300 19068 3320
rect 18928 3280 18948 3300
rect 18868 3260 18948 3280
rect 18398 3240 18808 3260
rect 18768 3200 18808 3240
rect 17728 3180 17828 3200
rect 17728 3140 17778 3180
rect 17818 3140 17828 3180
rect 17548 3120 17608 3140
rect 17768 3120 17828 3140
rect 17878 3180 17938 3200
rect 17878 3140 17888 3180
rect 17928 3140 17938 3180
rect 17878 3120 17938 3140
rect 17988 3180 18048 3200
rect 17988 3140 17998 3180
rect 18038 3140 18048 3180
rect 17988 3120 18048 3140
rect 18098 3180 18158 3200
rect 18098 3140 18108 3180
rect 18148 3140 18158 3180
rect 18098 3120 18158 3140
rect 18208 3180 18268 3200
rect 18208 3140 18218 3180
rect 18258 3140 18268 3180
rect 18308 3180 18488 3200
rect 18308 3160 18438 3180
rect 18208 3120 18268 3140
rect 18428 3140 18438 3160
rect 18478 3140 18488 3180
rect 18428 3120 18488 3140
rect 18538 3180 18598 3200
rect 18538 3140 18548 3180
rect 18588 3140 18598 3180
rect 18538 3120 18598 3140
rect 18648 3180 18718 3200
rect 18648 3140 18658 3180
rect 18698 3140 18718 3180
rect 18648 3120 18718 3140
rect 18758 3180 18818 3200
rect 18758 3140 18768 3180
rect 18808 3140 18818 3180
rect 18758 3120 18818 3140
rect 12398 3080 12438 3120
rect 12378 3060 12458 3080
rect 12378 3020 12398 3060
rect 12438 3020 12458 3060
rect 12378 3000 12458 3020
rect 12558 2970 12598 3120
rect 12778 2970 12818 3120
rect 13248 2970 13288 3120
rect 13328 3080 13408 3100
rect 13478 3080 13518 3120
rect 13328 3040 13348 3080
rect 13388 3040 13408 3080
rect 13328 3020 13408 3040
rect 13458 3070 13538 3080
rect 13458 3030 13478 3070
rect 13518 3030 13538 3070
rect 13458 3010 13538 3030
rect 13588 2970 13628 3120
rect 13808 2970 13848 3120
rect 14248 2970 14288 3120
rect 14398 3070 14478 3080
rect 14398 3030 14418 3070
rect 14458 3030 14478 3070
rect 14398 3010 14478 3030
rect 14928 2970 14968 3120
rect 15148 2970 15188 3120
rect 15618 2970 15658 3120
rect 15958 3070 16038 3080
rect 15958 3030 15978 3070
rect 16018 3030 16038 3070
rect 15958 3010 16038 3030
rect 16078 2970 16118 3120
rect 16428 2970 16468 3120
rect 16678 2970 16718 3120
rect 16898 2970 16938 3120
rect 17228 2970 17268 3120
rect 17888 2970 17928 3120
rect 18108 2970 18148 3120
rect 18572 3060 18638 3080
rect 18572 3020 18582 3060
rect 18622 3020 18638 3060
rect 18572 3000 18638 3020
rect 18678 2970 18718 3120
rect 19028 3110 19068 3300
rect 19118 3210 19198 3230
rect 19118 3170 19138 3210
rect 19178 3190 19198 3210
rect 19448 3190 19488 3440
rect 19708 3400 19748 3440
rect 19528 3380 19748 3400
rect 19528 3340 19548 3380
rect 19588 3360 19748 3380
rect 19588 3340 19648 3360
rect 19528 3320 19648 3340
rect 19178 3170 19558 3190
rect 19118 3150 19558 3170
rect 19298 3110 19338 3150
rect 19518 3110 19558 3150
rect 19608 3110 19648 3320
rect 19698 3210 19778 3230
rect 19698 3170 19718 3210
rect 19758 3190 19778 3210
rect 19848 3190 19888 3440
rect 20068 3190 20108 3440
rect 20328 3340 20368 3460
rect 20438 3440 20498 3460
rect 20548 3500 20688 3520
rect 20548 3460 20558 3500
rect 20598 3460 20638 3500
rect 20678 3460 20688 3500
rect 20548 3440 20688 3460
rect 20748 3500 20838 3520
rect 20748 3460 20788 3500
rect 20828 3460 20838 3500
rect 20748 3440 20838 3460
rect 20888 3500 20948 3520
rect 20888 3460 20898 3500
rect 20938 3460 20948 3500
rect 20888 3440 20948 3460
rect 20998 3500 21058 3520
rect 20998 3460 21008 3500
rect 21048 3460 21058 3500
rect 20998 3440 21058 3460
rect 21138 3500 21198 3520
rect 21138 3460 21148 3500
rect 21188 3460 21198 3500
rect 21138 3440 21198 3460
rect 21248 3500 21308 3520
rect 21248 3460 21258 3500
rect 21298 3460 21308 3500
rect 21248 3440 21308 3460
rect 21358 3500 21418 3520
rect 21738 3500 21798 3520
rect 21358 3460 21368 3500
rect 21408 3460 21418 3500
rect 21358 3440 21418 3460
rect 21628 3460 21748 3500
rect 21788 3460 21798 3500
rect 20168 3320 20368 3340
rect 20168 3280 20188 3320
rect 20228 3300 20368 3320
rect 20228 3280 20248 3300
rect 20168 3260 20248 3280
rect 19758 3170 20108 3190
rect 19698 3150 20108 3170
rect 20068 3110 20108 3150
rect 20328 3110 20368 3300
rect 20418 3210 20498 3230
rect 20418 3170 20438 3210
rect 20478 3190 20498 3210
rect 20748 3190 20788 3440
rect 21008 3400 21048 3440
rect 20828 3380 21048 3400
rect 20828 3340 20848 3380
rect 20888 3360 21048 3380
rect 20888 3340 20948 3360
rect 20828 3320 20948 3340
rect 20478 3170 20858 3190
rect 20418 3150 20858 3170
rect 20598 3110 20638 3150
rect 20818 3110 20858 3150
rect 20908 3110 20948 3320
rect 20998 3210 21078 3230
rect 20998 3170 21018 3210
rect 21058 3190 21078 3210
rect 21148 3190 21188 3440
rect 21368 3190 21408 3440
rect 21628 3340 21668 3460
rect 21738 3440 21798 3460
rect 21848 3500 21988 3520
rect 21848 3460 21858 3500
rect 21898 3460 21938 3500
rect 21978 3460 21988 3500
rect 21848 3440 21988 3460
rect 22048 3500 22138 3520
rect 22048 3460 22088 3500
rect 22128 3460 22138 3500
rect 22048 3440 22138 3460
rect 22188 3500 22248 3520
rect 22188 3460 22198 3500
rect 22238 3460 22248 3500
rect 22188 3440 22248 3460
rect 22298 3500 22358 3520
rect 22298 3460 22308 3500
rect 22348 3460 22358 3500
rect 22298 3440 22358 3460
rect 22438 3500 22498 3520
rect 22438 3460 22448 3500
rect 22488 3460 22498 3500
rect 22438 3440 22498 3460
rect 22548 3500 22608 3520
rect 22548 3460 22558 3500
rect 22598 3460 22608 3500
rect 22548 3440 22608 3460
rect 22658 3500 22718 3520
rect 22658 3460 22668 3500
rect 22708 3460 22718 3500
rect 22658 3440 22718 3460
rect 21468 3320 21668 3340
rect 21468 3280 21488 3320
rect 21528 3300 21668 3320
rect 21528 3280 21548 3300
rect 21468 3260 21548 3280
rect 21058 3170 21408 3190
rect 20998 3150 21408 3170
rect 21368 3110 21408 3150
rect 21628 3110 21668 3300
rect 21718 3210 21798 3230
rect 21718 3170 21738 3210
rect 21778 3190 21798 3210
rect 22048 3190 22088 3440
rect 22308 3400 22348 3440
rect 22128 3380 22348 3400
rect 22128 3340 22148 3380
rect 22188 3360 22348 3380
rect 22188 3340 22248 3360
rect 22128 3320 22248 3340
rect 21778 3170 22158 3190
rect 21718 3150 22158 3170
rect 21898 3110 21938 3150
rect 22118 3110 22158 3150
rect 22208 3110 22248 3320
rect 22298 3210 22378 3230
rect 22298 3170 22318 3210
rect 22358 3190 22378 3210
rect 22448 3190 22488 3440
rect 22668 3190 22708 3440
rect 23088 3420 23128 4730
rect 23208 4710 23268 4730
rect 23208 4670 23218 4710
rect 23258 4670 23268 4710
rect 23208 4610 23268 4670
rect 23208 4570 23218 4610
rect 23258 4570 23268 4610
rect 23208 4510 23268 4570
rect 23208 4470 23218 4510
rect 23258 4470 23268 4510
rect 23208 4410 23268 4470
rect 23208 4370 23218 4410
rect 23258 4370 23268 4410
rect 23208 4310 23268 4370
rect 23208 4270 23218 4310
rect 23258 4270 23268 4310
rect 23208 4210 23268 4270
rect 23208 4170 23218 4210
rect 23258 4170 23268 4210
rect 23208 4150 23268 4170
rect 23318 4710 23378 4730
rect 23318 4670 23328 4710
rect 23368 4670 23378 4710
rect 23318 4610 23378 4670
rect 23318 4570 23328 4610
rect 23368 4570 23378 4610
rect 23318 4510 23378 4570
rect 23318 4470 23328 4510
rect 23368 4470 23378 4510
rect 23318 4410 23378 4470
rect 23318 4370 23328 4410
rect 23368 4370 23378 4410
rect 23318 4310 23378 4370
rect 23318 4270 23328 4310
rect 23368 4270 23378 4310
rect 23318 4210 23378 4270
rect 23318 4170 23328 4210
rect 23368 4170 23378 4210
rect 23318 4150 23378 4170
rect 23728 4710 23788 4730
rect 23728 4670 23738 4710
rect 23778 4670 23788 4710
rect 23728 4610 23788 4670
rect 23728 4570 23738 4610
rect 23778 4570 23788 4610
rect 23728 4510 23788 4570
rect 23728 4470 23738 4510
rect 23778 4470 23788 4510
rect 23728 4410 23788 4470
rect 23728 4370 23738 4410
rect 23778 4370 23788 4410
rect 23728 4310 23788 4370
rect 23728 4270 23738 4310
rect 23778 4270 23788 4310
rect 23728 4210 23788 4270
rect 23728 4170 23738 4210
rect 23778 4170 23788 4210
rect 23728 4150 23788 4170
rect 23838 4710 23898 4730
rect 23838 4670 23848 4710
rect 23888 4670 23898 4710
rect 23838 4610 23898 4670
rect 23838 4570 23848 4610
rect 23888 4570 23898 4610
rect 23838 4510 23898 4570
rect 23838 4470 23848 4510
rect 23888 4470 23898 4510
rect 23838 4410 23898 4470
rect 23838 4370 23848 4410
rect 23888 4370 23898 4410
rect 23838 4310 23898 4370
rect 23838 4270 23848 4310
rect 23888 4270 23898 4310
rect 23838 4210 23898 4270
rect 23838 4170 23848 4210
rect 23888 4170 23898 4210
rect 23838 4150 23898 4170
rect 24248 4710 24308 4730
rect 24248 4670 24258 4710
rect 24298 4670 24308 4710
rect 24248 4610 24308 4670
rect 24248 4570 24258 4610
rect 24298 4570 24308 4610
rect 24248 4510 24308 4570
rect 24248 4470 24258 4510
rect 24298 4470 24308 4510
rect 24248 4410 24308 4470
rect 24248 4370 24258 4410
rect 24298 4370 24308 4410
rect 24248 4310 24308 4370
rect 24248 4270 24258 4310
rect 24298 4270 24308 4310
rect 24248 4210 24308 4270
rect 24248 4170 24258 4210
rect 24298 4170 24308 4210
rect 24248 4150 24308 4170
rect 24358 4710 24418 4730
rect 24358 4670 24368 4710
rect 24408 4670 24418 4710
rect 24358 4610 24418 4670
rect 24358 4570 24368 4610
rect 24408 4570 24418 4610
rect 24358 4510 24418 4570
rect 24358 4470 24368 4510
rect 24408 4470 24418 4510
rect 24358 4410 24418 4470
rect 24358 4370 24368 4410
rect 24408 4370 24418 4410
rect 24358 4310 24418 4370
rect 24358 4270 24368 4310
rect 24408 4270 24418 4310
rect 24358 4210 24418 4270
rect 24358 4170 24368 4210
rect 24408 4170 24418 4210
rect 24358 4150 24418 4170
rect 23278 4092 23336 4110
rect 23278 4058 23290 4092
rect 23324 4058 23336 4092
rect 23278 4040 23336 4058
rect 23798 4092 23856 4110
rect 23798 4058 23810 4092
rect 23844 4058 23856 4092
rect 23798 4040 23856 4058
rect 24318 4092 24376 4110
rect 24318 4058 24330 4092
rect 24364 4058 24376 4092
rect 24318 4040 24376 4058
rect 23206 3930 23266 3950
rect 23206 3890 23216 3930
rect 23256 3890 23266 3930
rect 23206 3830 23266 3890
rect 23206 3790 23216 3830
rect 23256 3790 23266 3830
rect 23206 3730 23266 3790
rect 23206 3690 23216 3730
rect 23256 3690 23266 3730
rect 23206 3630 23266 3690
rect 23206 3590 23216 3630
rect 23256 3590 23266 3630
rect 23206 3570 23266 3590
rect 23318 3930 23378 3950
rect 23318 3890 23328 3930
rect 23368 3890 23378 3930
rect 23318 3830 23378 3890
rect 23318 3790 23328 3830
rect 23368 3790 23378 3830
rect 23318 3730 23378 3790
rect 23318 3690 23328 3730
rect 23368 3690 23378 3730
rect 23318 3630 23378 3690
rect 23318 3590 23328 3630
rect 23368 3590 23378 3630
rect 23318 3570 23378 3590
rect 23726 3930 23786 3950
rect 23726 3890 23736 3930
rect 23776 3890 23786 3930
rect 23726 3830 23786 3890
rect 23726 3790 23736 3830
rect 23776 3790 23786 3830
rect 23726 3730 23786 3790
rect 23726 3690 23736 3730
rect 23776 3690 23786 3730
rect 23726 3630 23786 3690
rect 23726 3590 23736 3630
rect 23776 3590 23786 3630
rect 23726 3570 23786 3590
rect 23838 3930 23898 3950
rect 23838 3890 23848 3930
rect 23888 3890 23898 3930
rect 23838 3830 23898 3890
rect 23838 3790 23848 3830
rect 23888 3790 23898 3830
rect 23838 3730 23898 3790
rect 23838 3690 23848 3730
rect 23888 3690 23898 3730
rect 23838 3630 23898 3690
rect 23838 3590 23848 3630
rect 23888 3590 23898 3630
rect 23838 3570 23898 3590
rect 24246 3930 24306 3950
rect 24246 3890 24256 3930
rect 24296 3890 24306 3930
rect 24246 3830 24306 3890
rect 24246 3790 24256 3830
rect 24296 3790 24306 3830
rect 24246 3730 24306 3790
rect 24246 3690 24256 3730
rect 24296 3690 24306 3730
rect 24246 3630 24306 3690
rect 24246 3590 24256 3630
rect 24296 3590 24306 3630
rect 24246 3570 24306 3590
rect 24358 3930 24418 3950
rect 24358 3890 24368 3930
rect 24408 3890 24418 3930
rect 24358 3830 24418 3890
rect 24358 3790 24368 3830
rect 24408 3790 24418 3830
rect 24358 3730 24418 3790
rect 24358 3690 24368 3730
rect 24408 3690 24418 3730
rect 24358 3630 24418 3690
rect 24358 3590 24368 3630
rect 24408 3590 24418 3630
rect 24358 3570 24418 3590
rect 23250 3512 23308 3530
rect 23250 3478 23262 3512
rect 23296 3478 23308 3512
rect 23250 3460 23308 3478
rect 23770 3512 23828 3530
rect 23770 3478 23782 3512
rect 23816 3478 23828 3512
rect 23770 3460 23828 3478
rect 24290 3512 24348 3530
rect 24290 3478 24302 3512
rect 24336 3478 24348 3512
rect 24290 3460 24348 3478
rect 25278 3420 25318 4730
rect 23088 3380 24108 3420
rect 24268 3380 25318 3420
rect 22750 3322 22808 3340
rect 22750 3288 22762 3322
rect 22796 3288 22808 3322
rect 22750 3260 22808 3288
rect 22358 3170 22708 3190
rect 22298 3150 22708 3170
rect 22668 3110 22708 3150
rect 23088 3180 24228 3220
rect 24368 3180 25128 3220
rect 18928 3090 18988 3110
rect 18928 3050 18938 3090
rect 18978 3050 18988 3090
rect 19028 3090 19128 3110
rect 19028 3050 19078 3090
rect 19118 3050 19128 3090
rect 18928 3030 18988 3050
rect 19068 3030 19128 3050
rect 19178 3090 19238 3110
rect 19178 3050 19188 3090
rect 19228 3050 19238 3090
rect 19178 3030 19238 3050
rect 19288 3090 19348 3110
rect 19288 3050 19298 3090
rect 19338 3050 19348 3090
rect 19288 3030 19348 3050
rect 19398 3090 19458 3110
rect 19398 3050 19408 3090
rect 19448 3050 19458 3090
rect 19398 3030 19458 3050
rect 19508 3090 19568 3110
rect 19508 3050 19518 3090
rect 19558 3050 19568 3090
rect 19608 3090 19788 3110
rect 19608 3070 19738 3090
rect 19508 3030 19568 3050
rect 19728 3050 19738 3070
rect 19778 3050 19788 3090
rect 19728 3030 19788 3050
rect 19838 3090 19898 3110
rect 19838 3050 19848 3090
rect 19888 3050 19898 3090
rect 19838 3030 19898 3050
rect 19948 3090 20008 3110
rect 19948 3050 19958 3090
rect 19998 3050 20008 3090
rect 19948 3030 20008 3050
rect 20058 3090 20118 3110
rect 20058 3050 20068 3090
rect 20108 3050 20118 3090
rect 20058 3030 20118 3050
rect 20228 3090 20288 3110
rect 20228 3050 20238 3090
rect 20278 3050 20288 3090
rect 20328 3090 20428 3110
rect 20328 3050 20378 3090
rect 20418 3050 20428 3090
rect 20228 3030 20288 3050
rect 20368 3030 20428 3050
rect 20478 3090 20538 3110
rect 20478 3050 20488 3090
rect 20528 3050 20538 3090
rect 20478 3030 20538 3050
rect 20588 3090 20648 3110
rect 20588 3050 20598 3090
rect 20638 3050 20648 3090
rect 20588 3030 20648 3050
rect 20698 3090 20758 3110
rect 20698 3050 20708 3090
rect 20748 3050 20758 3090
rect 20698 3030 20758 3050
rect 20808 3090 20868 3110
rect 20808 3050 20818 3090
rect 20858 3050 20868 3090
rect 20908 3090 21088 3110
rect 20908 3070 21038 3090
rect 20808 3030 20868 3050
rect 21028 3050 21038 3070
rect 21078 3050 21088 3090
rect 21028 3030 21088 3050
rect 21138 3090 21198 3110
rect 21138 3050 21148 3090
rect 21188 3050 21198 3090
rect 21138 3030 21198 3050
rect 21248 3090 21308 3110
rect 21248 3050 21258 3090
rect 21298 3050 21308 3090
rect 21248 3030 21308 3050
rect 21358 3090 21418 3110
rect 21358 3050 21368 3090
rect 21408 3050 21418 3090
rect 21358 3030 21418 3050
rect 21528 3090 21588 3110
rect 21528 3050 21538 3090
rect 21578 3050 21588 3090
rect 21628 3090 21728 3110
rect 21628 3050 21678 3090
rect 21718 3050 21728 3090
rect 21528 3030 21588 3050
rect 21668 3030 21728 3050
rect 21778 3090 21838 3110
rect 21778 3050 21788 3090
rect 21828 3050 21838 3090
rect 21778 3030 21838 3050
rect 21888 3090 21948 3110
rect 21888 3050 21898 3090
rect 21938 3050 21948 3090
rect 21888 3030 21948 3050
rect 21998 3090 22058 3110
rect 21998 3050 22008 3090
rect 22048 3050 22058 3090
rect 21998 3030 22058 3050
rect 22108 3090 22168 3110
rect 22108 3050 22118 3090
rect 22158 3050 22168 3090
rect 22208 3090 22388 3110
rect 22208 3070 22338 3090
rect 22108 3030 22168 3050
rect 22328 3050 22338 3070
rect 22378 3050 22388 3090
rect 22328 3030 22388 3050
rect 22438 3090 22498 3110
rect 22438 3050 22448 3090
rect 22488 3050 22498 3090
rect 22438 3030 22498 3050
rect 22548 3090 22608 3110
rect 22548 3050 22558 3090
rect 22598 3050 22608 3090
rect 22548 3030 22608 3050
rect 22658 3090 22718 3110
rect 22658 3050 22668 3090
rect 22708 3050 22718 3090
rect 22658 3030 22718 3050
rect 18938 2970 18978 3030
rect 19188 2970 19228 3030
rect 19408 2970 19448 3030
rect 19958 2970 19998 3030
rect 20238 2970 20278 3030
rect 20488 2970 20528 3030
rect 20708 2970 20748 3030
rect 21258 2970 21298 3030
rect 21538 2970 21578 3030
rect 21788 2970 21828 3030
rect 22008 2970 22048 3030
rect 22558 2970 22598 3030
rect 12538 2950 12618 2970
rect 12538 2910 12558 2950
rect 12598 2910 12618 2950
rect 12538 2890 12618 2910
rect 12758 2950 12838 2970
rect 12758 2910 12778 2950
rect 12818 2910 12838 2950
rect 12758 2890 12838 2910
rect 13228 2950 13308 2970
rect 13228 2910 13248 2950
rect 13288 2910 13308 2950
rect 13228 2890 13308 2910
rect 13568 2950 13648 2970
rect 13568 2910 13588 2950
rect 13628 2910 13648 2950
rect 13568 2890 13648 2910
rect 13788 2950 13868 2970
rect 13788 2910 13808 2950
rect 13848 2910 13868 2950
rect 13788 2890 13868 2910
rect 14228 2950 14308 2970
rect 14228 2910 14248 2950
rect 14288 2910 14308 2950
rect 14228 2890 14308 2910
rect 14908 2950 14988 2970
rect 14908 2910 14928 2950
rect 14968 2910 14988 2950
rect 14908 2890 14988 2910
rect 15128 2950 15208 2970
rect 15128 2910 15148 2950
rect 15188 2910 15208 2950
rect 15128 2890 15208 2910
rect 15598 2950 15678 2970
rect 15598 2910 15618 2950
rect 15658 2910 15678 2950
rect 15598 2890 15678 2910
rect 16058 2950 16138 2970
rect 16058 2910 16078 2950
rect 16118 2910 16138 2950
rect 16058 2890 16138 2910
rect 16408 2950 16488 2970
rect 16408 2910 16428 2950
rect 16468 2910 16488 2950
rect 16408 2890 16488 2910
rect 16658 2950 16738 2970
rect 16658 2910 16678 2950
rect 16718 2910 16738 2950
rect 16658 2890 16738 2910
rect 16878 2950 16958 2970
rect 16878 2910 16898 2950
rect 16938 2910 16958 2950
rect 16878 2890 16958 2910
rect 17208 2950 17288 2970
rect 17208 2910 17228 2950
rect 17268 2910 17288 2950
rect 17208 2890 17288 2910
rect 17868 2950 17948 2970
rect 17868 2910 17888 2950
rect 17928 2910 17948 2950
rect 17868 2890 17948 2910
rect 18088 2950 18168 2970
rect 18088 2910 18108 2950
rect 18148 2910 18168 2950
rect 18088 2890 18168 2910
rect 18658 2950 18738 2970
rect 18658 2910 18678 2950
rect 18718 2910 18738 2950
rect 18658 2890 18738 2910
rect 18918 2950 18998 2970
rect 18918 2910 18938 2950
rect 18978 2910 18998 2950
rect 18918 2890 18998 2910
rect 19168 2950 19248 2970
rect 19168 2910 19188 2950
rect 19228 2910 19248 2950
rect 19168 2890 19248 2910
rect 19388 2950 19468 2970
rect 19388 2910 19408 2950
rect 19448 2910 19468 2950
rect 19388 2890 19468 2910
rect 19938 2950 20018 2970
rect 19938 2910 19958 2950
rect 19998 2910 20018 2950
rect 19938 2890 20018 2910
rect 20218 2950 20298 2970
rect 20218 2910 20238 2950
rect 20278 2910 20298 2950
rect 20218 2890 20298 2910
rect 20468 2950 20548 2970
rect 20468 2910 20488 2950
rect 20528 2910 20548 2950
rect 20468 2890 20548 2910
rect 20688 2950 20768 2970
rect 20688 2910 20708 2950
rect 20748 2910 20768 2950
rect 20688 2890 20768 2910
rect 21238 2950 21318 2970
rect 21238 2910 21258 2950
rect 21298 2910 21318 2950
rect 21238 2890 21318 2910
rect 21518 2950 21598 2970
rect 21518 2910 21538 2950
rect 21578 2910 21598 2950
rect 21518 2890 21598 2910
rect 21768 2950 21848 2970
rect 21768 2910 21788 2950
rect 21828 2910 21848 2950
rect 21768 2890 21848 2910
rect 21988 2950 22068 2970
rect 21988 2910 22008 2950
rect 22048 2910 22068 2950
rect 21988 2890 22068 2910
rect 22538 2950 22618 2970
rect 22538 2910 22558 2950
rect 22598 2910 22618 2950
rect 22538 2890 22618 2910
rect 23088 2660 23128 3180
rect 23250 3122 23308 3140
rect 23250 3088 23262 3122
rect 23296 3088 23308 3122
rect 23250 3070 23308 3088
rect 23770 3122 23828 3140
rect 23770 3088 23782 3122
rect 23816 3088 23828 3122
rect 23770 3070 23828 3088
rect 24290 3122 24348 3140
rect 24290 3088 24302 3122
rect 24336 3088 24348 3122
rect 24290 3070 24348 3088
rect 23206 3010 23266 3030
rect 23206 2970 23216 3010
rect 23256 2970 23266 3010
rect 23206 2910 23266 2970
rect 23206 2870 23216 2910
rect 23256 2870 23266 2910
rect 23206 2850 23266 2870
rect 23318 3010 23378 3030
rect 23318 2970 23328 3010
rect 23368 2970 23378 3010
rect 23318 2910 23378 2970
rect 23318 2870 23328 2910
rect 23368 2870 23378 2910
rect 23318 2850 23378 2870
rect 23726 3010 23786 3030
rect 23726 2970 23736 3010
rect 23776 2970 23786 3010
rect 23726 2910 23786 2970
rect 23726 2870 23736 2910
rect 23776 2870 23786 2910
rect 23726 2850 23786 2870
rect 23838 3010 23898 3030
rect 23838 2970 23848 3010
rect 23888 2970 23898 3010
rect 23838 2910 23898 2970
rect 23838 2870 23848 2910
rect 23888 2870 23898 2910
rect 23838 2850 23898 2870
rect 24246 3010 24306 3030
rect 24246 2970 24256 3010
rect 24296 2970 24306 3010
rect 24246 2910 24306 2970
rect 24246 2870 24256 2910
rect 24296 2870 24306 2910
rect 24246 2850 24306 2870
rect 24358 3010 24418 3030
rect 24358 2970 24368 3010
rect 24408 2970 24418 3010
rect 24358 2910 24418 2970
rect 24358 2870 24368 2910
rect 24408 2870 24418 2910
rect 24358 2850 24418 2870
rect 23278 2742 23336 2760
rect 23278 2708 23290 2742
rect 23324 2708 23336 2742
rect 23278 2690 23336 2708
rect 23798 2742 23856 2760
rect 23798 2708 23810 2742
rect 23844 2708 23856 2742
rect 23798 2690 23856 2708
rect 24318 2742 24376 2760
rect 24318 2708 24330 2742
rect 24364 2708 24376 2742
rect 24318 2690 24376 2708
rect 25088 2660 25128 3180
rect 23088 1920 23128 2450
rect 23208 2630 23268 2650
rect 23208 2590 23218 2630
rect 23258 2590 23268 2630
rect 23208 2530 23268 2590
rect 23208 2490 23218 2530
rect 23258 2490 23268 2530
rect 23208 2430 23268 2490
rect 23208 2390 23218 2430
rect 23258 2390 23268 2430
rect 23208 2370 23268 2390
rect 23318 2630 23378 2650
rect 23318 2590 23328 2630
rect 23368 2590 23378 2630
rect 23318 2530 23378 2590
rect 23318 2490 23328 2530
rect 23368 2490 23378 2530
rect 23318 2430 23378 2490
rect 23318 2390 23328 2430
rect 23368 2390 23378 2430
rect 23318 2370 23378 2390
rect 23728 2630 23788 2650
rect 23728 2590 23738 2630
rect 23778 2590 23788 2630
rect 23728 2530 23788 2590
rect 23728 2490 23738 2530
rect 23778 2490 23788 2530
rect 23728 2430 23788 2490
rect 23728 2390 23738 2430
rect 23778 2390 23788 2430
rect 23728 2370 23788 2390
rect 23838 2630 23898 2650
rect 23838 2590 23848 2630
rect 23888 2590 23898 2630
rect 23838 2530 23898 2590
rect 23838 2490 23848 2530
rect 23888 2490 23898 2530
rect 23838 2430 23898 2490
rect 23838 2390 23848 2430
rect 23888 2390 23898 2430
rect 23838 2370 23898 2390
rect 24248 2630 24308 2650
rect 24248 2590 24258 2630
rect 24298 2590 24308 2630
rect 24248 2530 24308 2590
rect 24248 2490 24258 2530
rect 24298 2490 24308 2530
rect 24248 2430 24308 2490
rect 24248 2390 24258 2430
rect 24298 2390 24308 2430
rect 24248 2370 24308 2390
rect 24358 2630 24418 2650
rect 24358 2590 24368 2630
rect 24408 2590 24418 2630
rect 24358 2530 24418 2590
rect 24358 2490 24368 2530
rect 24408 2490 24418 2530
rect 24358 2430 24418 2490
rect 24358 2390 24368 2430
rect 24408 2390 24418 2430
rect 24358 2370 24418 2390
rect 23264 2262 23322 2280
rect 23264 2228 23276 2262
rect 23310 2228 23322 2262
rect 23264 2210 23322 2228
rect 23784 2262 23842 2280
rect 23784 2228 23796 2262
rect 23830 2228 23842 2262
rect 23784 2210 23842 2228
rect 24304 2262 24362 2280
rect 24304 2228 24316 2262
rect 24350 2228 24362 2262
rect 24304 2210 24362 2228
rect 24872 2262 24930 2280
rect 24872 2228 24884 2262
rect 24918 2228 24930 2262
rect 24872 2210 24930 2228
rect 23208 2150 23268 2170
rect 23208 2110 23218 2150
rect 23258 2110 23268 2150
rect 23208 2050 23268 2110
rect 23208 2010 23218 2050
rect 23258 2010 23268 2050
rect 23208 1990 23268 2010
rect 23318 2150 23378 2170
rect 23318 2110 23328 2150
rect 23368 2110 23378 2150
rect 23318 2050 23378 2110
rect 23318 2010 23328 2050
rect 23368 2010 23378 2050
rect 23318 1990 23378 2010
rect 23728 2150 23788 2170
rect 23728 2110 23738 2150
rect 23778 2110 23788 2150
rect 23728 2050 23788 2110
rect 23728 2010 23738 2050
rect 23778 2010 23788 2050
rect 23728 1990 23788 2010
rect 23838 2150 23898 2170
rect 23838 2110 23848 2150
rect 23888 2110 23898 2150
rect 23838 2050 23898 2110
rect 23838 2010 23848 2050
rect 23888 2010 23898 2050
rect 23838 1990 23898 2010
rect 24248 2150 24308 2170
rect 24248 2110 24258 2150
rect 24298 2110 24308 2150
rect 24248 2050 24308 2110
rect 24248 2010 24258 2050
rect 24298 2010 24308 2050
rect 24248 1990 24308 2010
rect 24358 2150 24418 2170
rect 24358 2110 24368 2150
rect 24408 2110 24418 2150
rect 24358 2050 24418 2110
rect 24358 2010 24368 2050
rect 24408 2010 24418 2050
rect 24358 1990 24418 2010
rect 24848 2150 24908 2170
rect 24848 2110 24858 2150
rect 24898 2110 24908 2150
rect 24848 2050 24908 2110
rect 24848 2010 24858 2050
rect 24898 2010 24908 2050
rect 24848 1990 24908 2010
rect 24958 2150 25018 2170
rect 24958 2110 24968 2150
rect 25008 2110 25018 2150
rect 24958 2050 25018 2110
rect 24958 2010 24968 2050
rect 25008 2010 25018 2050
rect 24958 1990 25018 2010
rect 23308 1920 23388 1940
rect 23828 1920 23908 1940
rect 24348 1920 24428 1940
rect 24838 1920 24918 1940
rect 25088 1920 25128 2450
rect 23088 1880 23328 1920
rect 23368 1880 23848 1920
rect 23888 1880 24228 1920
rect 24408 1880 24858 1920
rect 24898 1880 25128 1920
rect 23308 1860 23388 1880
rect 23828 1860 23908 1880
rect 24348 1860 24428 1880
rect 24838 1860 24918 1880
<< viali >>
rect 16138 19663 16178 19680
rect 16138 19640 16178 19663
rect 15008 19452 15405 19490
rect 16911 19452 17308 19490
rect 13258 19030 13298 19070
rect 13258 18950 13298 18990
rect 13258 18870 13298 18910
rect 8468 18597 8508 18610
rect 9258 18600 9298 18610
rect 8468 18570 8508 18597
rect 8468 18043 8506 18440
rect 8468 17234 8506 17631
rect 9258 18570 9298 18600
rect 10698 18597 10738 18610
rect 9248 18060 9288 18450
rect 9588 16836 9628 17226
rect 10698 18570 10738 18597
rect 10698 18050 10738 18440
rect 10368 16310 10408 16700
rect 11658 18392 11664 18414
rect 11664 18392 11692 18414
rect 11658 18380 11692 18392
rect 11758 18380 11792 18414
rect 11858 18380 11892 18414
rect 11958 18392 11990 18414
rect 11990 18392 11992 18414
rect 12058 18392 12080 18414
rect 12080 18392 12092 18414
rect 12158 18392 12170 18414
rect 12170 18392 12192 18414
rect 11958 18380 11992 18392
rect 12058 18380 12092 18392
rect 12158 18380 12192 18392
rect 11658 18302 11664 18314
rect 11664 18302 11692 18314
rect 11658 18280 11692 18302
rect 11758 18280 11792 18314
rect 11858 18280 11892 18314
rect 11958 18302 11990 18314
rect 11990 18302 11992 18314
rect 12058 18302 12080 18314
rect 12080 18302 12092 18314
rect 12158 18302 12170 18314
rect 12170 18302 12192 18314
rect 11958 18280 11992 18302
rect 12058 18280 12092 18302
rect 12158 18280 12192 18302
rect 11658 18212 11664 18214
rect 11664 18212 11692 18214
rect 11658 18180 11692 18212
rect 11758 18180 11792 18214
rect 11858 18180 11892 18214
rect 11958 18212 11990 18214
rect 11990 18212 11992 18214
rect 12058 18212 12080 18214
rect 12080 18212 12092 18214
rect 12158 18212 12170 18214
rect 12170 18212 12192 18214
rect 11958 18180 11992 18212
rect 12058 18180 12092 18212
rect 12158 18180 12192 18212
rect 11658 18080 11692 18114
rect 11758 18080 11792 18114
rect 11858 18080 11892 18114
rect 11958 18080 11992 18114
rect 12058 18080 12092 18114
rect 12158 18080 12192 18114
rect 11658 17980 11692 18014
rect 11758 17980 11792 18014
rect 11858 17980 11892 18014
rect 11958 17980 11992 18014
rect 12058 17980 12092 18014
rect 12158 17980 12192 18014
rect 11658 17886 11692 17914
rect 11658 17880 11664 17886
rect 11664 17880 11692 17886
rect 11758 17880 11792 17914
rect 11858 17880 11892 17914
rect 11958 17886 11992 17914
rect 12058 17886 12092 17914
rect 12158 17886 12192 17914
rect 11958 17880 11990 17886
rect 11990 17880 11992 17886
rect 12058 17880 12080 17886
rect 12080 17880 12092 17886
rect 12158 17880 12170 17886
rect 12170 17880 12192 17886
rect 13018 18392 13024 18414
rect 13024 18392 13052 18414
rect 13018 18380 13052 18392
rect 13118 18380 13152 18414
rect 13218 18380 13252 18414
rect 13318 18392 13350 18414
rect 13350 18392 13352 18414
rect 13418 18392 13440 18414
rect 13440 18392 13452 18414
rect 13518 18392 13530 18414
rect 13530 18392 13552 18414
rect 13318 18380 13352 18392
rect 13418 18380 13452 18392
rect 13518 18380 13552 18392
rect 13018 18302 13024 18314
rect 13024 18302 13052 18314
rect 13018 18280 13052 18302
rect 13118 18280 13152 18314
rect 13218 18280 13252 18314
rect 13318 18302 13350 18314
rect 13350 18302 13352 18314
rect 13418 18302 13440 18314
rect 13440 18302 13452 18314
rect 13518 18302 13530 18314
rect 13530 18302 13552 18314
rect 13318 18280 13352 18302
rect 13418 18280 13452 18302
rect 13518 18280 13552 18302
rect 13018 18212 13024 18214
rect 13024 18212 13052 18214
rect 13018 18180 13052 18212
rect 13118 18180 13152 18214
rect 13218 18180 13252 18214
rect 13318 18212 13350 18214
rect 13350 18212 13352 18214
rect 13418 18212 13440 18214
rect 13440 18212 13452 18214
rect 13518 18212 13530 18214
rect 13530 18212 13552 18214
rect 13318 18180 13352 18212
rect 13418 18180 13452 18212
rect 13518 18180 13552 18212
rect 13018 18080 13052 18114
rect 13118 18080 13152 18114
rect 13218 18080 13252 18114
rect 13318 18080 13352 18114
rect 13418 18080 13452 18114
rect 13518 18080 13552 18114
rect 13018 17980 13052 18014
rect 13118 17980 13152 18014
rect 13218 17980 13252 18014
rect 13318 17980 13352 18014
rect 13418 17980 13452 18014
rect 13518 17980 13552 18014
rect 13018 17886 13052 17914
rect 13018 17880 13024 17886
rect 13024 17880 13052 17886
rect 13118 17880 13152 17914
rect 13218 17880 13252 17914
rect 13318 17886 13352 17914
rect 13418 17886 13452 17914
rect 13518 17886 13552 17914
rect 13318 17880 13350 17886
rect 13350 17880 13352 17886
rect 13418 17880 13440 17886
rect 13440 17880 13452 17886
rect 13518 17880 13530 17886
rect 13530 17880 13552 17886
rect 14378 18392 14384 18414
rect 14384 18392 14412 18414
rect 14378 18380 14412 18392
rect 14478 18380 14512 18414
rect 14578 18380 14612 18414
rect 14678 18392 14710 18414
rect 14710 18392 14712 18414
rect 14778 18392 14800 18414
rect 14800 18392 14812 18414
rect 14878 18392 14890 18414
rect 14890 18392 14912 18414
rect 14678 18380 14712 18392
rect 14778 18380 14812 18392
rect 14878 18380 14912 18392
rect 14378 18302 14384 18314
rect 14384 18302 14412 18314
rect 14378 18280 14412 18302
rect 14478 18280 14512 18314
rect 14578 18280 14612 18314
rect 14678 18302 14710 18314
rect 14710 18302 14712 18314
rect 14778 18302 14800 18314
rect 14800 18302 14812 18314
rect 14878 18302 14890 18314
rect 14890 18302 14912 18314
rect 14678 18280 14712 18302
rect 14778 18280 14812 18302
rect 14878 18280 14912 18302
rect 14378 18212 14384 18214
rect 14384 18212 14412 18214
rect 14378 18180 14412 18212
rect 14478 18180 14512 18214
rect 14578 18180 14612 18214
rect 14678 18212 14710 18214
rect 14710 18212 14712 18214
rect 14778 18212 14800 18214
rect 14800 18212 14812 18214
rect 14878 18212 14890 18214
rect 14890 18212 14912 18214
rect 14678 18180 14712 18212
rect 14778 18180 14812 18212
rect 14878 18180 14912 18212
rect 14378 18080 14412 18114
rect 14478 18080 14512 18114
rect 14578 18080 14612 18114
rect 14678 18080 14712 18114
rect 14778 18080 14812 18114
rect 14878 18080 14912 18114
rect 14378 17980 14412 18014
rect 14478 17980 14512 18014
rect 14578 17980 14612 18014
rect 14678 17980 14712 18014
rect 14778 17980 14812 18014
rect 14878 17980 14912 18014
rect 14378 17886 14412 17914
rect 14378 17880 14384 17886
rect 14384 17880 14412 17886
rect 14478 17880 14512 17914
rect 14578 17880 14612 17914
rect 14678 17886 14712 17914
rect 14778 17886 14812 17914
rect 14878 17886 14912 17914
rect 14678 17880 14710 17886
rect 14710 17880 14712 17886
rect 14778 17880 14800 17886
rect 14800 17880 14812 17886
rect 14878 17880 14890 17886
rect 14890 17880 14912 17886
rect 15688 18597 15728 18610
rect 15688 18570 15728 18597
rect 16798 18594 16838 18610
rect 17588 18597 17628 18610
rect 11658 17032 11664 17054
rect 11664 17032 11692 17054
rect 11658 17020 11692 17032
rect 11758 17020 11792 17054
rect 11858 17020 11892 17054
rect 11958 17032 11990 17054
rect 11990 17032 11992 17054
rect 12058 17032 12080 17054
rect 12080 17032 12092 17054
rect 12158 17032 12170 17054
rect 12170 17032 12192 17054
rect 11958 17020 11992 17032
rect 12058 17020 12092 17032
rect 12158 17020 12192 17032
rect 11658 16942 11664 16954
rect 11664 16942 11692 16954
rect 11658 16920 11692 16942
rect 11758 16920 11792 16954
rect 11858 16920 11892 16954
rect 11958 16942 11990 16954
rect 11990 16942 11992 16954
rect 12058 16942 12080 16954
rect 12080 16942 12092 16954
rect 12158 16942 12170 16954
rect 12170 16942 12192 16954
rect 11958 16920 11992 16942
rect 12058 16920 12092 16942
rect 12158 16920 12192 16942
rect 11658 16852 11664 16854
rect 11664 16852 11692 16854
rect 11658 16820 11692 16852
rect 11758 16820 11792 16854
rect 11858 16820 11892 16854
rect 11958 16852 11990 16854
rect 11990 16852 11992 16854
rect 12058 16852 12080 16854
rect 12080 16852 12092 16854
rect 12158 16852 12170 16854
rect 12170 16852 12192 16854
rect 11958 16820 11992 16852
rect 12058 16820 12092 16852
rect 12158 16820 12192 16852
rect 11658 16720 11692 16754
rect 11758 16720 11792 16754
rect 11858 16720 11892 16754
rect 11958 16720 11992 16754
rect 12058 16720 12092 16754
rect 12158 16720 12192 16754
rect 11658 16620 11692 16654
rect 11758 16620 11792 16654
rect 11858 16620 11892 16654
rect 11958 16620 11992 16654
rect 12058 16620 12092 16654
rect 12158 16620 12192 16654
rect 11658 16526 11692 16554
rect 11658 16520 11664 16526
rect 11664 16520 11692 16526
rect 11758 16520 11792 16554
rect 11858 16520 11892 16554
rect 11958 16526 11992 16554
rect 12058 16526 12092 16554
rect 12158 16526 12192 16554
rect 11958 16520 11990 16526
rect 11990 16520 11992 16526
rect 12058 16520 12080 16526
rect 12080 16520 12092 16526
rect 12158 16520 12170 16526
rect 12170 16520 12192 16526
rect 13018 17032 13024 17054
rect 13024 17032 13052 17054
rect 13018 17020 13052 17032
rect 13118 17020 13152 17054
rect 13218 17020 13252 17054
rect 13318 17032 13350 17054
rect 13350 17032 13352 17054
rect 13418 17032 13440 17054
rect 13440 17032 13452 17054
rect 13518 17032 13530 17054
rect 13530 17032 13552 17054
rect 13318 17020 13352 17032
rect 13418 17020 13452 17032
rect 13518 17020 13552 17032
rect 13018 16942 13024 16954
rect 13024 16942 13052 16954
rect 13018 16920 13052 16942
rect 13118 16920 13152 16954
rect 13218 16920 13252 16954
rect 13318 16942 13350 16954
rect 13350 16942 13352 16954
rect 13418 16942 13440 16954
rect 13440 16942 13452 16954
rect 13518 16942 13530 16954
rect 13530 16942 13552 16954
rect 13318 16920 13352 16942
rect 13418 16920 13452 16942
rect 13518 16920 13552 16942
rect 13018 16852 13024 16854
rect 13024 16852 13052 16854
rect 13018 16820 13052 16852
rect 13118 16820 13152 16854
rect 13218 16820 13252 16854
rect 13318 16852 13350 16854
rect 13350 16852 13352 16854
rect 13418 16852 13440 16854
rect 13440 16852 13452 16854
rect 13518 16852 13530 16854
rect 13530 16852 13552 16854
rect 13318 16820 13352 16852
rect 13418 16820 13452 16852
rect 13518 16820 13552 16852
rect 13018 16720 13052 16754
rect 13118 16720 13152 16754
rect 13218 16720 13252 16754
rect 13318 16720 13352 16754
rect 13418 16720 13452 16754
rect 13518 16720 13552 16754
rect 13018 16620 13052 16654
rect 13118 16620 13152 16654
rect 13218 16620 13252 16654
rect 13318 16620 13352 16654
rect 13418 16620 13452 16654
rect 13518 16620 13552 16654
rect 13018 16526 13052 16554
rect 13018 16520 13024 16526
rect 13024 16520 13052 16526
rect 13118 16520 13152 16554
rect 13218 16520 13252 16554
rect 13318 16526 13352 16554
rect 13418 16526 13452 16554
rect 13518 16526 13552 16554
rect 13318 16520 13350 16526
rect 13350 16520 13352 16526
rect 13418 16520 13440 16526
rect 13440 16520 13452 16526
rect 13518 16520 13530 16526
rect 13530 16520 13552 16526
rect 14378 17032 14384 17054
rect 14384 17032 14412 17054
rect 14378 17020 14412 17032
rect 14478 17020 14512 17054
rect 14578 17020 14612 17054
rect 14678 17032 14710 17054
rect 14710 17032 14712 17054
rect 14778 17032 14800 17054
rect 14800 17032 14812 17054
rect 14878 17032 14890 17054
rect 14890 17032 14912 17054
rect 14678 17020 14712 17032
rect 14778 17020 14812 17032
rect 14878 17020 14912 17032
rect 14378 16942 14384 16954
rect 14384 16942 14412 16954
rect 14378 16920 14412 16942
rect 14478 16920 14512 16954
rect 14578 16920 14612 16954
rect 14678 16942 14710 16954
rect 14710 16942 14712 16954
rect 14778 16942 14800 16954
rect 14800 16942 14812 16954
rect 14878 16942 14890 16954
rect 14890 16942 14912 16954
rect 14678 16920 14712 16942
rect 14778 16920 14812 16942
rect 14878 16920 14912 16942
rect 14378 16852 14384 16854
rect 14384 16852 14412 16854
rect 14378 16820 14412 16852
rect 14478 16820 14512 16854
rect 14578 16820 14612 16854
rect 14678 16852 14710 16854
rect 14710 16852 14712 16854
rect 14778 16852 14800 16854
rect 14800 16852 14812 16854
rect 14878 16852 14890 16854
rect 14890 16852 14912 16854
rect 14678 16820 14712 16852
rect 14778 16820 14812 16852
rect 14878 16820 14912 16852
rect 14378 16720 14412 16754
rect 14478 16720 14512 16754
rect 14578 16720 14612 16754
rect 14678 16720 14712 16754
rect 14778 16720 14812 16754
rect 14878 16720 14912 16754
rect 14378 16620 14412 16654
rect 14478 16620 14512 16654
rect 14578 16620 14612 16654
rect 14678 16620 14712 16654
rect 14778 16620 14812 16654
rect 14878 16620 14912 16654
rect 14378 16526 14412 16554
rect 14378 16520 14384 16526
rect 14384 16520 14412 16526
rect 14478 16520 14512 16554
rect 14578 16520 14612 16554
rect 14678 16526 14712 16554
rect 14778 16526 14812 16554
rect 14878 16526 14912 16554
rect 14678 16520 14710 16526
rect 14710 16520 14712 16526
rect 14778 16520 14800 16526
rect 14800 16520 14812 16526
rect 14878 16520 14890 16526
rect 14890 16520 14912 16526
rect 15688 18050 15728 18440
rect 16018 16310 16058 16700
rect 16798 18570 16838 18594
rect 16801 18040 16839 18437
rect 16801 17441 16839 17838
rect 17588 18570 17628 18597
rect 17588 18043 17626 18440
rect 17588 17234 17626 17631
rect 11658 15672 11664 15694
rect 11664 15672 11692 15694
rect 11658 15660 11692 15672
rect 11758 15660 11792 15694
rect 11858 15660 11892 15694
rect 11958 15672 11990 15694
rect 11990 15672 11992 15694
rect 12058 15672 12080 15694
rect 12080 15672 12092 15694
rect 12158 15672 12170 15694
rect 12170 15672 12192 15694
rect 11958 15660 11992 15672
rect 12058 15660 12092 15672
rect 12158 15660 12192 15672
rect 11658 15582 11664 15594
rect 11664 15582 11692 15594
rect 11658 15560 11692 15582
rect 11758 15560 11792 15594
rect 11858 15560 11892 15594
rect 11958 15582 11990 15594
rect 11990 15582 11992 15594
rect 12058 15582 12080 15594
rect 12080 15582 12092 15594
rect 12158 15582 12170 15594
rect 12170 15582 12192 15594
rect 11958 15560 11992 15582
rect 12058 15560 12092 15582
rect 12158 15560 12192 15582
rect 11658 15492 11664 15494
rect 11664 15492 11692 15494
rect 11658 15460 11692 15492
rect 11758 15460 11792 15494
rect 11858 15460 11892 15494
rect 11958 15492 11990 15494
rect 11990 15492 11992 15494
rect 12058 15492 12080 15494
rect 12080 15492 12092 15494
rect 12158 15492 12170 15494
rect 12170 15492 12192 15494
rect 11958 15460 11992 15492
rect 12058 15460 12092 15492
rect 12158 15460 12192 15492
rect 11658 15360 11692 15394
rect 11758 15360 11792 15394
rect 11858 15360 11892 15394
rect 11958 15360 11992 15394
rect 12058 15360 12092 15394
rect 12158 15360 12192 15394
rect 11658 15260 11692 15294
rect 11758 15260 11792 15294
rect 11858 15260 11892 15294
rect 11958 15260 11992 15294
rect 12058 15260 12092 15294
rect 12158 15260 12192 15294
rect 11658 15166 11692 15194
rect 11658 15160 11664 15166
rect 11664 15160 11692 15166
rect 11758 15160 11792 15194
rect 11858 15160 11892 15194
rect 11958 15166 11992 15194
rect 12058 15166 12092 15194
rect 12158 15166 12192 15194
rect 11958 15160 11990 15166
rect 11990 15160 11992 15166
rect 12058 15160 12080 15166
rect 12080 15160 12092 15166
rect 12158 15160 12170 15166
rect 12170 15160 12192 15166
rect 13018 15672 13024 15694
rect 13024 15672 13052 15694
rect 13018 15660 13052 15672
rect 13118 15660 13152 15694
rect 13218 15660 13252 15694
rect 13318 15672 13350 15694
rect 13350 15672 13352 15694
rect 13418 15672 13440 15694
rect 13440 15672 13452 15694
rect 13518 15672 13530 15694
rect 13530 15672 13552 15694
rect 13318 15660 13352 15672
rect 13418 15660 13452 15672
rect 13518 15660 13552 15672
rect 13018 15582 13024 15594
rect 13024 15582 13052 15594
rect 13018 15560 13052 15582
rect 13118 15560 13152 15594
rect 13218 15560 13252 15594
rect 13318 15582 13350 15594
rect 13350 15582 13352 15594
rect 13418 15582 13440 15594
rect 13440 15582 13452 15594
rect 13518 15582 13530 15594
rect 13530 15582 13552 15594
rect 13318 15560 13352 15582
rect 13418 15560 13452 15582
rect 13518 15560 13552 15582
rect 13018 15492 13024 15494
rect 13024 15492 13052 15494
rect 13018 15460 13052 15492
rect 13118 15460 13152 15494
rect 13218 15460 13252 15494
rect 13318 15492 13350 15494
rect 13350 15492 13352 15494
rect 13418 15492 13440 15494
rect 13440 15492 13452 15494
rect 13518 15492 13530 15494
rect 13530 15492 13552 15494
rect 13318 15460 13352 15492
rect 13418 15460 13452 15492
rect 13518 15460 13552 15492
rect 13018 15360 13052 15394
rect 13118 15360 13152 15394
rect 13218 15360 13252 15394
rect 13318 15360 13352 15394
rect 13418 15360 13452 15394
rect 13518 15360 13552 15394
rect 13018 15260 13052 15294
rect 13118 15260 13152 15294
rect 13218 15260 13252 15294
rect 13318 15260 13352 15294
rect 13418 15260 13452 15294
rect 13518 15260 13552 15294
rect 13018 15166 13052 15194
rect 13018 15160 13024 15166
rect 13024 15160 13052 15166
rect 13118 15160 13152 15194
rect 13218 15160 13252 15194
rect 13318 15166 13352 15194
rect 13418 15166 13452 15194
rect 13518 15166 13552 15194
rect 13318 15160 13350 15166
rect 13350 15160 13352 15166
rect 13418 15160 13440 15166
rect 13440 15160 13452 15166
rect 13518 15160 13530 15166
rect 13530 15160 13552 15166
rect 14378 15672 14384 15694
rect 14384 15672 14412 15694
rect 14378 15660 14412 15672
rect 14478 15660 14512 15694
rect 14578 15660 14612 15694
rect 14678 15672 14710 15694
rect 14710 15672 14712 15694
rect 14778 15672 14800 15694
rect 14800 15672 14812 15694
rect 14878 15672 14890 15694
rect 14890 15672 14912 15694
rect 14678 15660 14712 15672
rect 14778 15660 14812 15672
rect 14878 15660 14912 15672
rect 14378 15582 14384 15594
rect 14384 15582 14412 15594
rect 14378 15560 14412 15582
rect 14478 15560 14512 15594
rect 14578 15560 14612 15594
rect 14678 15582 14710 15594
rect 14710 15582 14712 15594
rect 14778 15582 14800 15594
rect 14800 15582 14812 15594
rect 14878 15582 14890 15594
rect 14890 15582 14912 15594
rect 14678 15560 14712 15582
rect 14778 15560 14812 15582
rect 14878 15560 14912 15582
rect 14378 15492 14384 15494
rect 14384 15492 14412 15494
rect 14378 15460 14412 15492
rect 14478 15460 14512 15494
rect 14578 15460 14612 15494
rect 14678 15492 14710 15494
rect 14710 15492 14712 15494
rect 14778 15492 14800 15494
rect 14800 15492 14812 15494
rect 14878 15492 14890 15494
rect 14890 15492 14912 15494
rect 14678 15460 14712 15492
rect 14778 15460 14812 15492
rect 14878 15460 14912 15492
rect 14378 15360 14412 15394
rect 14478 15360 14512 15394
rect 14578 15360 14612 15394
rect 14678 15360 14712 15394
rect 14778 15360 14812 15394
rect 14878 15360 14912 15394
rect 14378 15260 14412 15294
rect 14478 15260 14512 15294
rect 14578 15260 14612 15294
rect 14678 15260 14712 15294
rect 14778 15260 14812 15294
rect 14878 15260 14912 15294
rect 14378 15166 14412 15194
rect 14378 15160 14384 15166
rect 14384 15160 14412 15166
rect 14478 15160 14512 15194
rect 14578 15160 14612 15194
rect 14678 15166 14712 15194
rect 14778 15166 14812 15194
rect 14878 15166 14912 15194
rect 14678 15160 14710 15166
rect 14710 15160 14712 15166
rect 14778 15160 14800 15166
rect 14800 15160 14812 15166
rect 14878 15160 14890 15166
rect 14890 15160 14912 15166
rect 12560 14550 12610 14600
rect 13958 14550 14008 14600
rect 11098 14160 11138 14200
rect 15488 14200 15528 14240
rect 15488 14120 15528 14160
rect 11178 13990 11218 14030
rect 11338 13990 11378 14030
rect 11498 13990 11538 14030
rect 11658 13990 11698 14030
rect 11818 13990 11858 14030
rect 11978 13990 12018 14030
rect 12138 13990 12178 14030
rect 12298 13990 12338 14030
rect 12458 13990 12498 14030
rect 12618 13990 12658 14030
rect 12778 13990 12818 14030
rect 12938 13990 12978 14030
rect 13098 13990 13138 14030
rect 13258 13990 13298 14030
rect 13418 13990 13458 14030
rect 13578 13990 13618 14030
rect 13738 13990 13778 14030
rect 13898 13990 13938 14030
rect 14058 13990 14098 14030
rect 14218 13990 14258 14030
rect 14378 13990 14418 14030
rect 14538 13990 14578 14030
rect 14698 13990 14738 14030
rect 14858 13990 14898 14030
rect 15018 13990 15058 14030
rect 15178 13990 15218 14030
rect 11918 13720 11958 13760
rect 14598 13720 14638 13760
rect 10758 13120 10798 13160
rect 10938 13080 10978 13120
rect 11178 13080 11218 13120
rect 11418 13080 11458 13120
rect 11658 13080 11698 13120
rect 12298 13080 12338 13120
rect 12538 13080 12578 13120
rect 12778 13080 12818 13120
rect 13078 13110 13118 13150
rect 15758 13600 15798 13640
rect 15758 13500 15798 13540
rect 15758 13400 15798 13440
rect 23228 13450 23288 13510
rect 15758 13300 15798 13340
rect 15758 13200 15798 13240
rect 13438 13110 13478 13150
rect 13738 13080 13778 13120
rect 13978 13080 14018 13120
rect 14218 13080 14258 13120
rect 14858 13080 14898 13120
rect 15098 13080 15138 13120
rect 15338 13080 15378 13120
rect 15578 13080 15618 13120
rect 23028 13130 23031 13170
rect 23031 13130 23065 13170
rect 23065 13130 23068 13170
rect 11441 12708 11475 12742
rect 11801 12708 11835 12742
rect 11921 12708 11955 12742
rect 12281 12708 12315 12742
rect 12401 12708 12435 12742
rect 12818 12680 12858 12720
rect 11378 12590 11418 12630
rect 11498 12590 11538 12630
rect 11618 12590 11658 12630
rect 11738 12590 11778 12630
rect 11858 12590 11898 12630
rect 11978 12590 12018 12630
rect 12098 12590 12138 12630
rect 12218 12590 12258 12630
rect 12338 12590 12378 12630
rect 12458 12590 12498 12630
rect 12578 12590 12618 12630
rect 12818 12600 12858 12640
rect 11542 12478 11576 12512
rect 11700 12478 11734 12512
rect 12024 12478 12058 12512
rect 12178 12478 12212 12512
rect 12502 12478 12536 12512
rect 12818 12520 12858 12560
rect 13698 12680 13738 12720
rect 14121 12708 14155 12742
rect 14241 12708 14275 12742
rect 14601 12708 14635 12742
rect 14721 12708 14755 12742
rect 15081 12708 15115 12742
rect 20338 12740 20378 12780
rect 20738 12740 20778 12780
rect 13698 12600 13738 12640
rect 13938 12590 13978 12630
rect 14058 12590 14098 12630
rect 14178 12590 14218 12630
rect 14298 12590 14338 12630
rect 14418 12590 14458 12630
rect 14538 12590 14578 12630
rect 14658 12590 14698 12630
rect 14778 12590 14818 12630
rect 14898 12590 14938 12630
rect 15018 12590 15058 12630
rect 15138 12590 15178 12630
rect 19538 12620 19578 12660
rect 13698 12520 13738 12560
rect 14020 12478 14054 12512
rect 14344 12478 14378 12512
rect 14498 12478 14532 12512
rect 14822 12478 14856 12512
rect 14980 12478 15014 12512
rect 19538 12520 19578 12560
rect 19538 12420 19578 12460
rect 19538 12320 19578 12360
rect 19538 12220 19578 12260
rect 19738 12620 19778 12660
rect 19738 12520 19778 12560
rect 19738 12420 19778 12460
rect 19738 12320 19778 12360
rect 19738 12220 19778 12260
rect 19938 12620 19978 12660
rect 19938 12520 19978 12560
rect 19938 12420 19978 12460
rect 19938 12320 19978 12360
rect 19938 12220 19978 12260
rect 20138 12620 20178 12660
rect 20138 12520 20178 12560
rect 20138 12420 20178 12460
rect 20138 12320 20178 12360
rect 20138 12220 20178 12260
rect 20338 12620 20378 12660
rect 20338 12520 20378 12560
rect 20338 12420 20378 12460
rect 20338 12320 20378 12360
rect 20338 12220 20378 12260
rect 20538 12620 20578 12660
rect 20538 12520 20578 12560
rect 20538 12420 20578 12460
rect 20538 12320 20578 12360
rect 20538 12220 20578 12260
rect 20738 12620 20778 12660
rect 20738 12520 20778 12560
rect 20738 12420 20778 12460
rect 20738 12320 20778 12360
rect 20738 12220 20778 12260
rect 20938 12620 20978 12660
rect 20938 12520 20978 12560
rect 20938 12420 20978 12460
rect 20938 12320 20978 12360
rect 20938 12220 20978 12260
rect 21138 12620 21178 12660
rect 21138 12520 21178 12560
rect 21138 12420 21178 12460
rect 21138 12320 21178 12360
rect 21138 12220 21178 12260
rect 21338 12620 21378 12660
rect 21338 12520 21378 12560
rect 21338 12420 21378 12460
rect 21338 12320 21378 12360
rect 21338 12220 21378 12260
rect 21538 12620 21578 12660
rect 21538 12520 21578 12560
rect 21538 12420 21578 12460
rect 21538 12320 21578 12360
rect 21538 12220 21578 12260
rect 19538 12100 19578 12140
rect 21538 12100 21578 12140
rect 23238 12733 23276 13130
rect 23238 12106 23276 12503
rect 21018 11940 21058 11980
rect 10718 11880 10758 11920
rect 10898 11870 10938 11910
rect 11378 11870 11418 11910
rect 11618 11870 11658 11910
rect 12098 11870 12138 11910
rect 12338 11870 12378 11910
rect 12758 11870 12798 11910
rect 13758 11870 13798 11910
rect 14178 11870 14218 11910
rect 14418 11870 14458 11910
rect 14898 11870 14938 11910
rect 15138 11870 15178 11910
rect 15618 11870 15658 11910
rect 15798 11880 15838 11920
rect 22138 11940 22178 11980
rect 10538 11750 10578 11790
rect 10538 11650 10578 11690
rect 10658 11750 10698 11790
rect 10658 11650 10698 11690
rect 10778 11750 10818 11790
rect 10778 11650 10818 11690
rect 10898 11750 10938 11790
rect 10898 11650 10938 11690
rect 11018 11750 11058 11790
rect 11018 11650 11058 11690
rect 11138 11750 11178 11790
rect 11138 11650 11178 11690
rect 11258 11750 11298 11790
rect 11258 11650 11298 11690
rect 11378 11750 11418 11790
rect 11378 11650 11418 11690
rect 11498 11750 11538 11790
rect 11498 11650 11538 11690
rect 11618 11750 11658 11790
rect 11618 11650 11658 11690
rect 11738 11750 11778 11790
rect 11738 11650 11778 11690
rect 11858 11750 11898 11790
rect 11858 11650 11898 11690
rect 11978 11750 12018 11790
rect 11978 11650 12018 11690
rect 12098 11750 12138 11790
rect 12098 11650 12138 11690
rect 12218 11750 12258 11790
rect 12218 11650 12258 11690
rect 12338 11750 12378 11790
rect 12338 11650 12378 11690
rect 12458 11750 12498 11790
rect 12458 11650 12498 11690
rect 12578 11750 12618 11790
rect 12578 11650 12618 11690
rect 12698 11750 12738 11790
rect 12698 11650 12738 11690
rect 12818 11750 12858 11790
rect 12818 11650 12858 11690
rect 12938 11750 12978 11790
rect 12938 11650 12978 11690
rect 13578 11750 13618 11790
rect 13578 11650 13618 11690
rect 13698 11750 13738 11790
rect 13698 11650 13738 11690
rect 13818 11750 13858 11790
rect 13818 11650 13858 11690
rect 13938 11750 13978 11790
rect 13938 11650 13978 11690
rect 14058 11750 14098 11790
rect 14058 11650 14098 11690
rect 14178 11750 14218 11790
rect 14178 11650 14218 11690
rect 14298 11750 14338 11790
rect 14298 11650 14338 11690
rect 14418 11750 14458 11790
rect 14418 11650 14458 11690
rect 14538 11750 14578 11790
rect 14538 11650 14578 11690
rect 14658 11750 14698 11790
rect 14658 11650 14698 11690
rect 14778 11750 14818 11790
rect 14778 11650 14818 11690
rect 14898 11750 14938 11790
rect 14898 11650 14938 11690
rect 15018 11750 15058 11790
rect 15018 11650 15058 11690
rect 15138 11750 15178 11790
rect 15138 11650 15178 11690
rect 15258 11750 15298 11790
rect 15258 11650 15298 11690
rect 15378 11750 15418 11790
rect 15378 11650 15418 11690
rect 15498 11750 15538 11790
rect 15498 11650 15538 11690
rect 15618 11750 15658 11790
rect 15618 11650 15658 11690
rect 15738 11750 15778 11790
rect 15738 11650 15778 11690
rect 15858 11750 15898 11790
rect 15858 11650 15898 11690
rect 15978 11750 16018 11790
rect 19938 11830 19978 11870
rect 15978 11650 16018 11690
rect 19468 11670 19508 11710
rect 10538 11530 10578 11570
rect 12938 11530 12978 11570
rect 13578 11530 13618 11570
rect 15978 11530 16018 11570
rect 19468 11570 19508 11610
rect 19598 11670 19638 11710
rect 19598 11570 19638 11610
rect 19728 11670 19768 11710
rect 19728 11570 19768 11610
rect 19858 11670 19898 11710
rect 19858 11570 19898 11610
rect 19988 11670 20028 11710
rect 19988 11570 20028 11610
rect 20118 11670 20158 11710
rect 20118 11570 20158 11610
rect 20248 11670 20288 11710
rect 20248 11570 20288 11610
rect 20608 11670 20648 11710
rect 20608 11570 20648 11610
rect 20738 11670 20778 11710
rect 20738 11570 20778 11610
rect 20868 11670 20908 11710
rect 20868 11570 20908 11610
rect 20998 11670 21038 11710
rect 20998 11570 21038 11610
rect 21128 11670 21168 11710
rect 21128 11570 21168 11610
rect 21258 11670 21298 11710
rect 21258 11570 21298 11610
rect 21388 11670 21428 11710
rect 21388 11570 21428 11610
rect 19638 11450 19678 11490
rect 20078 11450 20118 11490
rect 20868 11440 20908 11480
rect 21918 11450 21958 11490
rect 23458 11510 23528 11580
rect 22758 11450 22798 11490
rect 21918 11230 21958 11270
rect 23628 11280 23668 11320
rect 19728 11110 19768 11150
rect 20778 11110 20818 11150
rect 21218 11110 21258 11150
rect 22758 11110 22798 11150
rect 19468 10990 19508 11030
rect 19598 10990 19638 11030
rect 19728 10990 19768 11030
rect 19858 10990 19898 11030
rect 19988 10990 20028 11030
rect 20118 10990 20158 11030
rect 20248 10990 20288 11030
rect 20608 10990 20648 11030
rect 20738 10990 20778 11030
rect 20868 10990 20908 11030
rect 20998 10990 21038 11030
rect 21128 10990 21168 11030
rect 21258 10990 21298 11030
rect 21388 10990 21428 11030
rect 23458 11000 23528 11070
rect 20998 10830 21038 10870
rect 11908 10710 11948 10750
rect 12088 10710 12128 10750
rect 12268 10710 12308 10750
rect 12448 10710 12488 10750
rect 12628 10710 12668 10750
rect 12808 10710 12848 10750
rect 12988 10710 13028 10750
rect 13168 10710 13208 10750
rect 13348 10710 13388 10750
rect 13528 10710 13568 10750
rect 13708 10710 13748 10750
rect 13888 10710 13928 10750
rect 14068 10710 14108 10750
rect 14248 10710 14288 10750
rect 14428 10710 14468 10750
rect 14608 10710 14648 10750
rect 19858 10720 19898 10760
rect 22138 10720 22178 10760
rect 11638 10590 11678 10630
rect 11638 10490 11678 10530
rect 11638 10390 11678 10430
rect 11638 10290 11678 10330
rect 11638 10190 11678 10230
rect 11638 10090 11678 10130
rect 11818 10590 11858 10630
rect 11818 10490 11858 10530
rect 11818 10390 11858 10430
rect 11818 10290 11858 10330
rect 11818 10190 11858 10230
rect 11818 10090 11858 10130
rect 11998 10590 12038 10630
rect 11998 10490 12038 10530
rect 11998 10390 12038 10430
rect 11998 10290 12038 10330
rect 11998 10190 12038 10230
rect 11998 10090 12038 10130
rect 12178 10590 12218 10630
rect 12178 10490 12218 10530
rect 12178 10390 12218 10430
rect 12178 10290 12218 10330
rect 12178 10190 12218 10230
rect 12178 10090 12218 10130
rect 12358 10590 12398 10630
rect 12358 10490 12398 10530
rect 12358 10390 12398 10430
rect 12358 10290 12398 10330
rect 12358 10190 12398 10230
rect 12358 10090 12398 10130
rect 12538 10590 12578 10630
rect 12538 10490 12578 10530
rect 12538 10390 12578 10430
rect 12538 10290 12578 10330
rect 12538 10190 12578 10230
rect 12538 10090 12578 10130
rect 12718 10590 12758 10630
rect 12718 10490 12758 10530
rect 12718 10390 12758 10430
rect 12718 10290 12758 10330
rect 12718 10190 12758 10230
rect 12718 10090 12758 10130
rect 12898 10590 12938 10630
rect 12898 10490 12938 10530
rect 12898 10390 12938 10430
rect 12898 10290 12938 10330
rect 12898 10190 12938 10230
rect 12898 10090 12938 10130
rect 13078 10590 13118 10630
rect 13078 10490 13118 10530
rect 13078 10390 13118 10430
rect 13078 10290 13118 10330
rect 13078 10190 13118 10230
rect 13078 10090 13118 10130
rect 13258 10590 13298 10630
rect 13258 10490 13298 10530
rect 13258 10390 13298 10430
rect 13258 10290 13298 10330
rect 13258 10190 13298 10230
rect 13258 10090 13298 10130
rect 13438 10590 13478 10630
rect 13438 10490 13478 10530
rect 13438 10390 13478 10430
rect 13438 10290 13478 10330
rect 13438 10190 13478 10230
rect 13438 10090 13478 10130
rect 13618 10590 13658 10630
rect 13618 10490 13658 10530
rect 13618 10390 13658 10430
rect 13618 10290 13658 10330
rect 13618 10190 13658 10230
rect 13618 10090 13658 10130
rect 13798 10590 13838 10630
rect 13798 10490 13838 10530
rect 13798 10390 13838 10430
rect 13798 10290 13838 10330
rect 13798 10190 13838 10230
rect 13798 10090 13838 10130
rect 13978 10590 14018 10630
rect 13978 10490 14018 10530
rect 13978 10390 14018 10430
rect 13978 10290 14018 10330
rect 13978 10190 14018 10230
rect 13978 10090 14018 10130
rect 14158 10590 14198 10630
rect 14158 10490 14198 10530
rect 14158 10390 14198 10430
rect 14158 10290 14198 10330
rect 14158 10190 14198 10230
rect 14158 10090 14198 10130
rect 14338 10590 14378 10630
rect 14338 10490 14378 10530
rect 14338 10390 14378 10430
rect 14338 10290 14378 10330
rect 14338 10190 14378 10230
rect 14338 10090 14378 10130
rect 14518 10590 14558 10630
rect 14518 10490 14558 10530
rect 14518 10390 14558 10430
rect 14518 10290 14558 10330
rect 14518 10190 14558 10230
rect 14518 10090 14558 10130
rect 14698 10590 14738 10630
rect 14698 10490 14738 10530
rect 14698 10390 14738 10430
rect 14698 10290 14738 10330
rect 14698 10190 14738 10230
rect 14698 10090 14738 10130
rect 14878 10590 14918 10630
rect 19418 10570 19458 10610
rect 20998 10610 21038 10650
rect 14878 10490 14918 10530
rect 15608 10510 15648 10550
rect 15728 10510 15768 10550
rect 21418 10570 21458 10610
rect 15848 10510 15888 10550
rect 14878 10390 14918 10430
rect 14878 10290 14918 10330
rect 15508 10390 15548 10430
rect 15508 10290 15548 10330
rect 15618 10390 15658 10430
rect 15618 10290 15658 10330
rect 15728 10390 15768 10430
rect 15728 10290 15768 10330
rect 15838 10390 15878 10430
rect 15838 10290 15878 10330
rect 15948 10390 15988 10430
rect 15948 10290 15988 10330
rect 19618 10440 19658 10490
rect 19618 10300 19658 10350
rect 20018 10440 20058 10490
rect 20018 10300 20058 10350
rect 20418 10440 20458 10490
rect 20418 10300 20458 10350
rect 20818 10440 20858 10490
rect 20818 10300 20858 10350
rect 21218 10440 21258 10490
rect 21218 10300 21258 10350
rect 14878 10190 14918 10230
rect 15508 10170 15548 10210
rect 15728 10170 15768 10210
rect 15948 10170 15988 10210
rect 14878 10090 14918 10130
rect 11638 9970 11678 10010
rect 11998 9970 12038 10010
rect 12358 9970 12398 10010
rect 12718 9970 12758 10010
rect 13078 9970 13118 10010
rect 13438 9970 13478 10010
rect 13798 9970 13838 10010
rect 14158 9970 14198 10010
rect 14518 9970 14558 10010
rect 14878 9970 14918 10010
rect 19158 9990 19198 10030
rect 11816 9708 11850 9742
rect 11926 9708 11960 9742
rect 12036 9708 12070 9742
rect 12146 9708 12180 9742
rect 12256 9708 12290 9742
rect 12366 9708 12400 9742
rect 12476 9708 12510 9742
rect 12586 9708 12620 9742
rect 12696 9708 12730 9742
rect 12806 9708 12840 9742
rect 13716 9708 13750 9742
rect 13826 9708 13860 9742
rect 13936 9708 13970 9742
rect 14046 9708 14080 9742
rect 14156 9708 14190 9742
rect 14266 9708 14300 9742
rect 14376 9708 14410 9742
rect 14486 9708 14520 9742
rect 14596 9708 14630 9742
rect 14706 9708 14740 9742
rect 11568 9590 11608 9630
rect 11648 9590 11688 9630
rect 11568 9490 11608 9530
rect 11648 9490 11688 9530
rect 11758 9590 11798 9630
rect 11758 9490 11798 9530
rect 11868 9590 11908 9630
rect 11868 9490 11908 9530
rect 11978 9590 12018 9630
rect 11978 9490 12018 9530
rect 12088 9590 12128 9630
rect 12088 9490 12128 9530
rect 12198 9590 12238 9630
rect 12198 9490 12238 9530
rect 12308 9590 12348 9630
rect 12308 9490 12348 9530
rect 12418 9590 12458 9630
rect 12418 9490 12458 9530
rect 12528 9590 12568 9630
rect 12528 9490 12568 9530
rect 12638 9590 12678 9630
rect 12638 9490 12678 9530
rect 12748 9590 12788 9630
rect 12748 9490 12788 9530
rect 12858 9590 12898 9630
rect 12858 9490 12898 9530
rect 12968 9590 13008 9630
rect 13048 9590 13088 9630
rect 12968 9490 13008 9530
rect 13048 9490 13088 9530
rect 13468 9590 13508 9630
rect 13548 9590 13588 9630
rect 13468 9490 13508 9530
rect 13548 9490 13588 9530
rect 13658 9590 13698 9630
rect 13658 9490 13698 9530
rect 13768 9590 13808 9630
rect 13768 9490 13808 9530
rect 13878 9590 13918 9630
rect 13878 9490 13918 9530
rect 13988 9590 14028 9630
rect 13988 9490 14028 9530
rect 14098 9590 14138 9630
rect 14098 9490 14138 9530
rect 14208 9590 14248 9630
rect 14208 9490 14248 9530
rect 14318 9590 14358 9630
rect 14318 9490 14358 9530
rect 14428 9590 14468 9630
rect 14428 9490 14468 9530
rect 14538 9590 14578 9630
rect 14538 9490 14578 9530
rect 14648 9590 14688 9630
rect 14648 9490 14688 9530
rect 14758 9590 14798 9630
rect 14758 9490 14798 9530
rect 14868 9590 14908 9630
rect 14948 9590 14988 9630
rect 23238 10213 23276 10610
rect 23028 9600 23031 9640
rect 23031 9600 23065 9640
rect 23065 9600 23068 9640
rect 23238 9642 23276 10039
rect 14868 9490 14908 9530
rect 14948 9490 14988 9530
rect 11648 9370 11688 9410
rect 12968 9370 13008 9410
rect 13548 9370 13588 9410
rect 14868 9370 14908 9410
rect 23228 9070 23288 9130
rect 23108 8310 23178 8380
rect 13268 8250 13308 8290
rect 13488 8250 13528 8290
rect 13788 8250 13828 8290
rect 14018 8250 14058 8290
rect 14168 8250 14208 8290
rect 14388 8250 14428 8290
rect 14688 8250 14728 8290
rect 14908 8250 14948 8290
rect 15308 8250 15348 8290
rect 15638 8250 15678 8290
rect 15968 8250 16008 8290
rect 16408 8250 16448 8290
rect 17188 8250 17228 8290
rect 17868 8250 17908 8290
rect 16918 8140 16958 8180
rect 17548 8140 17588 8180
rect 19358 8090 19398 8130
rect 22398 8090 22438 8130
rect 19358 7970 19398 8010
rect 13148 7760 13188 7800
rect 15068 7750 15108 7790
rect 16098 7750 16138 7790
rect 16248 7760 16288 7800
rect 19358 7870 19398 7910
rect 18018 7800 18058 7840
rect 19358 7770 19398 7810
rect 19358 7670 19398 7710
rect 19578 7970 19618 8010
rect 19578 7870 19618 7910
rect 19578 7770 19618 7810
rect 19578 7670 19618 7710
rect 19798 7970 19838 8010
rect 19798 7870 19838 7910
rect 19798 7770 19838 7810
rect 19798 7670 19838 7710
rect 20018 7970 20058 8010
rect 20018 7870 20058 7910
rect 20018 7770 20058 7810
rect 20018 7670 20058 7710
rect 20238 7970 20278 8010
rect 20338 7970 20378 8010
rect 20438 7970 20478 8010
rect 20238 7870 20278 7910
rect 20338 7870 20378 7910
rect 20438 7870 20478 7910
rect 20238 7770 20278 7810
rect 20338 7770 20378 7810
rect 20438 7770 20478 7810
rect 20238 7670 20278 7710
rect 20338 7670 20378 7710
rect 20438 7670 20478 7710
rect 20658 7970 20698 8010
rect 20658 7870 20698 7910
rect 20658 7770 20698 7810
rect 20658 7670 20698 7710
rect 20878 7970 20918 8010
rect 20878 7870 20918 7910
rect 20878 7770 20918 7810
rect 20878 7670 20918 7710
rect 21098 7970 21138 8010
rect 21098 7870 21138 7910
rect 21098 7770 21138 7810
rect 21098 7670 21138 7710
rect 21318 7970 21358 8010
rect 21418 7970 21458 8010
rect 21518 7970 21558 8010
rect 21318 7870 21358 7910
rect 21418 7870 21458 7910
rect 21518 7870 21558 7910
rect 21318 7770 21358 7810
rect 21418 7770 21458 7810
rect 21518 7770 21558 7810
rect 21318 7670 21358 7710
rect 21418 7670 21458 7710
rect 21518 7670 21558 7710
rect 21738 7970 21778 8010
rect 21738 7870 21778 7910
rect 21738 7770 21778 7810
rect 21738 7670 21778 7710
rect 21958 7970 21998 8010
rect 21958 7870 21998 7910
rect 21958 7770 21998 7810
rect 21958 7670 21998 7710
rect 22178 7970 22218 8010
rect 22178 7870 22218 7910
rect 22178 7770 22218 7810
rect 22178 7670 22218 7710
rect 22398 7970 22438 8010
rect 22398 7870 22438 7910
rect 22398 7770 22438 7810
rect 22398 7670 22438 7710
rect 19798 7560 19838 7600
rect 21828 7520 21868 7560
rect 22088 7520 22128 7560
rect 22758 7520 22828 7590
rect 13718 7180 13758 7220
rect 16838 7180 16878 7220
rect 17478 7180 17518 7220
rect 13268 7070 13308 7110
rect 14008 7070 14048 7110
rect 14168 7070 14208 7110
rect 14908 7070 14948 7110
rect 15158 7070 15198 7110
rect 15348 7070 15388 7110
rect 15428 7070 15468 7110
rect 15638 7070 15678 7110
rect 15968 7070 16008 7110
rect 16408 7070 16448 7110
rect 16798 7070 16838 7110
rect 17188 7070 17228 7110
rect 17868 7070 17908 7110
rect 15268 6960 15308 7000
rect 20218 6990 20258 7030
rect 21388 7020 21428 7060
rect 22088 7020 22128 7060
rect 22758 6990 22828 7060
rect 13148 6380 13188 6420
rect 19558 6870 19598 6910
rect 19558 6770 19598 6810
rect 19558 6670 19598 6710
rect 19558 6570 19598 6610
rect 19778 6870 19818 6910
rect 19778 6770 19818 6810
rect 19778 6670 19818 6710
rect 19778 6570 19818 6610
rect 19998 6870 20038 6910
rect 19998 6770 20038 6810
rect 19998 6670 20038 6710
rect 19998 6570 20038 6610
rect 20218 6870 20258 6910
rect 20218 6770 20258 6810
rect 20218 6670 20258 6710
rect 20218 6570 20258 6610
rect 20438 6870 20478 6910
rect 20438 6770 20478 6810
rect 20438 6670 20478 6710
rect 20438 6570 20478 6610
rect 20658 6870 20698 6910
rect 20658 6770 20698 6810
rect 20658 6670 20698 6710
rect 20658 6570 20698 6610
rect 20878 6870 20918 6910
rect 20978 6870 21018 6910
rect 21078 6870 21118 6910
rect 20878 6770 20918 6810
rect 20978 6770 21018 6810
rect 21078 6770 21118 6810
rect 20878 6670 20918 6710
rect 20978 6670 21018 6710
rect 21078 6670 21118 6710
rect 20878 6570 20918 6610
rect 20978 6570 21018 6610
rect 21078 6570 21118 6610
rect 21298 6870 21338 6910
rect 21298 6770 21338 6810
rect 21298 6670 21338 6710
rect 21298 6570 21338 6610
rect 21518 6870 21558 6910
rect 21518 6770 21558 6810
rect 21518 6670 21558 6710
rect 21518 6570 21558 6610
rect 21738 6870 21778 6910
rect 21738 6770 21778 6810
rect 21738 6670 21778 6710
rect 21738 6570 21778 6610
rect 21958 6870 21998 6910
rect 21958 6770 21998 6810
rect 21958 6670 21998 6710
rect 21958 6570 21998 6610
rect 22178 6870 22218 6910
rect 22178 6770 22218 6810
rect 22178 6670 22218 6710
rect 22178 6570 22218 6610
rect 22398 6870 22438 6910
rect 22398 6770 22438 6810
rect 22398 6670 22438 6710
rect 22398 6570 22438 6610
rect 15048 6350 15088 6390
rect 16138 6390 16178 6430
rect 16268 6360 16308 6400
rect 17708 6420 17748 6460
rect 19558 6450 19598 6490
rect 22398 6450 22438 6490
rect 18018 6340 18058 6380
rect 13678 6000 13718 6040
rect 15398 6000 15438 6040
rect 17478 6000 17518 6040
rect 13268 5890 13308 5930
rect 13488 5890 13528 5930
rect 13788 5890 13828 5930
rect 14008 5890 14048 5930
rect 14168 5890 14208 5930
rect 14388 5890 14428 5930
rect 14688 5890 14728 5930
rect 14908 5890 14948 5930
rect 15208 5890 15248 5930
rect 15648 5890 15688 5930
rect 15978 5890 16018 5930
rect 16408 5890 16448 5930
rect 16798 5890 16838 5930
rect 17188 5890 17228 5930
rect 22998 5810 23068 5880
rect 23598 5490 23638 5530
rect 24118 5490 24158 5530
rect 24638 5490 24678 5530
rect 25158 5490 25198 5530
rect 23218 5360 23258 5400
rect 23218 5260 23258 5300
rect 23218 5160 23258 5200
rect 23218 5060 23258 5100
rect 23598 5360 23638 5400
rect 23598 5260 23638 5300
rect 23598 5160 23638 5200
rect 23598 5060 23638 5100
rect 23738 5360 23778 5400
rect 23738 5260 23778 5300
rect 23738 5160 23778 5200
rect 23738 5060 23778 5100
rect 24118 5360 24158 5400
rect 24118 5260 24158 5300
rect 24118 5160 24158 5200
rect 24118 5060 24158 5100
rect 24258 5360 24298 5400
rect 24258 5260 24298 5300
rect 24258 5160 24298 5200
rect 24258 5060 24298 5100
rect 24638 5360 24678 5400
rect 24638 5260 24678 5300
rect 24638 5160 24678 5200
rect 24638 5060 24678 5100
rect 24778 5360 24818 5400
rect 24778 5260 24818 5300
rect 24778 5160 24818 5200
rect 24778 5060 24818 5100
rect 25158 5360 25198 5400
rect 25158 5260 25198 5300
rect 25158 5160 25198 5200
rect 25158 5060 25198 5100
rect 23408 4940 23448 4980
rect 23928 4940 23968 4980
rect 24448 4940 24488 4980
rect 24968 4940 25008 4980
rect 12718 3690 12758 3730
rect 13138 3690 13178 3730
rect 13808 3690 13848 3730
rect 14378 3690 14418 3730
rect 15088 3690 15128 3730
rect 15518 3690 15558 3730
rect 15958 3690 15998 3730
rect 16208 3690 16248 3730
rect 16428 3690 16468 3730
rect 16898 3690 16938 3730
rect 17338 3690 17378 3730
rect 17958 3690 17998 3730
rect 18298 3690 18338 3730
rect 18658 3690 18698 3730
rect 19258 3690 19298 3730
rect 19598 3690 19638 3730
rect 19958 3690 19998 3730
rect 20558 3690 20598 3730
rect 20898 3690 20938 3730
rect 21258 3690 21298 3730
rect 21858 3690 21898 3730
rect 22198 3690 22238 3730
rect 22558 3690 22598 3730
rect 13038 3580 13078 3620
rect 13228 3580 13268 3620
rect 13348 3560 13388 3600
rect 14158 3580 14198 3620
rect 14288 3580 14328 3620
rect 15418 3580 15458 3620
rect 15638 3580 15678 3620
rect 16768 3590 16808 3630
rect 17178 3590 17218 3630
rect 19128 3580 19168 3620
rect 19708 3580 19748 3620
rect 20428 3580 20468 3620
rect 21008 3580 21048 3620
rect 21728 3580 21768 3620
rect 22308 3580 22348 3620
rect 12338 3290 12378 3330
rect 14748 3460 14788 3500
rect 14008 3260 14048 3300
rect 14528 3260 14568 3300
rect 16248 3270 16288 3310
rect 12398 3020 12438 3060
rect 13348 3040 13388 3080
rect 13478 3030 13518 3070
rect 14418 3030 14458 3070
rect 15978 3030 16018 3070
rect 18582 3020 18622 3060
rect 23218 4670 23258 4710
rect 23218 4570 23258 4610
rect 23218 4470 23258 4510
rect 23218 4370 23258 4410
rect 23218 4270 23258 4310
rect 23218 4170 23258 4210
rect 23328 4670 23368 4710
rect 23328 4570 23368 4610
rect 23328 4470 23368 4510
rect 23328 4370 23368 4410
rect 23328 4270 23368 4310
rect 23328 4170 23368 4210
rect 23738 4670 23778 4710
rect 23738 4570 23778 4610
rect 23738 4470 23778 4510
rect 23738 4370 23778 4410
rect 23738 4270 23778 4310
rect 23738 4170 23778 4210
rect 23848 4670 23888 4710
rect 23848 4570 23888 4610
rect 23848 4470 23888 4510
rect 23848 4370 23888 4410
rect 23848 4270 23888 4310
rect 23848 4170 23888 4210
rect 24258 4670 24298 4710
rect 24258 4570 24298 4610
rect 24258 4470 24298 4510
rect 24258 4370 24298 4410
rect 24258 4270 24298 4310
rect 24258 4170 24298 4210
rect 24368 4670 24408 4710
rect 24368 4570 24408 4610
rect 24368 4470 24408 4510
rect 24368 4370 24408 4410
rect 24368 4270 24408 4310
rect 24368 4170 24408 4210
rect 23290 4058 23324 4092
rect 23810 4058 23844 4092
rect 24330 4058 24364 4092
rect 23216 3890 23256 3930
rect 23216 3790 23256 3830
rect 23216 3690 23256 3730
rect 23216 3590 23256 3630
rect 23328 3890 23368 3930
rect 23328 3790 23368 3830
rect 23328 3690 23368 3730
rect 23328 3590 23368 3630
rect 23736 3890 23776 3930
rect 23736 3790 23776 3830
rect 23736 3690 23776 3730
rect 23736 3590 23776 3630
rect 23848 3890 23888 3930
rect 23848 3790 23888 3830
rect 23848 3690 23888 3730
rect 23848 3590 23888 3630
rect 24256 3890 24296 3930
rect 24256 3790 24296 3830
rect 24256 3690 24296 3730
rect 24256 3590 24296 3630
rect 24368 3890 24408 3930
rect 24368 3790 24408 3830
rect 24368 3690 24408 3730
rect 24368 3590 24408 3630
rect 23262 3478 23296 3512
rect 23782 3478 23816 3512
rect 24302 3478 24336 3512
rect 22762 3288 22796 3322
rect 12558 2910 12598 2950
rect 12778 2910 12818 2950
rect 13248 2910 13288 2950
rect 13588 2910 13628 2950
rect 13808 2910 13848 2950
rect 14248 2910 14288 2950
rect 14928 2910 14968 2950
rect 15148 2910 15188 2950
rect 15618 2910 15658 2950
rect 16078 2910 16118 2950
rect 16428 2910 16468 2950
rect 16678 2910 16718 2950
rect 16898 2910 16938 2950
rect 17228 2910 17268 2950
rect 17888 2910 17928 2950
rect 18108 2910 18148 2950
rect 18678 2910 18718 2950
rect 18938 2910 18978 2950
rect 19188 2910 19228 2950
rect 19408 2910 19448 2950
rect 19958 2910 19998 2950
rect 20238 2910 20278 2950
rect 20488 2910 20528 2950
rect 20708 2910 20748 2950
rect 21258 2910 21298 2950
rect 21538 2910 21578 2950
rect 21788 2910 21828 2950
rect 22008 2910 22048 2950
rect 22558 2910 22598 2950
rect 23262 3088 23296 3122
rect 23782 3088 23816 3122
rect 24302 3088 24336 3122
rect 23216 2970 23256 3010
rect 23216 2870 23256 2910
rect 23328 2970 23368 3010
rect 23328 2870 23368 2910
rect 23736 2970 23776 3010
rect 23736 2870 23776 2910
rect 23848 2970 23888 3010
rect 23848 2870 23888 2910
rect 24256 2970 24296 3010
rect 24256 2870 24296 2910
rect 24368 2970 24408 3010
rect 24368 2870 24408 2910
rect 23290 2708 23324 2742
rect 23810 2708 23844 2742
rect 24330 2708 24364 2742
rect 23218 2590 23258 2630
rect 23218 2490 23258 2530
rect 23218 2390 23258 2430
rect 23328 2590 23368 2630
rect 23328 2490 23368 2530
rect 23328 2390 23368 2430
rect 23738 2590 23778 2630
rect 23738 2490 23778 2530
rect 23738 2390 23778 2430
rect 23848 2590 23888 2630
rect 23848 2490 23888 2530
rect 23848 2390 23888 2430
rect 24258 2590 24298 2630
rect 24258 2490 24298 2530
rect 24258 2390 24298 2430
rect 24368 2590 24408 2630
rect 24368 2490 24408 2530
rect 24368 2390 24408 2430
rect 23276 2228 23310 2262
rect 23796 2228 23830 2262
rect 24316 2228 24350 2262
rect 24884 2228 24918 2262
rect 23218 2110 23258 2150
rect 23218 2010 23258 2050
rect 23328 2110 23368 2150
rect 23328 2010 23368 2050
rect 23738 2110 23778 2150
rect 23738 2010 23778 2050
rect 23848 2110 23888 2150
rect 23848 2010 23888 2050
rect 24258 2110 24298 2150
rect 24258 2010 24298 2050
rect 24368 2110 24408 2150
rect 24368 2010 24408 2050
rect 24858 2110 24898 2150
rect 24858 2010 24898 2050
rect 24968 2110 25008 2150
rect 24968 2010 25008 2050
rect 23328 1880 23368 1920
rect 23848 1880 23888 1920
rect 24368 1880 24408 1920
rect 24858 1880 24898 1920
<< metal1 >>
rect 16118 19690 16198 19700
rect 16118 19630 16128 19690
rect 16188 19630 16198 19690
rect 16118 19620 16198 19630
rect 25988 19510 26088 19520
rect 14988 19500 15418 19510
rect 14988 19440 14998 19500
rect 15408 19440 15418 19500
rect 14988 19430 15418 19440
rect 16898 19500 17328 19510
rect 16898 19440 16908 19500
rect 17318 19440 17328 19500
rect 16898 19430 17328 19440
rect 25988 19500 26478 19510
rect 25988 19440 26008 19500
rect 26068 19440 26098 19500
rect 26158 19440 26198 19500
rect 26258 19440 26308 19500
rect 26368 19440 26408 19500
rect 26468 19440 26478 19500
rect 25988 19420 26478 19440
rect 8868 19190 8948 19200
rect 8868 19130 8878 19190
rect 8938 19130 8948 19190
rect 8448 19080 8528 19090
rect 8448 19020 8458 19080
rect 8518 19020 8528 19080
rect 8448 19000 8528 19020
rect 8448 18940 8458 19000
rect 8518 18940 8528 19000
rect 8448 18920 8528 18940
rect 8448 18860 8458 18920
rect 8518 18860 8528 18920
rect 8448 18610 8528 18860
rect 8448 18570 8468 18610
rect 8508 18570 8528 18610
rect 8448 18550 8528 18570
rect 8448 18440 8528 18460
rect 8448 18040 8458 18440
rect 8518 18040 8528 18440
rect 8448 18030 8528 18040
rect 8868 18450 8948 19130
rect 8868 18390 8878 18450
rect 8938 18390 8948 18450
rect 8868 18370 8948 18390
rect 8868 18310 8878 18370
rect 8938 18310 8948 18370
rect 8868 18280 8948 18310
rect 8868 18220 8878 18280
rect 8938 18220 8948 18280
rect 8868 18190 8948 18220
rect 8868 18130 8878 18190
rect 8938 18130 8948 18190
rect 8868 18110 8948 18130
rect 8868 18050 8878 18110
rect 8938 18050 8948 18110
rect 8868 18030 8948 18050
rect 9238 19080 9318 19090
rect 9238 19020 9248 19080
rect 9308 19020 9318 19080
rect 9238 19000 9318 19020
rect 9238 18940 9248 19000
rect 9308 18940 9318 19000
rect 9238 18920 9318 18940
rect 9238 18860 9248 18920
rect 9308 18860 9318 18920
rect 9238 18610 9318 18860
rect 9238 18570 9258 18610
rect 9298 18570 9318 18610
rect 9238 18450 9318 18570
rect 9238 18060 9248 18450
rect 9288 18060 9318 18450
rect 9238 18030 9318 18060
rect 10678 19080 10758 19090
rect 10678 19020 10688 19080
rect 10748 19020 10758 19080
rect 10678 19000 10758 19020
rect 10678 18940 10688 19000
rect 10748 18940 10758 19000
rect 10678 18920 10758 18940
rect 10678 18860 10688 18920
rect 10748 18860 10758 18920
rect 10678 18610 10758 18860
rect 10678 18570 10698 18610
rect 10738 18570 10758 18610
rect 10678 18440 10758 18570
rect 10678 18050 10698 18440
rect 10738 18050 10758 18440
rect 10678 18030 10758 18050
rect 8462 17631 8512 17643
rect 8462 17234 8468 17631
rect 8506 17234 8512 17631
rect 8462 17230 8512 17234
rect 8448 11580 8528 17230
rect 9568 17226 9648 17246
rect 9568 16836 9588 17226
rect 9628 16836 9648 17226
rect 8448 11520 8458 11580
rect 8518 11520 8528 11580
rect 8448 9760 8528 11520
rect 9458 14210 9538 14220
rect 9458 14150 9468 14210
rect 9528 14150 9538 14210
rect 9458 11090 9538 14150
rect 9568 12520 9648 16836
rect 10348 16700 10428 16720
rect 10348 16310 10368 16700
rect 10408 16310 10428 16700
rect 10348 14720 10428 16310
rect 10348 14660 10358 14720
rect 10418 14660 10428 14720
rect 10348 14650 10428 14660
rect 9568 12460 9578 12520
rect 9638 12460 9648 12520
rect 9568 11200 9648 12460
rect 9568 11140 9578 11200
rect 9638 11140 9648 11200
rect 9568 11130 9648 11140
rect 9678 14490 9758 14500
rect 9678 14430 9688 14490
rect 9748 14430 9758 14490
rect 9678 12750 9758 14430
rect 9678 12690 9688 12750
rect 9748 12690 9758 12750
rect 9458 11030 9468 11090
rect 9528 11030 9538 11090
rect 9458 11020 9538 11030
rect 8448 9700 8458 9760
rect 8518 9700 8528 9760
rect 8448 9690 8528 9700
rect 9678 9310 9758 12690
rect 10618 14380 10698 14390
rect 10618 14320 10628 14380
rect 10688 14320 10698 14380
rect 10618 12050 10698 14320
rect 11028 14380 11108 19200
rect 18188 19190 18268 19200
rect 18188 19130 18198 19190
rect 18258 19130 18268 19190
rect 13238 19080 13318 19090
rect 13238 19020 13248 19080
rect 13308 19020 13318 19080
rect 13238 19000 13318 19020
rect 13238 18940 13248 19000
rect 13308 18940 13318 19000
rect 13238 18920 13318 18940
rect 13238 18860 13248 18920
rect 13308 18860 13318 18920
rect 13238 18850 13318 18860
rect 15668 19080 15748 19090
rect 15668 19020 15678 19080
rect 15738 19020 15748 19080
rect 15668 19000 15748 19020
rect 15668 18940 15678 19000
rect 15738 18940 15748 19000
rect 15668 18920 15748 18940
rect 15668 18860 15678 18920
rect 15738 18860 15748 18920
rect 15668 18610 15748 18860
rect 15668 18570 15688 18610
rect 15728 18570 15748 18610
rect 11568 18414 14988 18490
rect 11568 18380 11658 18414
rect 11692 18380 11758 18414
rect 11792 18380 11858 18414
rect 11892 18380 11958 18414
rect 11992 18380 12058 18414
rect 12092 18380 12158 18414
rect 12192 18380 13018 18414
rect 13052 18380 13118 18414
rect 13152 18380 13218 18414
rect 13252 18380 13318 18414
rect 13352 18380 13418 18414
rect 13452 18380 13518 18414
rect 13552 18380 14378 18414
rect 14412 18380 14478 18414
rect 14512 18380 14578 18414
rect 14612 18380 14678 18414
rect 14712 18380 14778 18414
rect 14812 18380 14878 18414
rect 14912 18380 14988 18414
rect 11568 18314 14988 18380
rect 11568 18280 11658 18314
rect 11692 18280 11758 18314
rect 11792 18280 11858 18314
rect 11892 18280 11958 18314
rect 11992 18280 12058 18314
rect 12092 18280 12158 18314
rect 12192 18280 13018 18314
rect 13052 18280 13118 18314
rect 13152 18280 13218 18314
rect 13252 18280 13318 18314
rect 13352 18280 13418 18314
rect 13452 18280 13518 18314
rect 13552 18280 14378 18314
rect 14412 18280 14478 18314
rect 14512 18280 14578 18314
rect 14612 18280 14678 18314
rect 14712 18280 14778 18314
rect 14812 18280 14878 18314
rect 14912 18280 14988 18314
rect 11568 18214 14988 18280
rect 11568 18180 11658 18214
rect 11692 18180 11758 18214
rect 11792 18180 11858 18214
rect 11892 18180 11958 18214
rect 11992 18180 12058 18214
rect 12092 18180 12158 18214
rect 12192 18180 13018 18214
rect 13052 18180 13118 18214
rect 13152 18180 13218 18214
rect 13252 18180 13318 18214
rect 13352 18180 13418 18214
rect 13452 18180 13518 18214
rect 13552 18180 14378 18214
rect 14412 18180 14478 18214
rect 14512 18180 14578 18214
rect 14612 18180 14678 18214
rect 14712 18180 14778 18214
rect 14812 18180 14878 18214
rect 14912 18180 14988 18214
rect 11568 18114 14988 18180
rect 11568 18080 11658 18114
rect 11692 18080 11758 18114
rect 11792 18080 11858 18114
rect 11892 18080 11958 18114
rect 11992 18080 12058 18114
rect 12092 18080 12158 18114
rect 12192 18080 13018 18114
rect 13052 18080 13118 18114
rect 13152 18080 13218 18114
rect 13252 18080 13318 18114
rect 13352 18080 13418 18114
rect 13452 18080 13518 18114
rect 13552 18080 14378 18114
rect 14412 18080 14478 18114
rect 14512 18080 14578 18114
rect 14612 18080 14678 18114
rect 14712 18080 14778 18114
rect 14812 18080 14878 18114
rect 14912 18080 14988 18114
rect 11568 18014 14988 18080
rect 15668 18440 15748 18570
rect 15668 18050 15688 18440
rect 15728 18050 15748 18440
rect 15668 18030 15748 18050
rect 16778 19080 16858 19090
rect 16778 19020 16788 19080
rect 16848 19020 16858 19080
rect 16778 19000 16858 19020
rect 16778 18940 16788 19000
rect 16848 18940 16858 19000
rect 16778 18920 16858 18940
rect 16778 18860 16788 18920
rect 16848 18860 16858 18920
rect 16778 18610 16858 18860
rect 16778 18570 16798 18610
rect 16838 18570 16858 18610
rect 16778 18437 16858 18570
rect 17568 19080 17648 19090
rect 17568 19020 17578 19080
rect 17638 19020 17648 19080
rect 17568 19000 17648 19020
rect 17568 18940 17578 19000
rect 17638 18940 17648 19000
rect 17568 18920 17648 18940
rect 17568 18860 17578 18920
rect 17638 18860 17648 18920
rect 17568 18610 17648 18860
rect 18188 18850 18268 19130
rect 18188 18790 18198 18850
rect 18258 18790 18268 18850
rect 18188 18780 18268 18790
rect 17568 18570 17588 18610
rect 17628 18570 17648 18610
rect 17568 18550 17648 18570
rect 16778 18040 16801 18437
rect 16839 18040 16858 18437
rect 16778 18030 16858 18040
rect 17568 18440 17648 18460
rect 17568 18040 17578 18440
rect 17638 18040 17648 18440
rect 17568 18030 17648 18040
rect 17948 18450 18028 18460
rect 17948 18390 17958 18450
rect 18018 18390 18028 18450
rect 17948 18370 18028 18390
rect 17948 18310 17958 18370
rect 18018 18310 18028 18370
rect 17948 18280 18028 18310
rect 17948 18220 17958 18280
rect 18018 18220 18028 18280
rect 17948 18190 18028 18220
rect 17948 18130 17958 18190
rect 18018 18130 18028 18190
rect 17948 18110 18028 18130
rect 17948 18050 17958 18110
rect 18018 18050 18028 18110
rect 18638 18150 18738 18170
rect 18638 18090 18658 18150
rect 18718 18090 18738 18150
rect 18638 18070 18738 18090
rect 16795 18028 16845 18030
rect 11568 17980 11658 18014
rect 11692 17980 11758 18014
rect 11792 17980 11858 18014
rect 11892 17980 11958 18014
rect 11992 17980 12058 18014
rect 12092 17980 12158 18014
rect 12192 17980 13018 18014
rect 13052 17980 13118 18014
rect 13152 17980 13218 18014
rect 13252 17980 13318 18014
rect 13352 17980 13418 18014
rect 13452 17980 13518 18014
rect 13552 17980 14378 18014
rect 14412 17980 14478 18014
rect 14512 17980 14578 18014
rect 14612 17980 14678 18014
rect 14712 17980 14778 18014
rect 14812 17980 14878 18014
rect 14912 17980 14988 18014
rect 11568 17914 14988 17980
rect 11568 17880 11658 17914
rect 11692 17880 11758 17914
rect 11792 17880 11858 17914
rect 11892 17880 11958 17914
rect 11992 17880 12058 17914
rect 12092 17880 12158 17914
rect 12192 17880 13018 17914
rect 13052 17880 13118 17914
rect 13152 17880 13218 17914
rect 13252 17880 13318 17914
rect 13352 17880 13418 17914
rect 13452 17880 13518 17914
rect 13552 17880 14378 17914
rect 14412 17880 14478 17914
rect 14512 17880 14578 17914
rect 14612 17880 14678 17914
rect 14712 17880 14778 17914
rect 14812 17880 14878 17914
rect 14912 17880 14988 17914
rect 11568 17790 14988 17880
rect 11568 17054 12268 17790
rect 11568 17020 11658 17054
rect 11692 17020 11758 17054
rect 11792 17020 11858 17054
rect 11892 17020 11958 17054
rect 11992 17020 12058 17054
rect 12092 17020 12158 17054
rect 12192 17020 12268 17054
rect 11568 16954 12268 17020
rect 11568 16920 11658 16954
rect 11692 16920 11758 16954
rect 11792 16920 11858 16954
rect 11892 16920 11958 16954
rect 11992 16920 12058 16954
rect 12092 16920 12158 16954
rect 12192 16920 12268 16954
rect 11568 16854 12268 16920
rect 11568 16820 11658 16854
rect 11692 16820 11758 16854
rect 11792 16820 11858 16854
rect 11892 16820 11958 16854
rect 11992 16820 12058 16854
rect 12092 16820 12158 16854
rect 12192 16820 12268 16854
rect 11138 16810 11218 16820
rect 11138 16750 11148 16810
rect 11208 16750 11218 16810
rect 11138 14610 11218 16750
rect 11568 16810 12268 16820
rect 11568 16750 11578 16810
rect 11638 16754 12268 16810
rect 11638 16750 11658 16754
rect 11568 16720 11658 16750
rect 11692 16720 11758 16754
rect 11792 16720 11858 16754
rect 11892 16720 11958 16754
rect 11992 16720 12058 16754
rect 12092 16720 12158 16754
rect 12192 16720 12268 16754
rect 11568 16654 12268 16720
rect 11568 16620 11658 16654
rect 11692 16620 11758 16654
rect 11792 16620 11858 16654
rect 11892 16620 11958 16654
rect 11992 16620 12058 16654
rect 12092 16620 12158 16654
rect 12192 16620 12268 16654
rect 11568 16554 12268 16620
rect 11568 16520 11658 16554
rect 11692 16520 11758 16554
rect 11792 16520 11858 16554
rect 11892 16520 11958 16554
rect 11992 16520 12058 16554
rect 12092 16520 12158 16554
rect 12192 16520 12268 16554
rect 11568 15770 12268 16520
rect 12928 17054 13628 17130
rect 12928 17020 13018 17054
rect 13052 17020 13118 17054
rect 13152 17020 13218 17054
rect 13252 17020 13318 17054
rect 13352 17020 13418 17054
rect 13452 17020 13518 17054
rect 13552 17020 13628 17054
rect 12928 16954 13628 17020
rect 12928 16920 13018 16954
rect 13052 16920 13118 16954
rect 13152 16920 13218 16954
rect 13252 16920 13318 16954
rect 13352 16920 13418 16954
rect 13452 16920 13518 16954
rect 13552 16920 13628 16954
rect 12928 16854 13628 16920
rect 12928 16820 13018 16854
rect 13052 16820 13118 16854
rect 13152 16820 13218 16854
rect 13252 16820 13318 16854
rect 13352 16820 13418 16854
rect 13452 16820 13518 16854
rect 13552 16820 13628 16854
rect 12928 16810 13628 16820
rect 12928 16754 13248 16810
rect 13308 16754 13628 16810
rect 12928 16720 13018 16754
rect 13052 16720 13118 16754
rect 13152 16720 13218 16754
rect 13308 16750 13318 16754
rect 13252 16720 13318 16750
rect 13352 16720 13418 16754
rect 13452 16720 13518 16754
rect 13552 16720 13628 16754
rect 12928 16654 13628 16720
rect 12928 16620 13018 16654
rect 13052 16620 13118 16654
rect 13152 16620 13218 16654
rect 13252 16620 13318 16654
rect 13352 16620 13418 16654
rect 13452 16620 13518 16654
rect 13552 16620 13628 16654
rect 12928 16554 13628 16620
rect 12928 16520 13018 16554
rect 13052 16520 13118 16554
rect 13152 16520 13218 16554
rect 13252 16520 13318 16554
rect 13352 16520 13418 16554
rect 13452 16520 13518 16554
rect 13552 16520 13628 16554
rect 12928 16430 13628 16520
rect 14288 17054 14988 17790
rect 14288 17020 14378 17054
rect 14412 17020 14478 17054
rect 14512 17020 14578 17054
rect 14612 17020 14678 17054
rect 14712 17020 14778 17054
rect 14812 17020 14878 17054
rect 14912 17020 14988 17054
rect 14288 16954 14988 17020
rect 14288 16920 14378 16954
rect 14412 16920 14478 16954
rect 14512 16920 14578 16954
rect 14612 16920 14678 16954
rect 14712 16920 14778 16954
rect 14812 16920 14878 16954
rect 14912 16920 14988 16954
rect 14288 16854 14988 16920
rect 14288 16820 14378 16854
rect 14412 16820 14478 16854
rect 14512 16820 14578 16854
rect 14612 16820 14678 16854
rect 14712 16820 14778 16854
rect 14812 16820 14878 16854
rect 14912 16820 14988 16854
rect 16778 17838 16858 17850
rect 16778 17441 16801 17838
rect 16839 17441 16858 17838
rect 14288 16754 14988 16820
rect 14288 16720 14378 16754
rect 14412 16720 14478 16754
rect 14512 16720 14578 16754
rect 14612 16720 14678 16754
rect 14712 16720 14778 16754
rect 14812 16720 14878 16754
rect 14912 16720 14988 16754
rect 14288 16654 14988 16720
rect 14288 16620 14378 16654
rect 14412 16620 14478 16654
rect 14512 16620 14578 16654
rect 14612 16620 14678 16654
rect 14712 16620 14778 16654
rect 14812 16620 14878 16654
rect 14912 16620 14988 16654
rect 14288 16554 14988 16620
rect 14288 16520 14378 16554
rect 14412 16520 14478 16554
rect 14512 16520 14578 16554
rect 14612 16520 14678 16554
rect 14712 16520 14778 16554
rect 14812 16520 14878 16554
rect 14912 16520 14988 16554
rect 14288 15770 14988 16520
rect 11568 15694 14988 15770
rect 11568 15660 11658 15694
rect 11692 15660 11758 15694
rect 11792 15660 11858 15694
rect 11892 15660 11958 15694
rect 11992 15660 12058 15694
rect 12092 15660 12158 15694
rect 12192 15660 13018 15694
rect 13052 15660 13118 15694
rect 13152 15660 13218 15694
rect 13252 15660 13318 15694
rect 13352 15660 13418 15694
rect 13452 15660 13518 15694
rect 13552 15660 14378 15694
rect 14412 15660 14478 15694
rect 14512 15660 14578 15694
rect 14612 15660 14678 15694
rect 14712 15660 14778 15694
rect 14812 15660 14878 15694
rect 14912 15660 14988 15694
rect 11568 15594 14988 15660
rect 11568 15560 11658 15594
rect 11692 15560 11758 15594
rect 11792 15560 11858 15594
rect 11892 15560 11958 15594
rect 11992 15560 12058 15594
rect 12092 15560 12158 15594
rect 12192 15560 13018 15594
rect 13052 15560 13118 15594
rect 13152 15560 13218 15594
rect 13252 15560 13318 15594
rect 13352 15560 13418 15594
rect 13452 15560 13518 15594
rect 13552 15560 14378 15594
rect 14412 15560 14478 15594
rect 14512 15560 14578 15594
rect 14612 15560 14678 15594
rect 14712 15560 14778 15594
rect 14812 15560 14878 15594
rect 14912 15560 14988 15594
rect 11568 15494 14988 15560
rect 11568 15460 11658 15494
rect 11692 15460 11758 15494
rect 11792 15460 11858 15494
rect 11892 15460 11958 15494
rect 11992 15460 12058 15494
rect 12092 15460 12158 15494
rect 12192 15460 13018 15494
rect 13052 15460 13118 15494
rect 13152 15460 13218 15494
rect 13252 15460 13318 15494
rect 13352 15460 13418 15494
rect 13452 15460 13518 15494
rect 13552 15460 14378 15494
rect 14412 15460 14478 15494
rect 14512 15460 14578 15494
rect 14612 15460 14678 15494
rect 14712 15460 14778 15494
rect 14812 15460 14878 15494
rect 14912 15460 14988 15494
rect 11568 15394 14988 15460
rect 11568 15360 11658 15394
rect 11692 15360 11758 15394
rect 11792 15360 11858 15394
rect 11892 15360 11958 15394
rect 11992 15360 12058 15394
rect 12092 15360 12158 15394
rect 12192 15360 13018 15394
rect 13052 15360 13118 15394
rect 13152 15360 13218 15394
rect 13252 15360 13318 15394
rect 13352 15360 13418 15394
rect 13452 15360 13518 15394
rect 13552 15360 14378 15394
rect 14412 15360 14478 15394
rect 14512 15360 14578 15394
rect 14612 15360 14678 15394
rect 14712 15360 14778 15394
rect 14812 15360 14878 15394
rect 14912 15360 14988 15394
rect 11568 15294 14988 15360
rect 11568 15260 11658 15294
rect 11692 15260 11758 15294
rect 11792 15260 11858 15294
rect 11892 15260 11958 15294
rect 11992 15260 12058 15294
rect 12092 15260 12158 15294
rect 12192 15260 13018 15294
rect 13052 15260 13118 15294
rect 13152 15260 13218 15294
rect 13252 15260 13318 15294
rect 13352 15260 13418 15294
rect 13452 15260 13518 15294
rect 13552 15260 14378 15294
rect 14412 15260 14478 15294
rect 14512 15260 14578 15294
rect 14612 15260 14678 15294
rect 14712 15260 14778 15294
rect 14812 15260 14878 15294
rect 14912 15260 14988 15294
rect 11568 15194 14988 15260
rect 11568 15160 11658 15194
rect 11692 15160 11758 15194
rect 11792 15160 11858 15194
rect 11892 15160 11958 15194
rect 11992 15160 12058 15194
rect 12092 15160 12158 15194
rect 12192 15160 13018 15194
rect 13052 15160 13118 15194
rect 13152 15160 13218 15194
rect 13252 15160 13318 15194
rect 13352 15160 13418 15194
rect 13452 15160 13518 15194
rect 13552 15160 14378 15194
rect 14412 15160 14478 15194
rect 14512 15160 14578 15194
rect 14612 15160 14678 15194
rect 14712 15160 14778 15194
rect 14812 15160 14878 15194
rect 14912 15160 14988 15194
rect 11568 15070 14988 15160
rect 15338 16810 15418 16820
rect 15338 16750 15348 16810
rect 15408 16750 15418 16810
rect 15338 14800 15418 16750
rect 15338 14740 15348 14800
rect 15408 14740 15418 14800
rect 15338 14730 15418 14740
rect 15998 16700 16078 16720
rect 15998 16310 16018 16700
rect 16058 16310 16078 16700
rect 15998 14800 16078 16310
rect 16348 15350 16588 15370
rect 16348 15290 16358 15350
rect 16418 15290 16438 15350
rect 16498 15290 16518 15350
rect 16578 15290 16588 15350
rect 15998 14740 16008 14800
rect 16068 14740 16078 14800
rect 15998 14730 16078 14740
rect 16238 14800 16318 14810
rect 16238 14740 16248 14800
rect 16308 14740 16318 14800
rect 16238 14730 16318 14740
rect 13948 14720 14028 14730
rect 13948 14660 13958 14720
rect 14018 14660 14028 14720
rect 13948 14610 14028 14660
rect 11138 14550 11148 14610
rect 11208 14550 11218 14610
rect 11138 14540 11218 14550
rect 12540 14540 12550 14610
rect 12620 14540 12630 14610
rect 13938 14540 13948 14610
rect 14018 14540 14028 14610
rect 16148 14600 16228 14610
rect 16148 14540 16158 14600
rect 16218 14540 16228 14600
rect 16148 14530 16228 14540
rect 11028 14320 11038 14380
rect 11098 14320 11108 14380
rect 11028 14310 11108 14320
rect 15468 14250 15548 14260
rect 11078 14210 11158 14220
rect 11078 14150 11088 14210
rect 11148 14150 11158 14210
rect 11078 14140 11158 14150
rect 15468 14190 15478 14250
rect 15538 14190 15548 14250
rect 15468 14170 15548 14190
rect 15468 14110 15478 14170
rect 15538 14110 15548 14170
rect 15468 14100 15548 14110
rect 11158 14040 11238 14050
rect 11158 13980 11168 14040
rect 11228 13980 11238 14040
rect 11158 13970 11238 13980
rect 11318 14040 11398 14050
rect 11318 13980 11328 14040
rect 11388 13980 11398 14040
rect 11318 13970 11398 13980
rect 11478 14040 11558 14050
rect 11478 13980 11488 14040
rect 11548 13980 11558 14040
rect 11478 13970 11558 13980
rect 11638 14040 11718 14050
rect 11638 13980 11648 14040
rect 11708 13980 11718 14040
rect 11638 13970 11718 13980
rect 11798 14040 11878 14050
rect 11798 13980 11808 14040
rect 11868 13980 11878 14040
rect 11798 13970 11878 13980
rect 11958 14040 12038 14050
rect 11958 13980 11968 14040
rect 12028 13980 12038 14040
rect 11958 13970 12038 13980
rect 12118 14040 12198 14050
rect 12118 13980 12128 14040
rect 12188 13980 12198 14040
rect 12118 13970 12198 13980
rect 12278 14040 12358 14050
rect 12278 13980 12288 14040
rect 12348 13980 12358 14040
rect 12278 13970 12358 13980
rect 12438 14040 12518 14050
rect 12438 13980 12448 14040
rect 12508 13980 12518 14040
rect 12438 13970 12518 13980
rect 12598 14040 12678 14050
rect 12598 13980 12608 14040
rect 12668 13980 12678 14040
rect 12598 13970 12678 13980
rect 12758 14040 12838 14050
rect 12758 13980 12768 14040
rect 12828 13980 12838 14040
rect 12758 13970 12838 13980
rect 12918 14040 12998 14050
rect 12918 13980 12928 14040
rect 12988 13980 12998 14040
rect 12918 13970 12998 13980
rect 13078 14040 13158 14050
rect 13078 13980 13088 14040
rect 13148 13980 13158 14040
rect 13078 13970 13158 13980
rect 13238 14040 13318 14050
rect 13238 13980 13248 14040
rect 13308 13980 13318 14040
rect 13238 13970 13318 13980
rect 13398 14040 13478 14050
rect 13398 13980 13408 14040
rect 13468 13980 13478 14040
rect 13398 13970 13478 13980
rect 13558 14040 13638 14050
rect 13558 13980 13568 14040
rect 13628 13980 13638 14040
rect 13558 13970 13638 13980
rect 13718 14040 13798 14050
rect 13718 13980 13728 14040
rect 13788 13980 13798 14040
rect 13718 13970 13798 13980
rect 13878 14040 13958 14050
rect 13878 13980 13888 14040
rect 13948 13980 13958 14040
rect 13878 13970 13958 13980
rect 14038 14040 14118 14050
rect 14038 13980 14048 14040
rect 14108 13980 14118 14040
rect 14038 13970 14118 13980
rect 14198 14040 14278 14050
rect 14198 13980 14208 14040
rect 14268 13980 14278 14040
rect 14198 13970 14278 13980
rect 14358 14040 14438 14050
rect 14358 13980 14368 14040
rect 14428 13980 14438 14040
rect 14358 13970 14438 13980
rect 14518 14040 14598 14050
rect 14518 13980 14528 14040
rect 14588 13980 14598 14040
rect 14518 13970 14598 13980
rect 14678 14040 14758 14050
rect 14678 13980 14688 14040
rect 14748 13980 14758 14040
rect 14678 13970 14758 13980
rect 14838 14040 14918 14050
rect 14838 13980 14848 14040
rect 14908 13980 14918 14040
rect 14838 13970 14918 13980
rect 14998 14040 15078 14050
rect 14998 13980 15008 14040
rect 15068 13980 15078 14040
rect 14998 13970 15078 13980
rect 15158 14040 15238 14050
rect 15158 13980 15168 14040
rect 15228 13980 15238 14040
rect 15158 13970 15238 13980
rect 11898 13930 11978 13940
rect 11898 13870 11908 13930
rect 11968 13870 11978 13930
rect 11898 13850 11978 13870
rect 11898 13790 11908 13850
rect 11968 13790 11978 13850
rect 11898 13770 11978 13790
rect 11898 13710 11908 13770
rect 11968 13710 11978 13770
rect 11898 13700 11978 13710
rect 13158 13930 13398 13940
rect 13158 13870 13168 13930
rect 13228 13870 13248 13930
rect 13308 13870 13328 13930
rect 13388 13870 13398 13930
rect 13158 13850 13398 13870
rect 13158 13790 13168 13850
rect 13228 13790 13248 13850
rect 13308 13790 13328 13850
rect 13388 13790 13398 13850
rect 13158 13770 13398 13790
rect 13158 13710 13168 13770
rect 13228 13710 13248 13770
rect 13308 13710 13328 13770
rect 13388 13710 13398 13770
rect 10738 13160 10818 13180
rect 10738 13120 10758 13160
rect 10798 13120 10818 13160
rect 13068 13150 13128 13170
rect 10738 12860 10818 13120
rect 10918 13130 10998 13140
rect 10918 13070 10928 13130
rect 10988 13070 10998 13130
rect 10918 13050 10998 13070
rect 10918 12990 10928 13050
rect 10988 12990 10998 13050
rect 10918 12970 10998 12990
rect 10918 12910 10928 12970
rect 10988 12910 10998 12970
rect 10918 12900 10998 12910
rect 11158 13130 11238 13140
rect 11158 13070 11168 13130
rect 11228 13070 11238 13130
rect 11158 13050 11238 13070
rect 11158 12990 11168 13050
rect 11228 12990 11238 13050
rect 11158 12970 11238 12990
rect 11158 12910 11168 12970
rect 11228 12910 11238 12970
rect 11158 12900 11238 12910
rect 11398 13130 11478 13140
rect 11398 13070 11408 13130
rect 11468 13070 11478 13130
rect 11398 13050 11478 13070
rect 11398 12990 11408 13050
rect 11468 12990 11478 13050
rect 11398 12970 11478 12990
rect 11398 12910 11408 12970
rect 11468 12910 11478 12970
rect 11398 12900 11478 12910
rect 11638 13130 11718 13140
rect 11638 13070 11648 13130
rect 11708 13070 11718 13130
rect 11638 13050 11718 13070
rect 11638 12990 11648 13050
rect 11708 12990 11718 13050
rect 11638 12970 11718 12990
rect 11638 12910 11648 12970
rect 11708 12910 11718 12970
rect 11638 12900 11718 12910
rect 12278 13130 12358 13140
rect 12278 13070 12288 13130
rect 12348 13070 12358 13130
rect 12278 13050 12358 13070
rect 12278 12990 12288 13050
rect 12348 12990 12358 13050
rect 12278 12970 12358 12990
rect 12278 12910 12288 12970
rect 12348 12910 12358 12970
rect 12278 12900 12358 12910
rect 12518 13130 12598 13140
rect 12518 13070 12528 13130
rect 12588 13070 12598 13130
rect 12518 13050 12598 13070
rect 12518 12990 12528 13050
rect 12588 12990 12598 13050
rect 12518 12970 12598 12990
rect 12518 12910 12528 12970
rect 12588 12910 12598 12970
rect 12518 12900 12598 12910
rect 12758 13130 12838 13140
rect 12758 13070 12768 13130
rect 12828 13070 12838 13130
rect 12758 13050 12838 13070
rect 12758 12990 12768 13050
rect 12828 12990 12838 13050
rect 12758 12970 12838 12990
rect 12758 12910 12768 12970
rect 12828 12910 12838 12970
rect 12758 12900 12838 12910
rect 13068 13110 13078 13150
rect 13118 13110 13128 13150
rect 10738 12800 10748 12860
rect 10808 12800 10818 12860
rect 10738 12790 10818 12800
rect 11488 12860 11568 12870
rect 11488 12800 11498 12860
rect 11558 12800 11568 12860
rect 11488 12790 11568 12800
rect 11708 12860 11788 12870
rect 11708 12800 11718 12860
rect 11778 12800 11788 12860
rect 11708 12790 11788 12800
rect 11968 12860 12048 12870
rect 11968 12800 11978 12860
rect 12038 12800 12048 12860
rect 11968 12790 12048 12800
rect 12188 12860 12268 12870
rect 12188 12800 12198 12860
rect 12258 12800 12268 12860
rect 12188 12790 12268 12800
rect 12448 12860 12528 12870
rect 12448 12800 12458 12860
rect 12518 12800 12528 12860
rect 12448 12790 12528 12800
rect 11429 12750 11487 12760
rect 11429 12698 11431 12750
rect 11483 12698 11487 12750
rect 11429 12690 11487 12698
rect 11518 12650 11548 12790
rect 11728 12650 11758 12790
rect 11789 12750 11847 12760
rect 11789 12698 11791 12750
rect 11843 12698 11847 12750
rect 11789 12690 11847 12698
rect 11909 12750 11967 12760
rect 11909 12698 11911 12750
rect 11963 12698 11967 12750
rect 11909 12690 11967 12698
rect 11998 12650 12028 12790
rect 12208 12650 12238 12790
rect 12269 12750 12327 12760
rect 12269 12698 12271 12750
rect 12323 12698 12327 12750
rect 12269 12690 12327 12698
rect 12389 12750 12447 12760
rect 12389 12698 12391 12750
rect 12443 12698 12447 12750
rect 12389 12690 12447 12698
rect 12478 12650 12508 12790
rect 12798 12730 12878 12740
rect 12798 12670 12808 12730
rect 12868 12670 12878 12730
rect 12798 12650 12878 12670
rect 11368 12630 11428 12650
rect 11368 12590 11378 12630
rect 11418 12590 11428 12630
rect 11368 12320 11428 12590
rect 11488 12630 11548 12650
rect 11488 12590 11498 12630
rect 11538 12590 11548 12630
rect 11488 12570 11548 12590
rect 11608 12630 11668 12650
rect 11608 12590 11618 12630
rect 11658 12590 11668 12630
rect 11608 12570 11668 12590
rect 11728 12630 11788 12650
rect 11728 12590 11738 12630
rect 11778 12590 11788 12630
rect 11728 12570 11788 12590
rect 11848 12630 11908 12650
rect 11848 12590 11858 12630
rect 11898 12590 11908 12630
rect 11848 12570 11908 12590
rect 11968 12630 12028 12650
rect 11968 12590 11978 12630
rect 12018 12590 12028 12630
rect 11968 12570 12028 12590
rect 12088 12630 12148 12650
rect 12088 12590 12098 12630
rect 12138 12590 12148 12630
rect 12088 12570 12148 12590
rect 12208 12630 12268 12650
rect 12208 12590 12218 12630
rect 12258 12590 12268 12630
rect 12208 12570 12268 12590
rect 12328 12630 12388 12650
rect 12328 12590 12338 12630
rect 12378 12590 12388 12630
rect 12328 12570 12388 12590
rect 12448 12630 12508 12650
rect 12448 12590 12458 12630
rect 12498 12590 12508 12630
rect 12448 12570 12508 12590
rect 12568 12630 12628 12650
rect 12568 12590 12578 12630
rect 12618 12590 12628 12630
rect 12568 12570 12628 12590
rect 12798 12590 12808 12650
rect 12868 12590 12878 12650
rect 12798 12570 12878 12590
rect 11530 12522 11588 12530
rect 11530 12470 11534 12522
rect 11586 12470 11588 12522
rect 11530 12460 11588 12470
rect 11618 12430 11658 12570
rect 11688 12522 11746 12530
rect 11688 12470 11692 12522
rect 11744 12470 11746 12522
rect 11688 12460 11746 12470
rect 11598 12420 11678 12430
rect 11598 12360 11608 12420
rect 11668 12360 11678 12420
rect 11358 12310 11438 12320
rect 11358 12250 11368 12310
rect 11428 12250 11438 12310
rect 10618 12040 10778 12050
rect 10618 11980 10628 12040
rect 10688 11980 10708 12040
rect 10768 11980 10778 12040
rect 10618 11970 10778 11980
rect 11118 12040 11198 12050
rect 11118 11980 11128 12040
rect 11188 11980 11198 12040
rect 11118 11970 11198 11980
rect 11358 12040 11438 12250
rect 11358 11980 11368 12040
rect 11428 11980 11438 12040
rect 11358 11970 11438 11980
rect 10708 11920 10768 11970
rect 10708 11880 10718 11920
rect 10758 11880 10768 11920
rect 10708 11860 10768 11880
rect 10878 11920 10958 11930
rect 10878 11860 10888 11920
rect 10948 11860 10958 11920
rect 10878 11850 10958 11860
rect 10528 11790 10588 11810
rect 10528 11750 10538 11790
rect 10578 11750 10588 11790
rect 10528 11690 10588 11750
rect 10528 11650 10538 11690
rect 10578 11650 10588 11690
rect 10528 11570 10588 11650
rect 10648 11790 10708 11810
rect 10648 11750 10658 11790
rect 10698 11750 10708 11790
rect 10648 11690 10708 11750
rect 10648 11650 10658 11690
rect 10698 11650 10708 11690
rect 10648 11590 10708 11650
rect 10768 11790 10828 11810
rect 10768 11750 10778 11790
rect 10818 11750 10828 11790
rect 10768 11690 10828 11750
rect 10768 11650 10778 11690
rect 10818 11650 10828 11690
rect 10528 11530 10538 11570
rect 10578 11530 10588 11570
rect 10528 11480 10588 11530
rect 10638 11580 10718 11590
rect 10638 11520 10648 11580
rect 10708 11520 10718 11580
rect 10638 11510 10718 11520
rect 10768 11480 10828 11650
rect 10888 11790 10948 11850
rect 10888 11750 10898 11790
rect 10938 11750 10948 11790
rect 10888 11690 10948 11750
rect 10888 11650 10898 11690
rect 10938 11650 10948 11690
rect 10888 11630 10948 11650
rect 11008 11790 11068 11810
rect 11008 11750 11018 11790
rect 11058 11750 11068 11790
rect 11008 11690 11068 11750
rect 11008 11650 11018 11690
rect 11058 11650 11068 11690
rect 11008 11480 11068 11650
rect 11128 11790 11188 11970
rect 11368 11910 11428 11970
rect 11368 11870 11378 11910
rect 11418 11870 11428 11910
rect 11368 11850 11428 11870
rect 11598 11920 11678 12360
rect 11858 12320 11898 12570
rect 12012 12522 12070 12530
rect 12012 12470 12016 12522
rect 12068 12470 12070 12522
rect 12012 12460 12070 12470
rect 12098 12430 12138 12570
rect 12166 12522 12224 12530
rect 12166 12470 12170 12522
rect 12222 12470 12224 12522
rect 12166 12460 12224 12470
rect 12078 12420 12158 12430
rect 12078 12360 12088 12420
rect 12148 12360 12158 12420
rect 12078 12350 12158 12360
rect 12338 12320 12378 12570
rect 12490 12522 12548 12530
rect 12490 12470 12494 12522
rect 12546 12470 12548 12522
rect 12490 12460 12548 12470
rect 12578 12430 12618 12570
rect 12798 12510 12808 12570
rect 12868 12510 12878 12570
rect 12798 12500 12878 12510
rect 12558 12420 12638 12430
rect 12558 12360 12568 12420
rect 12628 12360 12638 12420
rect 12558 12350 12638 12360
rect 11838 12310 11918 12320
rect 11838 12250 11848 12310
rect 11908 12250 11918 12310
rect 11838 12240 11918 12250
rect 12318 12310 12398 12320
rect 12318 12250 12328 12310
rect 12388 12250 12398 12310
rect 12318 12240 12398 12250
rect 11838 12040 11918 12050
rect 11838 11980 11848 12040
rect 11908 11980 11918 12040
rect 11838 11970 11918 11980
rect 12078 12040 12158 12050
rect 12078 11980 12088 12040
rect 12148 11980 12158 12040
rect 12078 11970 12158 11980
rect 12558 12040 12638 12050
rect 12558 11980 12568 12040
rect 12628 11980 12638 12040
rect 12558 11970 12638 11980
rect 12738 12040 12818 12050
rect 12738 11980 12748 12040
rect 12808 11980 12818 12040
rect 12738 11970 12818 11980
rect 11598 11860 11608 11920
rect 11668 11860 11678 11920
rect 11598 11850 11678 11860
rect 11128 11750 11138 11790
rect 11178 11750 11188 11790
rect 11128 11690 11188 11750
rect 11128 11650 11138 11690
rect 11178 11650 11188 11690
rect 11128 11630 11188 11650
rect 11248 11790 11308 11810
rect 11248 11750 11258 11790
rect 11298 11750 11308 11790
rect 11248 11690 11308 11750
rect 11248 11650 11258 11690
rect 11298 11650 11308 11690
rect 11248 11480 11308 11650
rect 11368 11790 11428 11810
rect 11368 11750 11378 11790
rect 11418 11750 11428 11790
rect 11368 11690 11428 11750
rect 11368 11650 11378 11690
rect 11418 11650 11428 11690
rect 11368 11590 11428 11650
rect 11488 11790 11548 11810
rect 11488 11750 11498 11790
rect 11538 11750 11548 11790
rect 11488 11690 11548 11750
rect 11488 11650 11498 11690
rect 11538 11650 11548 11690
rect 11358 11580 11438 11590
rect 11358 11520 11368 11580
rect 11428 11520 11438 11580
rect 11358 11510 11438 11520
rect 11488 11480 11548 11650
rect 11608 11790 11668 11850
rect 11608 11750 11618 11790
rect 11658 11750 11668 11790
rect 11608 11690 11668 11750
rect 11608 11650 11618 11690
rect 11658 11650 11668 11690
rect 11608 11630 11668 11650
rect 11728 11790 11788 11810
rect 11728 11750 11738 11790
rect 11778 11750 11788 11790
rect 11728 11690 11788 11750
rect 11728 11650 11738 11690
rect 11778 11650 11788 11690
rect 11728 11480 11788 11650
rect 11848 11790 11908 11970
rect 12088 11910 12148 11970
rect 12088 11870 12098 11910
rect 12138 11870 12148 11910
rect 12088 11850 12148 11870
rect 12318 11920 12398 11930
rect 12318 11860 12328 11920
rect 12388 11860 12398 11920
rect 12318 11850 12398 11860
rect 11848 11750 11858 11790
rect 11898 11750 11908 11790
rect 11848 11690 11908 11750
rect 11848 11650 11858 11690
rect 11898 11650 11908 11690
rect 11848 11630 11908 11650
rect 11968 11790 12028 11810
rect 11968 11750 11978 11790
rect 12018 11750 12028 11790
rect 11968 11690 12028 11750
rect 11968 11650 11978 11690
rect 12018 11650 12028 11690
rect 11968 11480 12028 11650
rect 12088 11790 12148 11810
rect 12088 11750 12098 11790
rect 12138 11750 12148 11790
rect 12088 11690 12148 11750
rect 12088 11650 12098 11690
rect 12138 11650 12148 11690
rect 12088 11590 12148 11650
rect 12208 11790 12268 11810
rect 12208 11750 12218 11790
rect 12258 11750 12268 11790
rect 12208 11690 12268 11750
rect 12208 11650 12218 11690
rect 12258 11650 12268 11690
rect 12078 11580 12158 11590
rect 12078 11520 12088 11580
rect 12148 11520 12158 11580
rect 12078 11510 12158 11520
rect 12208 11480 12268 11650
rect 12328 11790 12388 11850
rect 12328 11750 12338 11790
rect 12378 11750 12388 11790
rect 12328 11690 12388 11750
rect 12328 11650 12338 11690
rect 12378 11650 12388 11690
rect 12328 11630 12388 11650
rect 12448 11790 12508 11810
rect 12448 11750 12458 11790
rect 12498 11750 12508 11790
rect 12448 11690 12508 11750
rect 12448 11650 12458 11690
rect 12498 11650 12508 11690
rect 12448 11480 12508 11650
rect 12568 11790 12628 11970
rect 12748 11910 12808 11970
rect 12748 11870 12758 11910
rect 12798 11870 12808 11910
rect 12748 11850 12808 11870
rect 12568 11750 12578 11790
rect 12618 11750 12628 11790
rect 12568 11690 12628 11750
rect 12568 11650 12578 11690
rect 12618 11650 12628 11690
rect 12568 11630 12628 11650
rect 12688 11790 12748 11810
rect 12688 11750 12698 11790
rect 12738 11750 12748 11790
rect 12688 11690 12748 11750
rect 12688 11650 12698 11690
rect 12738 11650 12748 11690
rect 12688 11480 12748 11650
rect 12808 11790 12868 11810
rect 12808 11750 12818 11790
rect 12858 11750 12868 11790
rect 12808 11690 12868 11750
rect 12808 11650 12818 11690
rect 12858 11650 12868 11690
rect 12808 11590 12868 11650
rect 12928 11790 12988 11810
rect 12928 11750 12938 11790
rect 12978 11750 12988 11790
rect 12928 11690 12988 11750
rect 12928 11650 12938 11690
rect 12978 11650 12988 11690
rect 12798 11580 12878 11590
rect 12798 11520 12808 11580
rect 12868 11520 12878 11580
rect 12798 11510 12878 11520
rect 12928 11570 12988 11650
rect 13068 11590 13128 13110
rect 13158 12730 13398 13710
rect 14578 13930 14658 13940
rect 14578 13870 14588 13930
rect 14648 13870 14658 13930
rect 14578 13850 14658 13870
rect 14578 13790 14588 13850
rect 14648 13790 14658 13850
rect 14578 13770 14658 13790
rect 14578 13710 14588 13770
rect 14648 13710 14658 13770
rect 14578 13700 14658 13710
rect 15748 13640 15808 13660
rect 15748 13600 15758 13640
rect 15798 13600 15808 13640
rect 15748 13540 15808 13600
rect 15748 13500 15758 13540
rect 15798 13500 15808 13540
rect 15748 13440 15808 13500
rect 15748 13400 15758 13440
rect 15798 13400 15808 13440
rect 15748 13340 15808 13400
rect 15748 13300 15758 13340
rect 15798 13300 15808 13340
rect 15748 13240 15808 13300
rect 15748 13200 15758 13240
rect 15798 13200 15808 13240
rect 13158 12670 13168 12730
rect 13228 12670 13248 12730
rect 13308 12670 13328 12730
rect 13388 12670 13398 12730
rect 13158 12650 13398 12670
rect 13158 12590 13168 12650
rect 13228 12590 13248 12650
rect 13308 12590 13328 12650
rect 13388 12590 13398 12650
rect 13158 12570 13398 12590
rect 13158 12510 13168 12570
rect 13228 12510 13248 12570
rect 13308 12510 13328 12570
rect 13388 12510 13398 12570
rect 13158 12500 13398 12510
rect 13428 13150 13488 13170
rect 13428 13110 13438 13150
rect 13478 13110 13488 13150
rect 13428 11590 13488 13110
rect 13718 13130 13798 13140
rect 13718 13070 13728 13130
rect 13788 13070 13798 13130
rect 13718 13050 13798 13070
rect 13718 12990 13728 13050
rect 13788 12990 13798 13050
rect 13718 12970 13798 12990
rect 13718 12910 13728 12970
rect 13788 12910 13798 12970
rect 13718 12900 13798 12910
rect 13958 13130 14038 13140
rect 13958 13070 13968 13130
rect 14028 13070 14038 13130
rect 13958 13050 14038 13070
rect 13958 12990 13968 13050
rect 14028 12990 14038 13050
rect 13958 12970 14038 12990
rect 13958 12910 13968 12970
rect 14028 12910 14038 12970
rect 13958 12900 14038 12910
rect 14198 13130 14278 13140
rect 14198 13070 14208 13130
rect 14268 13070 14278 13130
rect 14198 13050 14278 13070
rect 14198 12990 14208 13050
rect 14268 12990 14278 13050
rect 14198 12970 14278 12990
rect 14198 12910 14208 12970
rect 14268 12910 14278 12970
rect 14198 12900 14278 12910
rect 14838 13130 14918 13140
rect 14838 13070 14848 13130
rect 14908 13070 14918 13130
rect 14838 13050 14918 13070
rect 14838 12990 14848 13050
rect 14908 12990 14918 13050
rect 14838 12970 14918 12990
rect 14838 12910 14848 12970
rect 14908 12910 14918 12970
rect 14838 12900 14918 12910
rect 15078 13130 15158 13140
rect 15078 13070 15088 13130
rect 15148 13070 15158 13130
rect 15078 13050 15158 13070
rect 15078 12990 15088 13050
rect 15148 12990 15158 13050
rect 15078 12970 15158 12990
rect 15078 12910 15088 12970
rect 15148 12910 15158 12970
rect 15078 12900 15158 12910
rect 15318 13130 15398 13140
rect 15318 13070 15328 13130
rect 15388 13070 15398 13130
rect 15318 13050 15398 13070
rect 15318 12990 15328 13050
rect 15388 12990 15398 13050
rect 15318 12970 15398 12990
rect 15318 12910 15328 12970
rect 15388 12910 15398 12970
rect 15318 12900 15398 12910
rect 15558 13130 15638 13140
rect 15558 13070 15568 13130
rect 15628 13070 15638 13130
rect 15558 13050 15638 13070
rect 15558 12990 15568 13050
rect 15628 12990 15638 13050
rect 15558 12970 15638 12990
rect 15558 12910 15568 12970
rect 15628 12910 15638 12970
rect 15558 12900 15638 12910
rect 15748 12870 15808 13200
rect 14028 12860 14108 12870
rect 14028 12800 14038 12860
rect 14098 12800 14108 12860
rect 14028 12790 14108 12800
rect 14288 12860 14368 12870
rect 14288 12800 14298 12860
rect 14358 12800 14368 12860
rect 14288 12790 14368 12800
rect 14508 12860 14588 12870
rect 14508 12800 14518 12860
rect 14578 12800 14588 12860
rect 14508 12790 14588 12800
rect 14768 12860 14848 12870
rect 14768 12800 14778 12860
rect 14838 12800 14848 12860
rect 14768 12790 14848 12800
rect 14988 12860 15068 12870
rect 14988 12800 14998 12860
rect 15058 12800 15068 12860
rect 14988 12790 15068 12800
rect 15738 12860 15818 12870
rect 15738 12800 15748 12860
rect 15808 12800 15818 12860
rect 15738 12790 15818 12800
rect 13678 12730 13758 12740
rect 13678 12670 13688 12730
rect 13748 12670 13758 12730
rect 13678 12650 13758 12670
rect 14048 12650 14078 12790
rect 14109 12750 14167 12760
rect 14109 12698 14113 12750
rect 14165 12698 14167 12750
rect 14109 12690 14167 12698
rect 14229 12750 14287 12760
rect 14229 12698 14233 12750
rect 14285 12698 14287 12750
rect 14229 12690 14287 12698
rect 14318 12650 14348 12790
rect 14528 12650 14558 12790
rect 14589 12750 14647 12760
rect 14589 12698 14593 12750
rect 14645 12698 14647 12750
rect 14589 12690 14647 12698
rect 14709 12750 14767 12760
rect 14709 12698 14713 12750
rect 14765 12698 14767 12750
rect 14709 12690 14767 12698
rect 14798 12650 14828 12790
rect 15008 12650 15038 12790
rect 16168 12760 16208 14530
rect 15069 12750 15127 12760
rect 15069 12698 15073 12750
rect 15125 12698 15127 12750
rect 15069 12690 15127 12698
rect 16148 12750 16228 12760
rect 16148 12690 16158 12750
rect 16218 12690 16228 12750
rect 16148 12680 16228 12690
rect 13678 12590 13688 12650
rect 13748 12590 13758 12650
rect 13678 12570 13758 12590
rect 13928 12630 13988 12650
rect 13928 12590 13938 12630
rect 13978 12590 13988 12630
rect 13928 12570 13988 12590
rect 14048 12630 14108 12650
rect 14048 12590 14058 12630
rect 14098 12590 14108 12630
rect 14048 12570 14108 12590
rect 14168 12630 14228 12650
rect 14168 12590 14178 12630
rect 14218 12590 14228 12630
rect 14168 12570 14228 12590
rect 14288 12630 14348 12650
rect 14288 12590 14298 12630
rect 14338 12590 14348 12630
rect 14288 12570 14348 12590
rect 14408 12630 14468 12650
rect 14408 12590 14418 12630
rect 14458 12590 14468 12630
rect 14408 12570 14468 12590
rect 14528 12630 14588 12650
rect 14528 12590 14538 12630
rect 14578 12590 14588 12630
rect 14528 12570 14588 12590
rect 14648 12630 14708 12650
rect 14648 12590 14658 12630
rect 14698 12590 14708 12630
rect 14648 12570 14708 12590
rect 14768 12630 14828 12650
rect 14768 12590 14778 12630
rect 14818 12590 14828 12630
rect 14768 12570 14828 12590
rect 14888 12630 14948 12650
rect 14888 12590 14898 12630
rect 14938 12590 14948 12630
rect 14888 12570 14948 12590
rect 15008 12630 15068 12650
rect 15008 12590 15018 12630
rect 15058 12590 15068 12630
rect 15008 12570 15068 12590
rect 15128 12630 15188 12650
rect 15128 12590 15138 12630
rect 15178 12590 15188 12630
rect 13678 12510 13688 12570
rect 13748 12510 13758 12570
rect 13678 12500 13758 12510
rect 13938 12430 13978 12570
rect 14008 12522 14066 12530
rect 14008 12470 14010 12522
rect 14062 12470 14066 12522
rect 14008 12460 14066 12470
rect 13918 12420 13998 12430
rect 13918 12360 13928 12420
rect 13988 12360 13998 12420
rect 13918 12350 13998 12360
rect 14178 12320 14218 12570
rect 14332 12522 14390 12530
rect 14332 12470 14334 12522
rect 14386 12470 14390 12522
rect 14332 12460 14390 12470
rect 14418 12430 14458 12570
rect 14486 12522 14544 12530
rect 14486 12470 14488 12522
rect 14540 12470 14544 12522
rect 14486 12460 14544 12470
rect 14398 12420 14478 12430
rect 14398 12360 14408 12420
rect 14468 12360 14478 12420
rect 14398 12350 14478 12360
rect 14658 12320 14698 12570
rect 14810 12522 14868 12530
rect 14810 12470 14812 12522
rect 14864 12470 14868 12522
rect 14810 12460 14868 12470
rect 14898 12430 14938 12570
rect 14968 12522 15026 12530
rect 14968 12470 14970 12522
rect 15022 12470 15026 12522
rect 14968 12460 15026 12470
rect 14878 12420 14958 12430
rect 14878 12360 14888 12420
rect 14948 12360 14958 12420
rect 14158 12310 14238 12320
rect 14158 12250 14168 12310
rect 14228 12250 14238 12310
rect 14158 12240 14238 12250
rect 14638 12310 14718 12320
rect 14638 12250 14648 12310
rect 14708 12250 14718 12310
rect 14638 12240 14718 12250
rect 13738 12200 13818 12210
rect 13738 12140 13748 12200
rect 13808 12140 13818 12200
rect 13738 12120 13818 12140
rect 13738 12060 13748 12120
rect 13808 12060 13818 12120
rect 13738 12040 13818 12060
rect 13738 11980 13748 12040
rect 13808 11980 13818 12040
rect 13738 11970 13818 11980
rect 13918 12200 13998 12210
rect 13918 12140 13928 12200
rect 13988 12140 13998 12200
rect 13918 12120 13998 12140
rect 13918 12060 13928 12120
rect 13988 12060 13998 12120
rect 13918 12040 13998 12060
rect 13918 11980 13928 12040
rect 13988 11980 13998 12040
rect 13918 11970 13998 11980
rect 14158 12200 14238 12210
rect 14158 12140 14168 12200
rect 14228 12140 14238 12200
rect 14158 12120 14238 12140
rect 14158 12060 14168 12120
rect 14228 12060 14238 12120
rect 14158 12040 14238 12060
rect 14158 11980 14168 12040
rect 14228 11980 14238 12040
rect 14158 11970 14238 11980
rect 14398 12200 14478 12210
rect 14398 12140 14408 12200
rect 14468 12140 14478 12200
rect 14398 12120 14478 12140
rect 14398 12060 14408 12120
rect 14468 12060 14478 12120
rect 14398 12040 14478 12060
rect 14398 11980 14408 12040
rect 14468 11980 14478 12040
rect 14398 11970 14478 11980
rect 14638 12200 14718 12210
rect 14638 12140 14648 12200
rect 14708 12140 14718 12200
rect 14638 12120 14718 12140
rect 14638 12060 14648 12120
rect 14708 12060 14718 12120
rect 14638 12040 14718 12060
rect 14638 11980 14648 12040
rect 14708 11980 14718 12040
rect 14638 11970 14718 11980
rect 13748 11910 13808 11970
rect 13748 11870 13758 11910
rect 13798 11870 13808 11910
rect 13748 11850 13808 11870
rect 13568 11790 13628 11810
rect 13568 11750 13578 11790
rect 13618 11750 13628 11790
rect 13568 11690 13628 11750
rect 13568 11650 13578 11690
rect 13618 11650 13628 11690
rect 12928 11530 12938 11570
rect 12978 11530 12988 11570
rect 12928 11480 12988 11530
rect 13058 11580 13138 11590
rect 13058 11520 13068 11580
rect 13128 11520 13138 11580
rect 13058 11510 13138 11520
rect 13418 11580 13498 11590
rect 13418 11520 13428 11580
rect 13488 11520 13498 11580
rect 10518 11470 10598 11480
rect 10518 11410 10528 11470
rect 10588 11410 10598 11470
rect 10518 11390 10598 11410
rect 10518 11330 10528 11390
rect 10588 11330 10598 11390
rect 10518 11310 10598 11330
rect 10518 11250 10528 11310
rect 10588 11250 10598 11310
rect 10518 11240 10598 11250
rect 10758 11470 10838 11480
rect 10758 11410 10768 11470
rect 10828 11410 10838 11470
rect 10758 11390 10838 11410
rect 10758 11330 10768 11390
rect 10828 11330 10838 11390
rect 10758 11310 10838 11330
rect 10758 11250 10768 11310
rect 10828 11250 10838 11310
rect 10758 11240 10838 11250
rect 10998 11470 11078 11480
rect 10998 11410 11008 11470
rect 11068 11410 11078 11470
rect 10998 11390 11078 11410
rect 10998 11330 11008 11390
rect 11068 11330 11078 11390
rect 10998 11310 11078 11330
rect 10998 11250 11008 11310
rect 11068 11250 11078 11310
rect 10998 11240 11078 11250
rect 11238 11470 11318 11480
rect 11238 11410 11248 11470
rect 11308 11410 11318 11470
rect 11238 11390 11318 11410
rect 11238 11330 11248 11390
rect 11308 11330 11318 11390
rect 11238 11310 11318 11330
rect 11238 11250 11248 11310
rect 11308 11250 11318 11310
rect 11238 11240 11318 11250
rect 11478 11470 11558 11480
rect 11478 11410 11488 11470
rect 11548 11410 11558 11470
rect 11478 11390 11558 11410
rect 11478 11330 11488 11390
rect 11548 11330 11558 11390
rect 11478 11310 11558 11330
rect 11478 11250 11488 11310
rect 11548 11250 11558 11310
rect 11478 11240 11558 11250
rect 11718 11470 11798 11480
rect 11718 11410 11728 11470
rect 11788 11410 11798 11470
rect 11718 11390 11798 11410
rect 11718 11330 11728 11390
rect 11788 11330 11798 11390
rect 11718 11310 11798 11330
rect 11718 11250 11728 11310
rect 11788 11250 11798 11310
rect 11718 11240 11798 11250
rect 11958 11470 12038 11480
rect 11958 11410 11968 11470
rect 12028 11410 12038 11470
rect 11958 11390 12038 11410
rect 11958 11330 11968 11390
rect 12028 11330 12038 11390
rect 11958 11310 12038 11330
rect 11958 11250 11968 11310
rect 12028 11250 12038 11310
rect 11958 11240 12038 11250
rect 12198 11470 12278 11480
rect 12198 11410 12208 11470
rect 12268 11410 12278 11470
rect 12198 11390 12278 11410
rect 12198 11330 12208 11390
rect 12268 11330 12278 11390
rect 12198 11310 12278 11330
rect 12198 11250 12208 11310
rect 12268 11250 12278 11310
rect 12198 11240 12278 11250
rect 12438 11470 12518 11480
rect 12438 11410 12448 11470
rect 12508 11410 12518 11470
rect 12438 11390 12518 11410
rect 12438 11330 12448 11390
rect 12508 11330 12518 11390
rect 12438 11310 12518 11330
rect 12438 11250 12448 11310
rect 12508 11250 12518 11310
rect 12438 11240 12518 11250
rect 12678 11470 12758 11480
rect 12678 11410 12688 11470
rect 12748 11410 12758 11470
rect 12678 11390 12758 11410
rect 12678 11330 12688 11390
rect 12748 11330 12758 11390
rect 12678 11310 12758 11330
rect 12678 11250 12688 11310
rect 12748 11250 12758 11310
rect 12678 11240 12758 11250
rect 12918 11470 12998 11480
rect 12918 11410 12928 11470
rect 12988 11410 12998 11470
rect 12918 11390 12998 11410
rect 12918 11330 12928 11390
rect 12988 11330 12998 11390
rect 12918 11310 12998 11330
rect 12918 11250 12928 11310
rect 12988 11250 12998 11310
rect 12918 11240 12998 11250
rect 11798 11200 11878 11210
rect 11798 11140 11808 11200
rect 11868 11140 11878 11200
rect 11798 11130 11878 11140
rect 13238 11200 13318 11210
rect 13238 11140 13248 11200
rect 13308 11140 13318 11200
rect 13238 11130 13318 11140
rect 11628 10630 11688 10650
rect 11628 10590 11638 10630
rect 11678 10590 11688 10630
rect 11628 10530 11688 10590
rect 11628 10490 11638 10530
rect 11678 10490 11688 10530
rect 11628 10430 11688 10490
rect 11628 10390 11638 10430
rect 11678 10390 11688 10430
rect 11628 10330 11688 10390
rect 11628 10290 11638 10330
rect 11678 10290 11688 10330
rect 11628 10230 11688 10290
rect 11628 10190 11638 10230
rect 11678 10190 11688 10230
rect 11628 10130 11688 10190
rect 11628 10090 11638 10130
rect 11678 10090 11688 10130
rect 11628 10070 11688 10090
rect 11808 10630 11868 11130
rect 12158 11090 12238 11100
rect 12158 11030 12168 11090
rect 12228 11030 12238 11090
rect 12158 11020 12238 11030
rect 11898 10760 11968 10770
rect 11958 10700 11968 10760
rect 11898 10690 11968 10700
rect 12068 10760 12148 10770
rect 12068 10700 12078 10760
rect 12138 10700 12148 10760
rect 12068 10690 12148 10700
rect 12178 10650 12218 11020
rect 12518 10980 12598 10990
rect 12518 10920 12528 10980
rect 12588 10920 12598 10980
rect 12518 10910 12598 10920
rect 12248 10760 12328 10770
rect 12248 10700 12258 10760
rect 12318 10700 12328 10760
rect 12248 10690 12328 10700
rect 12428 10760 12508 10770
rect 12428 10700 12438 10760
rect 12498 10700 12508 10760
rect 12428 10690 12508 10700
rect 12538 10650 12578 10910
rect 12878 10870 12958 10880
rect 12878 10810 12888 10870
rect 12948 10810 12958 10870
rect 12878 10800 12958 10810
rect 12608 10760 12688 10770
rect 12608 10700 12618 10760
rect 12678 10700 12688 10760
rect 12608 10690 12688 10700
rect 12788 10760 12868 10770
rect 12788 10700 12798 10760
rect 12858 10700 12868 10760
rect 12788 10690 12868 10700
rect 12898 10650 12938 10800
rect 12968 10760 13048 10770
rect 12968 10700 12978 10760
rect 13038 10700 13048 10760
rect 12968 10690 13048 10700
rect 13148 10760 13218 10770
rect 13148 10700 13158 10760
rect 13148 10690 13218 10700
rect 11808 10590 11818 10630
rect 11858 10590 11868 10630
rect 11808 10530 11868 10590
rect 11808 10490 11818 10530
rect 11858 10490 11868 10530
rect 11808 10430 11868 10490
rect 11808 10390 11818 10430
rect 11858 10390 11868 10430
rect 11808 10330 11868 10390
rect 11808 10290 11818 10330
rect 11858 10290 11868 10330
rect 11808 10230 11868 10290
rect 11808 10190 11818 10230
rect 11858 10190 11868 10230
rect 11808 10130 11868 10190
rect 11808 10090 11818 10130
rect 11858 10090 11868 10130
rect 11808 10070 11868 10090
rect 11988 10630 12048 10650
rect 11988 10590 11998 10630
rect 12038 10590 12048 10630
rect 11988 10530 12048 10590
rect 11988 10490 11998 10530
rect 12038 10490 12048 10530
rect 11988 10430 12048 10490
rect 11988 10390 11998 10430
rect 12038 10390 12048 10430
rect 11988 10330 12048 10390
rect 11988 10290 11998 10330
rect 12038 10290 12048 10330
rect 11988 10230 12048 10290
rect 11988 10190 11998 10230
rect 12038 10190 12048 10230
rect 11988 10130 12048 10190
rect 11988 10090 11998 10130
rect 12038 10090 12048 10130
rect 11988 10070 12048 10090
rect 12168 10630 12228 10650
rect 12168 10590 12178 10630
rect 12218 10590 12228 10630
rect 12168 10530 12228 10590
rect 12168 10490 12178 10530
rect 12218 10490 12228 10530
rect 12168 10430 12228 10490
rect 12168 10390 12178 10430
rect 12218 10390 12228 10430
rect 12168 10330 12228 10390
rect 12168 10290 12178 10330
rect 12218 10290 12228 10330
rect 12168 10230 12228 10290
rect 12168 10190 12178 10230
rect 12218 10190 12228 10230
rect 12168 10130 12228 10190
rect 12168 10090 12178 10130
rect 12218 10090 12228 10130
rect 12168 10070 12228 10090
rect 12348 10630 12408 10650
rect 12348 10590 12358 10630
rect 12398 10590 12408 10630
rect 12348 10530 12408 10590
rect 12348 10490 12358 10530
rect 12398 10490 12408 10530
rect 12348 10430 12408 10490
rect 12348 10390 12358 10430
rect 12398 10390 12408 10430
rect 12348 10330 12408 10390
rect 12348 10290 12358 10330
rect 12398 10290 12408 10330
rect 12348 10230 12408 10290
rect 12348 10190 12358 10230
rect 12398 10190 12408 10230
rect 12348 10130 12408 10190
rect 12348 10090 12358 10130
rect 12398 10090 12408 10130
rect 12348 10070 12408 10090
rect 12528 10630 12588 10650
rect 12528 10590 12538 10630
rect 12578 10590 12588 10630
rect 12528 10530 12588 10590
rect 12528 10490 12538 10530
rect 12578 10490 12588 10530
rect 12528 10430 12588 10490
rect 12528 10390 12538 10430
rect 12578 10390 12588 10430
rect 12528 10330 12588 10390
rect 12528 10290 12538 10330
rect 12578 10290 12588 10330
rect 12528 10230 12588 10290
rect 12528 10190 12538 10230
rect 12578 10190 12588 10230
rect 12528 10130 12588 10190
rect 12528 10090 12538 10130
rect 12578 10090 12588 10130
rect 12528 10070 12588 10090
rect 12708 10630 12768 10650
rect 12708 10590 12718 10630
rect 12758 10590 12768 10630
rect 12708 10530 12768 10590
rect 12708 10490 12718 10530
rect 12758 10490 12768 10530
rect 12708 10430 12768 10490
rect 12708 10390 12718 10430
rect 12758 10390 12768 10430
rect 12708 10330 12768 10390
rect 12708 10290 12718 10330
rect 12758 10290 12768 10330
rect 12708 10230 12768 10290
rect 12708 10190 12718 10230
rect 12758 10190 12768 10230
rect 12708 10130 12768 10190
rect 12708 10090 12718 10130
rect 12758 10090 12768 10130
rect 12708 10070 12768 10090
rect 12888 10630 12948 10650
rect 12888 10590 12898 10630
rect 12938 10590 12948 10630
rect 12888 10530 12948 10590
rect 12888 10490 12898 10530
rect 12938 10490 12948 10530
rect 12888 10430 12948 10490
rect 12888 10390 12898 10430
rect 12938 10390 12948 10430
rect 12888 10330 12948 10390
rect 12888 10290 12898 10330
rect 12938 10290 12948 10330
rect 12888 10230 12948 10290
rect 12888 10190 12898 10230
rect 12938 10190 12948 10230
rect 12888 10130 12948 10190
rect 12888 10090 12898 10130
rect 12938 10090 12948 10130
rect 12888 10070 12948 10090
rect 13068 10630 13128 10650
rect 13068 10590 13078 10630
rect 13118 10590 13128 10630
rect 13068 10530 13128 10590
rect 13068 10490 13078 10530
rect 13118 10490 13128 10530
rect 13068 10430 13128 10490
rect 13068 10390 13078 10430
rect 13118 10390 13128 10430
rect 13068 10330 13128 10390
rect 13068 10290 13078 10330
rect 13118 10290 13128 10330
rect 13068 10230 13128 10290
rect 13068 10190 13078 10230
rect 13118 10190 13128 10230
rect 13068 10130 13128 10190
rect 13068 10090 13078 10130
rect 13118 10090 13128 10130
rect 13068 10070 13128 10090
rect 13248 10630 13308 11130
rect 13418 10770 13498 11520
rect 13568 11570 13628 11650
rect 13688 11790 13748 11810
rect 13688 11750 13698 11790
rect 13738 11750 13748 11790
rect 13688 11690 13748 11750
rect 13688 11650 13698 11690
rect 13738 11650 13748 11690
rect 13688 11590 13748 11650
rect 13808 11790 13868 11810
rect 13808 11750 13818 11790
rect 13858 11750 13868 11790
rect 13808 11690 13868 11750
rect 13808 11650 13818 11690
rect 13858 11650 13868 11690
rect 13568 11530 13578 11570
rect 13618 11530 13628 11570
rect 13568 11480 13628 11530
rect 13678 11580 13758 11590
rect 13678 11520 13688 11580
rect 13748 11520 13758 11580
rect 13678 11510 13758 11520
rect 13808 11480 13868 11650
rect 13928 11790 13988 11970
rect 14158 11920 14238 11930
rect 14158 11860 14168 11920
rect 14228 11860 14238 11920
rect 14158 11850 14238 11860
rect 14408 11910 14468 11970
rect 14408 11870 14418 11910
rect 14458 11870 14468 11910
rect 14408 11850 14468 11870
rect 13928 11750 13938 11790
rect 13978 11750 13988 11790
rect 13928 11690 13988 11750
rect 13928 11650 13938 11690
rect 13978 11650 13988 11690
rect 13928 11630 13988 11650
rect 14048 11790 14108 11810
rect 14048 11750 14058 11790
rect 14098 11750 14108 11790
rect 14048 11690 14108 11750
rect 14048 11650 14058 11690
rect 14098 11650 14108 11690
rect 14048 11480 14108 11650
rect 14168 11790 14228 11850
rect 14168 11750 14178 11790
rect 14218 11750 14228 11790
rect 14168 11690 14228 11750
rect 14168 11650 14178 11690
rect 14218 11650 14228 11690
rect 14168 11630 14228 11650
rect 14288 11790 14348 11810
rect 14288 11750 14298 11790
rect 14338 11750 14348 11790
rect 14288 11690 14348 11750
rect 14288 11650 14298 11690
rect 14338 11650 14348 11690
rect 14288 11480 14348 11650
rect 14408 11790 14468 11810
rect 14408 11750 14418 11790
rect 14458 11750 14468 11790
rect 14408 11690 14468 11750
rect 14408 11650 14418 11690
rect 14458 11650 14468 11690
rect 14408 11590 14468 11650
rect 14528 11790 14588 11810
rect 14528 11750 14538 11790
rect 14578 11750 14588 11790
rect 14528 11690 14588 11750
rect 14528 11650 14538 11690
rect 14578 11650 14588 11690
rect 14398 11580 14478 11590
rect 14398 11520 14408 11580
rect 14468 11520 14478 11580
rect 14398 11510 14478 11520
rect 14528 11480 14588 11650
rect 14648 11790 14708 11970
rect 14878 11920 14958 12360
rect 15128 12320 15188 12590
rect 15118 12310 15198 12320
rect 15118 12250 15128 12310
rect 15188 12250 15198 12310
rect 15118 12200 15198 12250
rect 15118 12140 15128 12200
rect 15188 12140 15198 12200
rect 15118 12120 15198 12140
rect 15118 12060 15128 12120
rect 15188 12060 15198 12120
rect 15118 12040 15198 12060
rect 15118 11980 15128 12040
rect 15188 11980 15198 12040
rect 15118 11970 15198 11980
rect 15358 12200 15438 12210
rect 15358 12140 15368 12200
rect 15428 12140 15438 12200
rect 15358 12120 15438 12140
rect 15358 12060 15368 12120
rect 15428 12060 15438 12120
rect 15358 12040 15438 12060
rect 15358 11980 15368 12040
rect 15428 11980 15438 12040
rect 15358 11970 15438 11980
rect 15778 12200 15858 12210
rect 15778 12140 15788 12200
rect 15848 12140 15858 12200
rect 15778 12120 15858 12140
rect 15778 12060 15788 12120
rect 15848 12060 15858 12120
rect 15778 12040 15858 12060
rect 15778 11980 15788 12040
rect 15848 11980 15858 12040
rect 15778 11970 15858 11980
rect 14878 11860 14888 11920
rect 14948 11860 14958 11920
rect 14878 11850 14958 11860
rect 15128 11910 15188 11970
rect 15128 11870 15138 11910
rect 15178 11870 15188 11910
rect 15128 11850 15188 11870
rect 14648 11750 14658 11790
rect 14698 11750 14708 11790
rect 14648 11690 14708 11750
rect 14648 11650 14658 11690
rect 14698 11650 14708 11690
rect 14648 11630 14708 11650
rect 14768 11790 14828 11810
rect 14768 11750 14778 11790
rect 14818 11750 14828 11790
rect 14768 11690 14828 11750
rect 14768 11650 14778 11690
rect 14818 11650 14828 11690
rect 14768 11480 14828 11650
rect 14888 11790 14948 11850
rect 14888 11750 14898 11790
rect 14938 11750 14948 11790
rect 14888 11690 14948 11750
rect 14888 11650 14898 11690
rect 14938 11650 14948 11690
rect 14888 11630 14948 11650
rect 15008 11790 15068 11810
rect 15008 11750 15018 11790
rect 15058 11750 15068 11790
rect 15008 11690 15068 11750
rect 15008 11650 15018 11690
rect 15058 11650 15068 11690
rect 15008 11480 15068 11650
rect 15128 11790 15188 11810
rect 15128 11750 15138 11790
rect 15178 11750 15188 11790
rect 15128 11690 15188 11750
rect 15128 11650 15138 11690
rect 15178 11650 15188 11690
rect 15128 11590 15188 11650
rect 15248 11790 15308 11810
rect 15248 11750 15258 11790
rect 15298 11750 15308 11790
rect 15248 11690 15308 11750
rect 15248 11650 15258 11690
rect 15298 11650 15308 11690
rect 15118 11580 15198 11590
rect 15118 11520 15128 11580
rect 15188 11520 15198 11580
rect 15118 11510 15198 11520
rect 15248 11480 15308 11650
rect 15368 11790 15428 11970
rect 15598 11920 15678 11930
rect 15598 11860 15608 11920
rect 15668 11860 15678 11920
rect 15788 11920 15848 11970
rect 15788 11880 15798 11920
rect 15838 11880 15848 11920
rect 15788 11860 15848 11880
rect 15598 11850 15678 11860
rect 15368 11750 15378 11790
rect 15418 11750 15428 11790
rect 15368 11690 15428 11750
rect 15368 11650 15378 11690
rect 15418 11650 15428 11690
rect 15368 11630 15428 11650
rect 15488 11790 15548 11810
rect 15488 11750 15498 11790
rect 15538 11750 15548 11790
rect 15488 11690 15548 11750
rect 15488 11650 15498 11690
rect 15538 11650 15548 11690
rect 15488 11480 15548 11650
rect 15608 11790 15668 11850
rect 15608 11750 15618 11790
rect 15658 11750 15668 11790
rect 15608 11690 15668 11750
rect 15608 11650 15618 11690
rect 15658 11650 15668 11690
rect 15608 11630 15668 11650
rect 15728 11790 15788 11810
rect 15728 11750 15738 11790
rect 15778 11750 15788 11790
rect 15728 11690 15788 11750
rect 15728 11650 15738 11690
rect 15778 11650 15788 11690
rect 15728 11480 15788 11650
rect 15848 11790 15908 11810
rect 15848 11750 15858 11790
rect 15898 11750 15908 11790
rect 15848 11690 15908 11750
rect 15848 11650 15858 11690
rect 15898 11650 15908 11690
rect 15848 11590 15908 11650
rect 15968 11790 16028 11810
rect 15968 11750 15978 11790
rect 16018 11750 16028 11790
rect 15968 11690 16028 11750
rect 15968 11650 15978 11690
rect 16018 11650 16028 11690
rect 15838 11580 15918 11590
rect 15838 11520 15848 11580
rect 15908 11520 15918 11580
rect 13558 11470 13638 11480
rect 13558 11410 13568 11470
rect 13628 11410 13638 11470
rect 13558 11390 13638 11410
rect 13558 11330 13568 11390
rect 13628 11330 13638 11390
rect 13558 11310 13638 11330
rect 13558 11250 13568 11310
rect 13628 11250 13638 11310
rect 13558 11240 13638 11250
rect 13798 11470 13878 11480
rect 13798 11410 13808 11470
rect 13868 11410 13878 11470
rect 13798 11390 13878 11410
rect 13798 11330 13808 11390
rect 13868 11330 13878 11390
rect 13798 11310 13878 11330
rect 13798 11250 13808 11310
rect 13868 11250 13878 11310
rect 13798 11240 13878 11250
rect 14038 11470 14118 11480
rect 14038 11410 14048 11470
rect 14108 11410 14118 11470
rect 14038 11390 14118 11410
rect 14038 11330 14048 11390
rect 14108 11330 14118 11390
rect 14038 11310 14118 11330
rect 14038 11250 14048 11310
rect 14108 11250 14118 11310
rect 14038 11240 14118 11250
rect 14278 11470 14358 11480
rect 14278 11410 14288 11470
rect 14348 11410 14358 11470
rect 14278 11390 14358 11410
rect 14278 11330 14288 11390
rect 14348 11330 14358 11390
rect 14278 11310 14358 11330
rect 14278 11250 14288 11310
rect 14348 11250 14358 11310
rect 14278 11240 14358 11250
rect 14518 11470 14598 11480
rect 14518 11410 14528 11470
rect 14588 11410 14598 11470
rect 14518 11390 14598 11410
rect 14518 11330 14528 11390
rect 14588 11330 14598 11390
rect 14518 11310 14598 11330
rect 14518 11250 14528 11310
rect 14588 11250 14598 11310
rect 14518 11240 14598 11250
rect 14758 11470 14838 11480
rect 14758 11410 14768 11470
rect 14828 11410 14838 11470
rect 14758 11390 14838 11410
rect 14758 11330 14768 11390
rect 14828 11330 14838 11390
rect 14758 11310 14838 11330
rect 14758 11250 14768 11310
rect 14828 11250 14838 11310
rect 14758 11240 14838 11250
rect 14998 11470 15078 11480
rect 14998 11410 15008 11470
rect 15068 11410 15078 11470
rect 14998 11390 15078 11410
rect 14998 11330 15008 11390
rect 15068 11330 15078 11390
rect 14998 11310 15078 11330
rect 14998 11250 15008 11310
rect 15068 11250 15078 11310
rect 14998 11240 15078 11250
rect 15238 11470 15318 11480
rect 15238 11410 15248 11470
rect 15308 11410 15318 11470
rect 15238 11390 15318 11410
rect 15238 11330 15248 11390
rect 15308 11330 15318 11390
rect 15238 11310 15318 11330
rect 15238 11250 15248 11310
rect 15308 11250 15318 11310
rect 15238 11240 15318 11250
rect 15478 11470 15558 11480
rect 15478 11410 15488 11470
rect 15548 11410 15558 11470
rect 15478 11390 15558 11410
rect 15478 11330 15488 11390
rect 15548 11330 15558 11390
rect 15478 11310 15558 11330
rect 15478 11250 15488 11310
rect 15548 11250 15558 11310
rect 15478 11240 15558 11250
rect 15718 11470 15798 11480
rect 15718 11410 15728 11470
rect 15788 11410 15798 11470
rect 15718 11390 15798 11410
rect 15718 11330 15728 11390
rect 15788 11330 15798 11390
rect 15718 11310 15798 11330
rect 15718 11250 15728 11310
rect 15788 11250 15798 11310
rect 15718 11240 15798 11250
rect 14678 11200 14758 11210
rect 14678 11140 14688 11200
rect 14748 11140 14758 11200
rect 14678 11130 14758 11140
rect 14318 11090 14398 11100
rect 14318 11030 14328 11090
rect 14388 11030 14398 11090
rect 14318 11020 14398 11030
rect 13958 10980 14038 10990
rect 13958 10920 13968 10980
rect 14028 10920 14038 10980
rect 13958 10910 14038 10920
rect 13598 10870 13678 10880
rect 13598 10810 13608 10870
rect 13668 10810 13678 10870
rect 13598 10800 13678 10810
rect 13338 10760 13588 10770
rect 13398 10700 13428 10760
rect 13488 10700 13518 10760
rect 13578 10700 13588 10760
rect 13338 10690 13588 10700
rect 13618 10650 13658 10800
rect 13688 10760 13768 10770
rect 13688 10700 13698 10760
rect 13758 10700 13768 10760
rect 13688 10690 13768 10700
rect 13868 10760 13948 10770
rect 13868 10700 13878 10760
rect 13938 10700 13948 10760
rect 13868 10690 13948 10700
rect 13978 10650 14018 10910
rect 14048 10760 14128 10770
rect 14048 10700 14058 10760
rect 14118 10700 14128 10760
rect 14048 10690 14128 10700
rect 14228 10760 14308 10770
rect 14228 10700 14238 10760
rect 14298 10700 14308 10760
rect 14228 10690 14308 10700
rect 14338 10650 14378 11020
rect 14408 10760 14488 10770
rect 14408 10700 14418 10760
rect 14478 10700 14488 10760
rect 14408 10690 14488 10700
rect 14588 10760 14658 10770
rect 14588 10700 14598 10760
rect 14588 10690 14658 10700
rect 13248 10590 13258 10630
rect 13298 10590 13308 10630
rect 13248 10530 13308 10590
rect 13248 10490 13258 10530
rect 13298 10490 13308 10530
rect 13248 10430 13308 10490
rect 13248 10390 13258 10430
rect 13298 10390 13308 10430
rect 13248 10330 13308 10390
rect 13248 10290 13258 10330
rect 13298 10290 13308 10330
rect 13248 10230 13308 10290
rect 13248 10190 13258 10230
rect 13298 10190 13308 10230
rect 13248 10130 13308 10190
rect 13248 10090 13258 10130
rect 13298 10090 13308 10130
rect 13248 10070 13308 10090
rect 13428 10630 13488 10650
rect 13428 10590 13438 10630
rect 13478 10590 13488 10630
rect 13428 10530 13488 10590
rect 13428 10490 13438 10530
rect 13478 10490 13488 10530
rect 13428 10430 13488 10490
rect 13428 10390 13438 10430
rect 13478 10390 13488 10430
rect 13428 10330 13488 10390
rect 13428 10290 13438 10330
rect 13478 10290 13488 10330
rect 13428 10230 13488 10290
rect 13428 10190 13438 10230
rect 13478 10190 13488 10230
rect 13428 10130 13488 10190
rect 13428 10090 13438 10130
rect 13478 10090 13488 10130
rect 13428 10070 13488 10090
rect 13608 10630 13668 10650
rect 13608 10590 13618 10630
rect 13658 10590 13668 10630
rect 13608 10530 13668 10590
rect 13608 10490 13618 10530
rect 13658 10490 13668 10530
rect 13608 10430 13668 10490
rect 13608 10390 13618 10430
rect 13658 10390 13668 10430
rect 13608 10330 13668 10390
rect 13608 10290 13618 10330
rect 13658 10290 13668 10330
rect 13608 10230 13668 10290
rect 13608 10190 13618 10230
rect 13658 10190 13668 10230
rect 13608 10130 13668 10190
rect 13608 10090 13618 10130
rect 13658 10090 13668 10130
rect 13608 10070 13668 10090
rect 13788 10630 13848 10650
rect 13788 10590 13798 10630
rect 13838 10590 13848 10630
rect 13788 10530 13848 10590
rect 13788 10490 13798 10530
rect 13838 10490 13848 10530
rect 13788 10430 13848 10490
rect 13788 10390 13798 10430
rect 13838 10390 13848 10430
rect 13788 10330 13848 10390
rect 13788 10290 13798 10330
rect 13838 10290 13848 10330
rect 13788 10230 13848 10290
rect 13788 10190 13798 10230
rect 13838 10190 13848 10230
rect 13788 10130 13848 10190
rect 13788 10090 13798 10130
rect 13838 10090 13848 10130
rect 13788 10070 13848 10090
rect 13968 10630 14028 10650
rect 13968 10590 13978 10630
rect 14018 10590 14028 10630
rect 13968 10530 14028 10590
rect 13968 10490 13978 10530
rect 14018 10490 14028 10530
rect 13968 10430 14028 10490
rect 13968 10390 13978 10430
rect 14018 10390 14028 10430
rect 13968 10330 14028 10390
rect 13968 10290 13978 10330
rect 14018 10290 14028 10330
rect 13968 10230 14028 10290
rect 13968 10190 13978 10230
rect 14018 10190 14028 10230
rect 13968 10130 14028 10190
rect 13968 10090 13978 10130
rect 14018 10090 14028 10130
rect 13968 10070 14028 10090
rect 14148 10630 14208 10650
rect 14148 10590 14158 10630
rect 14198 10590 14208 10630
rect 14148 10530 14208 10590
rect 14148 10490 14158 10530
rect 14198 10490 14208 10530
rect 14148 10430 14208 10490
rect 14148 10390 14158 10430
rect 14198 10390 14208 10430
rect 14148 10330 14208 10390
rect 14148 10290 14158 10330
rect 14198 10290 14208 10330
rect 14148 10230 14208 10290
rect 14148 10190 14158 10230
rect 14198 10190 14208 10230
rect 14148 10130 14208 10190
rect 14148 10090 14158 10130
rect 14198 10090 14208 10130
rect 14148 10070 14208 10090
rect 14328 10630 14388 10650
rect 14328 10590 14338 10630
rect 14378 10590 14388 10630
rect 14328 10530 14388 10590
rect 14328 10490 14338 10530
rect 14378 10490 14388 10530
rect 14328 10430 14388 10490
rect 14328 10390 14338 10430
rect 14378 10390 14388 10430
rect 14328 10330 14388 10390
rect 14328 10290 14338 10330
rect 14378 10290 14388 10330
rect 14328 10230 14388 10290
rect 14328 10190 14338 10230
rect 14378 10190 14388 10230
rect 14328 10130 14388 10190
rect 14328 10090 14338 10130
rect 14378 10090 14388 10130
rect 14328 10070 14388 10090
rect 14508 10630 14568 10650
rect 14508 10590 14518 10630
rect 14558 10590 14568 10630
rect 14508 10530 14568 10590
rect 14508 10490 14518 10530
rect 14558 10490 14568 10530
rect 14508 10430 14568 10490
rect 14508 10390 14518 10430
rect 14558 10390 14568 10430
rect 14508 10330 14568 10390
rect 14508 10290 14518 10330
rect 14558 10290 14568 10330
rect 14508 10230 14568 10290
rect 14508 10190 14518 10230
rect 14558 10190 14568 10230
rect 14508 10130 14568 10190
rect 14508 10090 14518 10130
rect 14558 10090 14568 10130
rect 14508 10070 14568 10090
rect 14688 10630 14748 11130
rect 15708 11090 15788 11100
rect 15708 11030 15718 11090
rect 15778 11030 15788 11090
rect 15238 10980 15318 10990
rect 15238 10920 15248 10980
rect 15308 10920 15318 10980
rect 15238 10910 15318 10920
rect 14688 10590 14698 10630
rect 14738 10590 14748 10630
rect 14688 10530 14748 10590
rect 14688 10490 14698 10530
rect 14738 10490 14748 10530
rect 14688 10430 14748 10490
rect 14688 10390 14698 10430
rect 14738 10390 14748 10430
rect 14688 10330 14748 10390
rect 14688 10290 14698 10330
rect 14738 10290 14748 10330
rect 14688 10230 14748 10290
rect 14688 10190 14698 10230
rect 14738 10190 14748 10230
rect 14688 10130 14748 10190
rect 14688 10090 14698 10130
rect 14738 10090 14748 10130
rect 14688 10070 14748 10090
rect 14868 10630 14928 10650
rect 14868 10590 14878 10630
rect 14918 10590 14928 10630
rect 14868 10530 14928 10590
rect 14868 10490 14878 10530
rect 14918 10490 14928 10530
rect 14868 10430 14928 10490
rect 14868 10390 14878 10430
rect 14918 10390 14928 10430
rect 14868 10330 14928 10390
rect 14868 10290 14878 10330
rect 14918 10290 14928 10330
rect 14868 10230 14928 10290
rect 15258 10230 15298 10910
rect 15588 10560 15668 10570
rect 15588 10500 15598 10560
rect 15658 10500 15668 10560
rect 15588 10490 15668 10500
rect 15708 10550 15788 11030
rect 15838 10570 15918 11520
rect 15968 11570 16028 11650
rect 15968 11530 15978 11570
rect 16018 11530 16028 11570
rect 15968 11480 16028 11530
rect 15958 11470 16038 11480
rect 15958 11410 15968 11470
rect 16028 11410 16038 11470
rect 15958 11390 16038 11410
rect 15958 11330 15968 11390
rect 16028 11330 16038 11390
rect 15958 11310 16038 11330
rect 15958 11250 15968 11310
rect 16028 11250 16038 11310
rect 15958 11240 16038 11250
rect 16168 10880 16208 12680
rect 16258 12530 16298 14730
rect 16238 12520 16318 12530
rect 16238 12460 16248 12520
rect 16308 12460 16318 12520
rect 16238 12450 16318 12460
rect 16258 10990 16298 12450
rect 16348 12200 16588 15290
rect 16778 14490 16858 17441
rect 16778 14430 16788 14490
rect 16848 14430 16858 14490
rect 16778 14420 16858 14430
rect 17568 17631 17648 17650
rect 17568 17234 17588 17631
rect 17626 17234 17648 17631
rect 17568 16750 17648 17234
rect 17568 16690 17578 16750
rect 17638 16690 17648 16750
rect 16348 12140 16358 12200
rect 16418 12140 16438 12200
rect 16498 12140 16518 12200
rect 16578 12140 16588 12200
rect 16348 12120 16588 12140
rect 16348 12060 16358 12120
rect 16418 12060 16438 12120
rect 16498 12060 16518 12120
rect 16578 12060 16588 12120
rect 16348 12040 16588 12060
rect 16348 11980 16358 12040
rect 16418 11980 16438 12040
rect 16498 11980 16518 12040
rect 16578 11980 16588 12040
rect 16348 11970 16588 11980
rect 17568 11580 17648 16690
rect 17948 16050 18028 18050
rect 17948 15990 17958 16050
rect 18018 15990 18028 16050
rect 17948 15980 18028 15990
rect 18118 17450 18198 17460
rect 18118 17390 18128 17450
rect 18188 17390 18198 17450
rect 18118 13440 18198 17390
rect 18648 14380 18728 18070
rect 18778 16750 18878 16770
rect 18778 16690 18798 16750
rect 18858 16690 18878 16750
rect 18778 16670 18878 16690
rect 18778 15350 18878 15370
rect 18778 15290 18798 15350
rect 18858 15290 18878 15350
rect 18778 15270 18878 15290
rect 18648 14320 18658 14380
rect 18718 14320 18728 14380
rect 18648 14310 18728 14320
rect 23208 13510 23308 13530
rect 23208 13450 23228 13510
rect 23288 13450 23308 13510
rect 18038 13420 18278 13440
rect 23208 13430 23308 13450
rect 18038 13360 18078 13420
rect 18138 13360 18178 13420
rect 18238 13360 18278 13420
rect 18038 13340 18278 13360
rect 23008 13180 23088 13190
rect 23008 13120 23018 13180
rect 23078 13120 23088 13180
rect 23008 13110 23088 13120
rect 23218 13130 23298 13430
rect 17568 11520 17578 11580
rect 17638 11520 17648 11580
rect 17568 11510 17648 11520
rect 19138 12790 19218 12800
rect 19138 12730 19148 12790
rect 19208 12730 19218 12790
rect 19028 11410 19108 11420
rect 19028 11350 19038 11410
rect 19098 11350 19108 11410
rect 18918 11250 18998 11260
rect 18918 11190 18928 11250
rect 18988 11190 18998 11250
rect 16238 10980 16318 10990
rect 16238 10920 16248 10980
rect 16308 10920 16318 10980
rect 16238 10910 16318 10920
rect 16148 10870 16228 10880
rect 16148 10810 16158 10870
rect 16218 10810 16228 10870
rect 16148 10800 16228 10810
rect 15708 10510 15728 10550
rect 15768 10510 15788 10550
rect 15708 10490 15788 10510
rect 15828 10560 15908 10570
rect 15828 10500 15838 10560
rect 15898 10500 15908 10560
rect 15828 10490 15908 10500
rect 15498 10430 15558 10450
rect 15498 10390 15508 10430
rect 15548 10390 15558 10430
rect 15498 10330 15558 10390
rect 15498 10290 15508 10330
rect 15548 10290 15558 10330
rect 15498 10230 15558 10290
rect 15608 10430 15668 10490
rect 15608 10390 15618 10430
rect 15658 10390 15668 10430
rect 15608 10330 15668 10390
rect 15608 10290 15618 10330
rect 15658 10290 15668 10330
rect 15608 10270 15668 10290
rect 15718 10430 15778 10450
rect 15718 10390 15728 10430
rect 15768 10390 15778 10430
rect 15718 10330 15778 10390
rect 15718 10290 15728 10330
rect 15768 10290 15778 10330
rect 15718 10230 15778 10290
rect 15828 10430 15888 10490
rect 15828 10390 15838 10430
rect 15878 10390 15888 10430
rect 15828 10330 15888 10390
rect 15828 10290 15838 10330
rect 15878 10290 15888 10330
rect 15828 10270 15888 10290
rect 15938 10430 15998 10450
rect 15938 10390 15948 10430
rect 15988 10390 15998 10430
rect 15938 10330 15998 10390
rect 15938 10290 15948 10330
rect 15988 10290 15998 10330
rect 15938 10230 15998 10290
rect 14868 10190 14878 10230
rect 14918 10190 14928 10230
rect 14868 10130 14928 10190
rect 15238 10220 15318 10230
rect 15238 10160 15248 10220
rect 15308 10160 15318 10220
rect 15238 10150 15318 10160
rect 15488 10210 15568 10230
rect 15488 10170 15508 10210
rect 15548 10170 15568 10210
rect 15488 10150 15568 10170
rect 15708 10220 15788 10230
rect 15708 10160 15718 10220
rect 15778 10160 15788 10220
rect 15708 10150 15788 10160
rect 15928 10210 16008 10230
rect 15928 10170 15948 10210
rect 15988 10170 16008 10210
rect 15928 10150 16008 10170
rect 14868 10090 14878 10130
rect 14918 10090 14928 10130
rect 14868 10070 14928 10090
rect 15498 10030 15558 10150
rect 15938 10030 15998 10150
rect 11618 10020 11698 10030
rect 11618 9960 11628 10020
rect 11688 9960 11698 10020
rect 11618 9940 11698 9960
rect 11618 9880 11628 9940
rect 11688 9880 11698 9940
rect 11618 9860 11698 9880
rect 11618 9800 11628 9860
rect 11688 9800 11698 9860
rect 11618 9790 11698 9800
rect 11978 10020 12058 10030
rect 11978 9960 11988 10020
rect 12048 9960 12058 10020
rect 11978 9940 12058 9960
rect 11978 9880 11988 9940
rect 12048 9880 12058 9940
rect 11978 9860 12058 9880
rect 11978 9800 11988 9860
rect 12048 9800 12058 9860
rect 11978 9790 12058 9800
rect 12338 10020 12418 10030
rect 12338 9960 12348 10020
rect 12408 9960 12418 10020
rect 12338 9940 12418 9960
rect 12338 9880 12348 9940
rect 12408 9880 12418 9940
rect 12338 9860 12418 9880
rect 12338 9800 12348 9860
rect 12408 9800 12418 9860
rect 12338 9790 12418 9800
rect 12698 10020 12778 10030
rect 12698 9960 12708 10020
rect 12768 9960 12778 10020
rect 12698 9940 12778 9960
rect 12698 9880 12708 9940
rect 12768 9880 12778 9940
rect 12698 9860 12778 9880
rect 12698 9800 12708 9860
rect 12768 9800 12778 9860
rect 12698 9790 12778 9800
rect 13058 10020 13138 10030
rect 13058 9960 13068 10020
rect 13128 9960 13138 10020
rect 13058 9940 13138 9960
rect 13058 9880 13068 9940
rect 13128 9880 13138 9940
rect 13058 9860 13138 9880
rect 13058 9800 13068 9860
rect 13128 9800 13138 9860
rect 13058 9790 13138 9800
rect 13418 10020 13498 10030
rect 13418 9960 13428 10020
rect 13488 9960 13498 10020
rect 13418 9940 13498 9960
rect 13418 9880 13428 9940
rect 13488 9880 13498 9940
rect 13418 9860 13498 9880
rect 13418 9800 13428 9860
rect 13488 9800 13498 9860
rect 13418 9790 13498 9800
rect 13778 10020 13858 10030
rect 13778 9960 13788 10020
rect 13848 9960 13858 10020
rect 13778 9940 13858 9960
rect 13778 9880 13788 9940
rect 13848 9880 13858 9940
rect 13778 9860 13858 9880
rect 13778 9800 13788 9860
rect 13848 9800 13858 9860
rect 13778 9790 13858 9800
rect 14138 10020 14218 10030
rect 14138 9960 14148 10020
rect 14208 9960 14218 10020
rect 14138 9940 14218 9960
rect 14138 9880 14148 9940
rect 14208 9880 14218 9940
rect 14138 9860 14218 9880
rect 14138 9800 14148 9860
rect 14208 9800 14218 9860
rect 14138 9790 14218 9800
rect 14498 10020 14578 10030
rect 14498 9960 14508 10020
rect 14568 9960 14578 10020
rect 14498 9940 14578 9960
rect 14498 9880 14508 9940
rect 14568 9880 14578 9940
rect 14498 9860 14578 9880
rect 14498 9800 14508 9860
rect 14568 9800 14578 9860
rect 14498 9790 14578 9800
rect 14858 10020 14938 10030
rect 14858 9960 14868 10020
rect 14928 9960 14938 10020
rect 14858 9940 14938 9960
rect 14858 9880 14868 9940
rect 14928 9880 14938 9940
rect 14858 9860 14938 9880
rect 14858 9800 14868 9860
rect 14928 9800 14938 9860
rect 14858 9790 14938 9800
rect 15488 10020 15568 10030
rect 15488 9960 15498 10020
rect 15558 9960 15568 10020
rect 15488 9940 15568 9960
rect 15488 9880 15498 9940
rect 15558 9880 15568 9940
rect 15488 9860 15568 9880
rect 15488 9800 15498 9860
rect 15558 9800 15568 9860
rect 15488 9790 15568 9800
rect 15928 10020 16008 10030
rect 15928 9960 15938 10020
rect 15998 9960 16008 10020
rect 15928 9940 16008 9960
rect 15928 9880 15938 9940
rect 15998 9880 16008 9940
rect 15928 9860 16008 9880
rect 15928 9800 15938 9860
rect 15998 9800 16008 9860
rect 15928 9790 16008 9800
rect 11804 9750 11862 9760
rect 11804 9698 11806 9750
rect 11858 9698 11862 9750
rect 11804 9690 11862 9698
rect 11914 9750 11972 9760
rect 11914 9698 11916 9750
rect 11968 9698 11972 9750
rect 11914 9690 11972 9698
rect 12024 9750 12082 9760
rect 12024 9698 12026 9750
rect 12078 9698 12082 9750
rect 12024 9690 12082 9698
rect 12134 9750 12192 9760
rect 12134 9698 12136 9750
rect 12188 9698 12192 9750
rect 12134 9690 12192 9698
rect 12244 9750 12302 9760
rect 12244 9698 12246 9750
rect 12298 9698 12302 9750
rect 12244 9690 12302 9698
rect 12354 9750 12412 9760
rect 12354 9698 12356 9750
rect 12408 9698 12412 9750
rect 12354 9690 12412 9698
rect 12464 9750 12522 9760
rect 12464 9698 12466 9750
rect 12518 9698 12522 9750
rect 12464 9690 12522 9698
rect 12574 9750 12632 9760
rect 12574 9698 12576 9750
rect 12628 9698 12632 9750
rect 12574 9690 12632 9698
rect 12684 9750 12742 9760
rect 12684 9698 12686 9750
rect 12738 9698 12742 9750
rect 12684 9690 12742 9698
rect 12794 9750 12852 9760
rect 12794 9698 12796 9750
rect 12848 9698 12852 9750
rect 12794 9690 12852 9698
rect 13704 9750 13762 9760
rect 13704 9698 13706 9750
rect 13758 9698 13762 9750
rect 13704 9690 13762 9698
rect 13814 9750 13872 9760
rect 13814 9698 13816 9750
rect 13868 9698 13872 9750
rect 13814 9690 13872 9698
rect 13924 9750 13982 9760
rect 13924 9698 13926 9750
rect 13978 9698 13982 9750
rect 13924 9690 13982 9698
rect 14034 9750 14092 9760
rect 14034 9698 14036 9750
rect 14088 9698 14092 9750
rect 14034 9690 14092 9698
rect 14144 9750 14202 9760
rect 14144 9698 14146 9750
rect 14198 9698 14202 9750
rect 14144 9690 14202 9698
rect 14254 9750 14312 9760
rect 14254 9698 14256 9750
rect 14308 9698 14312 9750
rect 14254 9690 14312 9698
rect 14364 9750 14422 9760
rect 14364 9698 14366 9750
rect 14418 9698 14422 9750
rect 14364 9690 14422 9698
rect 14474 9750 14532 9760
rect 14474 9698 14476 9750
rect 14528 9698 14532 9750
rect 14474 9690 14532 9698
rect 14584 9750 14642 9760
rect 14584 9698 14586 9750
rect 14638 9698 14642 9750
rect 14584 9690 14642 9698
rect 14694 9750 14752 9760
rect 14694 9698 14696 9750
rect 14748 9698 14752 9750
rect 14694 9690 14752 9698
rect 11558 9630 11698 9650
rect 11558 9590 11568 9630
rect 11608 9590 11648 9630
rect 11688 9590 11698 9630
rect 11558 9530 11698 9590
rect 11558 9490 11568 9530
rect 11608 9490 11648 9530
rect 11688 9490 11698 9530
rect 11558 9470 11698 9490
rect 11638 9430 11698 9470
rect 11748 9630 11808 9650
rect 11748 9590 11758 9630
rect 11798 9590 11808 9630
rect 11748 9530 11808 9590
rect 11748 9490 11758 9530
rect 11798 9490 11808 9530
rect 11628 9420 11708 9430
rect 11628 9360 11638 9420
rect 11698 9360 11708 9420
rect 11628 9350 11708 9360
rect 11748 9320 11808 9490
rect 11858 9630 11918 9650
rect 11858 9590 11868 9630
rect 11908 9590 11918 9630
rect 11858 9530 11918 9590
rect 11858 9490 11868 9530
rect 11908 9490 11918 9530
rect 11858 9430 11918 9490
rect 11968 9630 12028 9650
rect 11968 9590 11978 9630
rect 12018 9590 12028 9630
rect 11968 9530 12028 9590
rect 11968 9490 11978 9530
rect 12018 9490 12028 9530
rect 11848 9420 11928 9430
rect 11848 9360 11858 9420
rect 11918 9360 11928 9420
rect 11848 9350 11928 9360
rect 11968 9320 12028 9490
rect 12078 9630 12138 9650
rect 12078 9590 12088 9630
rect 12128 9590 12138 9630
rect 12078 9530 12138 9590
rect 12078 9490 12088 9530
rect 12128 9490 12138 9530
rect 12078 9430 12138 9490
rect 12188 9630 12248 9650
rect 12188 9590 12198 9630
rect 12238 9590 12248 9630
rect 12188 9530 12248 9590
rect 12188 9490 12198 9530
rect 12238 9490 12248 9530
rect 12068 9420 12148 9430
rect 12068 9360 12078 9420
rect 12138 9360 12148 9420
rect 12068 9350 12148 9360
rect 12188 9320 12248 9490
rect 12298 9630 12358 9650
rect 12298 9590 12308 9630
rect 12348 9590 12358 9630
rect 12298 9530 12358 9590
rect 12298 9490 12308 9530
rect 12348 9490 12358 9530
rect 12298 9430 12358 9490
rect 12408 9630 12468 9650
rect 12408 9590 12418 9630
rect 12458 9590 12468 9630
rect 12408 9530 12468 9590
rect 12408 9490 12418 9530
rect 12458 9490 12468 9530
rect 12288 9420 12368 9430
rect 12288 9360 12298 9420
rect 12358 9360 12368 9420
rect 12288 9350 12368 9360
rect 12408 9320 12468 9490
rect 12518 9630 12578 9650
rect 12518 9590 12528 9630
rect 12568 9590 12578 9630
rect 12518 9530 12578 9590
rect 12518 9490 12528 9530
rect 12568 9490 12578 9530
rect 12518 9430 12578 9490
rect 12628 9630 12688 9650
rect 12628 9590 12638 9630
rect 12678 9590 12688 9630
rect 12628 9530 12688 9590
rect 12628 9490 12638 9530
rect 12678 9490 12688 9530
rect 12508 9420 12588 9430
rect 12508 9360 12518 9420
rect 12578 9360 12588 9420
rect 12508 9350 12588 9360
rect 12628 9320 12688 9490
rect 12738 9630 12798 9650
rect 12738 9590 12748 9630
rect 12788 9590 12798 9630
rect 12738 9530 12798 9590
rect 12738 9490 12748 9530
rect 12788 9490 12798 9530
rect 12738 9430 12798 9490
rect 12848 9630 12908 9650
rect 12848 9590 12858 9630
rect 12898 9590 12908 9630
rect 12848 9530 12908 9590
rect 12848 9490 12858 9530
rect 12898 9490 12908 9530
rect 12728 9420 12808 9430
rect 12728 9360 12738 9420
rect 12798 9360 12808 9420
rect 12728 9350 12808 9360
rect 12848 9320 12908 9490
rect 12958 9630 13098 9650
rect 12958 9590 12968 9630
rect 13008 9590 13048 9630
rect 13088 9590 13098 9630
rect 12958 9530 13098 9590
rect 12958 9490 12968 9530
rect 13008 9490 13048 9530
rect 13088 9490 13098 9530
rect 12958 9470 13098 9490
rect 13458 9630 13598 9650
rect 13458 9590 13468 9630
rect 13508 9590 13548 9630
rect 13588 9590 13598 9630
rect 13458 9530 13598 9590
rect 13458 9490 13468 9530
rect 13508 9490 13548 9530
rect 13588 9490 13598 9530
rect 13458 9470 13598 9490
rect 12958 9430 13018 9470
rect 13538 9430 13598 9470
rect 13648 9630 13708 9650
rect 13648 9590 13658 9630
rect 13698 9590 13708 9630
rect 13648 9530 13708 9590
rect 13648 9490 13658 9530
rect 13698 9490 13708 9530
rect 12948 9420 13028 9430
rect 12948 9360 12958 9420
rect 13018 9360 13028 9420
rect 12948 9350 13028 9360
rect 13528 9420 13608 9430
rect 13528 9360 13538 9420
rect 13598 9360 13608 9420
rect 13528 9350 13608 9360
rect 9678 9250 9688 9310
rect 9748 9250 9758 9310
rect 9678 9240 9758 9250
rect 11738 9310 11818 9320
rect 11738 9250 11748 9310
rect 11808 9250 11818 9310
rect 11738 9240 11818 9250
rect 11958 9310 12038 9320
rect 11958 9250 11968 9310
rect 12028 9250 12038 9310
rect 11958 9240 12038 9250
rect 12178 9310 12258 9320
rect 12178 9250 12188 9310
rect 12248 9250 12258 9310
rect 12178 9240 12258 9250
rect 12398 9310 12478 9320
rect 12398 9250 12408 9310
rect 12468 9250 12478 9310
rect 12398 9240 12478 9250
rect 12618 9310 12698 9320
rect 12618 9250 12628 9310
rect 12688 9250 12698 9310
rect 12618 9240 12698 9250
rect 12838 9310 12918 9320
rect 13648 9310 13708 9490
rect 13758 9630 13818 9650
rect 13758 9590 13768 9630
rect 13808 9590 13818 9630
rect 13758 9530 13818 9590
rect 13758 9490 13768 9530
rect 13808 9490 13818 9530
rect 13758 9430 13818 9490
rect 13868 9630 13928 9650
rect 13868 9590 13878 9630
rect 13918 9590 13928 9630
rect 13868 9530 13928 9590
rect 13868 9490 13878 9530
rect 13918 9490 13928 9530
rect 13748 9420 13828 9430
rect 13748 9360 13758 9420
rect 13818 9360 13828 9420
rect 13748 9350 13828 9360
rect 13868 9310 13928 9490
rect 13978 9630 14038 9650
rect 13978 9590 13988 9630
rect 14028 9590 14038 9630
rect 13978 9530 14038 9590
rect 13978 9490 13988 9530
rect 14028 9490 14038 9530
rect 13978 9430 14038 9490
rect 14088 9630 14148 9650
rect 14088 9590 14098 9630
rect 14138 9590 14148 9630
rect 14088 9530 14148 9590
rect 14088 9490 14098 9530
rect 14138 9490 14148 9530
rect 13968 9420 14048 9430
rect 13968 9360 13978 9420
rect 14038 9360 14048 9420
rect 13968 9350 14048 9360
rect 14088 9310 14148 9490
rect 14198 9630 14258 9650
rect 14198 9590 14208 9630
rect 14248 9590 14258 9630
rect 14198 9530 14258 9590
rect 14198 9490 14208 9530
rect 14248 9490 14258 9530
rect 14198 9430 14258 9490
rect 14308 9630 14368 9650
rect 14308 9590 14318 9630
rect 14358 9590 14368 9630
rect 14308 9530 14368 9590
rect 14308 9490 14318 9530
rect 14358 9490 14368 9530
rect 14188 9420 14268 9430
rect 14188 9360 14198 9420
rect 14258 9360 14268 9420
rect 14188 9350 14268 9360
rect 14308 9310 14368 9490
rect 14418 9630 14478 9650
rect 14418 9590 14428 9630
rect 14468 9590 14478 9630
rect 14418 9530 14478 9590
rect 14418 9490 14428 9530
rect 14468 9490 14478 9530
rect 14418 9430 14478 9490
rect 14528 9630 14588 9650
rect 14528 9590 14538 9630
rect 14578 9590 14588 9630
rect 14528 9530 14588 9590
rect 14528 9490 14538 9530
rect 14578 9490 14588 9530
rect 14408 9420 14488 9430
rect 14408 9360 14418 9420
rect 14478 9360 14488 9420
rect 14408 9350 14488 9360
rect 14528 9310 14588 9490
rect 14638 9630 14698 9650
rect 14638 9590 14648 9630
rect 14688 9590 14698 9630
rect 14638 9530 14698 9590
rect 14638 9490 14648 9530
rect 14688 9490 14698 9530
rect 14638 9430 14698 9490
rect 14748 9630 14808 9650
rect 14748 9590 14758 9630
rect 14798 9590 14808 9630
rect 14748 9530 14808 9590
rect 14748 9490 14758 9530
rect 14798 9490 14808 9530
rect 14628 9420 14708 9430
rect 14628 9360 14638 9420
rect 14698 9360 14708 9420
rect 14628 9350 14708 9360
rect 14748 9310 14808 9490
rect 14858 9630 14998 9650
rect 14858 9590 14868 9630
rect 14908 9590 14948 9630
rect 14988 9590 14998 9630
rect 14858 9530 14998 9590
rect 14858 9490 14868 9530
rect 14908 9490 14948 9530
rect 14988 9490 14998 9530
rect 14858 9470 14998 9490
rect 14858 9430 14918 9470
rect 14848 9420 14928 9430
rect 14848 9360 14858 9420
rect 14918 9360 14928 9420
rect 14848 9350 14928 9360
rect 12838 9250 12848 9310
rect 12908 9250 12918 9310
rect 12838 9240 12918 9250
rect 13638 9300 13718 9310
rect 13638 9240 13648 9300
rect 13708 9240 13718 9300
rect 13638 9220 13718 9240
rect 13638 9160 13648 9220
rect 13708 9160 13718 9220
rect 13638 9140 13718 9160
rect 13638 9080 13648 9140
rect 13708 9080 13718 9140
rect 13638 9070 13718 9080
rect 13858 9300 13938 9310
rect 13858 9240 13868 9300
rect 13928 9240 13938 9300
rect 13858 9220 13938 9240
rect 13858 9160 13868 9220
rect 13928 9160 13938 9220
rect 13858 9140 13938 9160
rect 13858 9080 13868 9140
rect 13928 9080 13938 9140
rect 13858 9070 13938 9080
rect 14078 9300 14158 9310
rect 14078 9240 14088 9300
rect 14148 9240 14158 9300
rect 14078 9220 14158 9240
rect 14078 9160 14088 9220
rect 14148 9160 14158 9220
rect 14078 9140 14158 9160
rect 14078 9080 14088 9140
rect 14148 9080 14158 9140
rect 14078 9070 14158 9080
rect 14298 9300 14378 9310
rect 14298 9240 14308 9300
rect 14368 9240 14378 9300
rect 14298 9220 14378 9240
rect 14298 9160 14308 9220
rect 14368 9160 14378 9220
rect 14298 9140 14378 9160
rect 14298 9080 14308 9140
rect 14368 9080 14378 9140
rect 14298 9070 14378 9080
rect 14518 9300 14598 9310
rect 14518 9240 14528 9300
rect 14588 9240 14598 9300
rect 14518 9220 14598 9240
rect 14518 9160 14528 9220
rect 14588 9160 14598 9220
rect 14518 9140 14598 9160
rect 14518 9080 14528 9140
rect 14588 9080 14598 9140
rect 14518 9070 14598 9080
rect 14738 9300 14818 9310
rect 14738 9240 14748 9300
rect 14808 9240 14818 9300
rect 14738 9220 14818 9240
rect 14738 9160 14748 9220
rect 14808 9160 14818 9220
rect 14738 9140 14818 9160
rect 14738 9080 14748 9140
rect 14808 9080 14818 9140
rect 14738 9070 14818 9080
rect 18648 9300 18888 9310
rect 18648 9240 18658 9300
rect 18718 9240 18738 9300
rect 18798 9240 18818 9300
rect 18878 9240 18888 9300
rect 18648 9220 18888 9240
rect 18648 9160 18658 9220
rect 18718 9160 18738 9220
rect 18798 9160 18818 9220
rect 18878 9160 18888 9220
rect 18648 9140 18888 9160
rect 18648 9080 18658 9140
rect 18718 9080 18738 9140
rect 18798 9080 18818 9140
rect 18878 9080 18888 9140
rect 18098 8370 18178 8380
rect 18098 8310 18108 8370
rect 18168 8310 18178 8370
rect 13248 8300 13328 8310
rect 13248 8240 13258 8300
rect 13318 8240 13328 8300
rect 13248 8230 13328 8240
rect 13468 8300 13548 8310
rect 13468 8240 13478 8300
rect 13538 8240 13548 8300
rect 13468 8230 13548 8240
rect 13768 8300 13848 8310
rect 13768 8240 13778 8300
rect 13838 8240 13848 8300
rect 13768 8230 13848 8240
rect 13998 8300 14078 8310
rect 13998 8240 14008 8300
rect 14068 8240 14078 8300
rect 13998 8230 14078 8240
rect 14148 8300 14228 8310
rect 14148 8240 14158 8300
rect 14218 8240 14228 8300
rect 14148 8230 14228 8240
rect 14368 8300 14448 8310
rect 14368 8240 14378 8300
rect 14438 8240 14448 8300
rect 14368 8230 14448 8240
rect 14668 8300 14748 8310
rect 14668 8240 14678 8300
rect 14738 8240 14748 8300
rect 14668 8230 14748 8240
rect 14888 8300 14968 8310
rect 14888 8240 14898 8300
rect 14958 8240 14968 8300
rect 14888 8230 14968 8240
rect 15288 8300 15368 8310
rect 15288 8240 15298 8300
rect 15358 8240 15368 8300
rect 15288 8230 15368 8240
rect 15618 8300 15698 8310
rect 15618 8240 15628 8300
rect 15688 8240 15698 8300
rect 15618 8230 15698 8240
rect 15948 8300 16028 8310
rect 15948 8240 15958 8300
rect 16018 8240 16028 8300
rect 15948 8230 16028 8240
rect 16388 8300 16468 8310
rect 16388 8240 16398 8300
rect 16458 8240 16468 8300
rect 16388 8230 16468 8240
rect 16648 8300 16728 8310
rect 16648 8240 16658 8300
rect 16718 8240 16728 8300
rect 16648 8230 16728 8240
rect 17168 8300 17248 8310
rect 17168 8240 17178 8300
rect 17238 8240 17248 8300
rect 17168 8230 17248 8240
rect 17848 8300 17928 8310
rect 17848 8240 17858 8300
rect 17918 8240 17928 8300
rect 17848 8230 17928 8240
rect 12108 7810 12188 7820
rect 12108 7750 12118 7810
rect 12178 7750 12188 7810
rect 11938 6430 12018 6440
rect 11938 6370 11948 6430
rect 12008 6370 12018 6430
rect 11938 1330 12018 6370
rect 12108 3340 12188 7750
rect 13128 7810 13208 7820
rect 13128 7750 13138 7810
rect 13198 7750 13208 7810
rect 13128 7740 13208 7750
rect 15048 7800 15128 7810
rect 15048 7740 15058 7800
rect 15118 7740 15128 7800
rect 15048 7730 15128 7740
rect 16078 7800 16198 7810
rect 16078 7740 16088 7800
rect 16148 7740 16198 7800
rect 16078 7730 16198 7740
rect 13698 7230 13778 7240
rect 13698 7170 13708 7230
rect 13768 7170 13778 7230
rect 13698 7160 13778 7170
rect 13248 7120 13328 7130
rect 13248 7060 13258 7120
rect 13318 7060 13328 7120
rect 13248 7050 13328 7060
rect 13988 7120 14068 7130
rect 13988 7060 13998 7120
rect 14058 7060 14068 7120
rect 13988 7050 14068 7060
rect 14148 7120 14228 7130
rect 14148 7060 14158 7120
rect 14218 7060 14228 7120
rect 14148 7050 14228 7060
rect 14888 7120 14968 7130
rect 14888 7060 14898 7120
rect 14958 7060 14968 7120
rect 14888 7050 14968 7060
rect 13128 6430 13208 6440
rect 13128 6370 13138 6430
rect 13198 6370 13208 6430
rect 15068 6410 15108 7730
rect 15228 7230 15308 7240
rect 15228 7170 15238 7230
rect 15298 7170 15308 7230
rect 15228 7160 15308 7170
rect 15138 7120 15218 7130
rect 15138 7060 15148 7120
rect 15208 7060 15218 7120
rect 15138 7050 15218 7060
rect 15248 7010 15288 7160
rect 15328 7120 15488 7130
rect 15328 7060 15338 7120
rect 15398 7060 15418 7120
rect 15478 7060 15488 7120
rect 15328 7050 15488 7060
rect 15618 7120 15698 7130
rect 15618 7060 15628 7120
rect 15688 7060 15698 7120
rect 15618 7050 15698 7060
rect 15948 7120 16028 7130
rect 15948 7060 15958 7120
rect 16018 7060 16028 7120
rect 15948 7050 16028 7060
rect 15248 6950 15258 7010
rect 15318 6950 15328 7010
rect 15248 6940 15328 6950
rect 16158 6450 16198 7730
rect 16228 7800 16308 7820
rect 16228 7760 16248 7800
rect 16288 7760 16308 7800
rect 16228 7740 16308 7760
rect 16228 7250 16268 7740
rect 16228 7240 16308 7250
rect 16228 7180 16238 7240
rect 16298 7180 16308 7240
rect 16668 7230 16708 8230
rect 16898 8190 17048 8200
rect 16898 8130 16908 8190
rect 16968 8130 17048 8190
rect 16898 8120 17048 8130
rect 17528 8190 17608 8200
rect 17528 8130 17538 8190
rect 17598 8130 17608 8190
rect 17528 8120 17608 8130
rect 18098 8190 18178 8310
rect 18098 8130 18108 8190
rect 18168 8130 18178 8190
rect 18098 8120 18178 8130
rect 16818 7230 16898 7240
rect 16228 7170 16308 7180
rect 16648 7170 16658 7230
rect 16718 7170 16728 7230
rect 16818 7170 16828 7230
rect 16888 7170 16898 7230
rect 17008 7130 17048 8120
rect 17998 7850 18078 7860
rect 17998 7790 18008 7850
rect 18068 7790 18078 7850
rect 17998 7780 18078 7790
rect 18178 7850 18258 7860
rect 18178 7790 18188 7850
rect 18248 7790 18258 7850
rect 18178 7490 18258 7790
rect 18178 7430 18188 7490
rect 18248 7430 18258 7490
rect 18178 7420 18258 7430
rect 18178 7380 18258 7390
rect 18178 7320 18188 7380
rect 18248 7320 18258 7380
rect 17458 7230 17538 7240
rect 17458 7170 17468 7230
rect 17528 7170 17538 7230
rect 17458 7160 17538 7170
rect 18178 7230 18258 7320
rect 18648 7380 18888 9080
rect 18648 7320 18658 7380
rect 18718 7320 18738 7380
rect 18798 7320 18818 7380
rect 18878 7320 18888 7380
rect 18648 7310 18888 7320
rect 18178 7170 18188 7230
rect 18248 7170 18258 7230
rect 18178 7160 18258 7170
rect 18288 7270 18368 7280
rect 18288 7210 18298 7270
rect 18358 7210 18368 7270
rect 16388 7120 16468 7130
rect 16388 7060 16398 7120
rect 16458 7060 16468 7120
rect 16388 7050 16468 7060
rect 16778 7120 16858 7130
rect 16778 7060 16788 7120
rect 16848 7060 16858 7120
rect 16778 7050 16858 7060
rect 16988 7120 17068 7130
rect 16988 7060 16998 7120
rect 17058 7060 17068 7120
rect 16988 7050 17068 7060
rect 17168 7120 17248 7130
rect 17168 7060 17178 7120
rect 17238 7060 17248 7120
rect 17168 7050 17248 7060
rect 17848 7120 17928 7130
rect 17848 7060 17858 7120
rect 17918 7060 17928 7120
rect 17848 7050 17928 7060
rect 13128 6360 13208 6370
rect 15028 6400 15108 6410
rect 15028 6340 15038 6400
rect 15098 6340 15108 6400
rect 16118 6440 16198 6450
rect 16118 6380 16128 6440
rect 16188 6380 16198 6440
rect 17688 6470 17768 6480
rect 16118 6370 16198 6380
rect 16248 6400 16328 6420
rect 15028 6330 15108 6340
rect 16248 6360 16268 6400
rect 16308 6360 16328 6400
rect 16248 6340 16328 6360
rect 17688 6410 17698 6470
rect 17758 6410 17768 6470
rect 16248 6080 16288 6340
rect 16228 6070 16308 6080
rect 13658 6050 13738 6060
rect 13658 5990 13668 6050
rect 13728 5990 13738 6050
rect 13658 5980 13738 5990
rect 15378 6050 15458 6060
rect 15378 5990 15388 6050
rect 15448 5990 15458 6050
rect 16228 6010 16238 6070
rect 16298 6010 16308 6070
rect 16228 6000 16308 6010
rect 17458 6050 17538 6060
rect 15378 5980 15458 5990
rect 17458 5990 17468 6050
rect 17528 5990 17538 6050
rect 17458 5980 17538 5990
rect 13248 5940 13328 5950
rect 13248 5880 13258 5940
rect 13318 5880 13328 5940
rect 13248 5870 13328 5880
rect 13468 5940 13548 5950
rect 13468 5880 13478 5940
rect 13538 5880 13548 5940
rect 13468 5870 13548 5880
rect 13768 5940 13848 5950
rect 13768 5880 13778 5940
rect 13838 5880 13848 5940
rect 13768 5870 13848 5880
rect 13988 5940 14068 5950
rect 13988 5880 13998 5940
rect 14058 5880 14068 5940
rect 13988 5870 14068 5880
rect 14148 5940 14228 5950
rect 14148 5880 14158 5940
rect 14218 5880 14228 5940
rect 14148 5870 14228 5880
rect 14368 5940 14448 5950
rect 14368 5880 14378 5940
rect 14438 5880 14448 5940
rect 14368 5870 14448 5880
rect 14668 5940 14748 5950
rect 14668 5880 14678 5940
rect 14738 5880 14748 5940
rect 14668 5870 14748 5880
rect 14888 5940 14968 5950
rect 14888 5880 14898 5940
rect 14958 5880 14968 5940
rect 14888 5870 14968 5880
rect 15188 5940 15268 5950
rect 15188 5880 15198 5940
rect 15258 5880 15268 5940
rect 15188 5870 15268 5880
rect 15628 5940 15708 5950
rect 15628 5880 15638 5940
rect 15698 5880 15708 5940
rect 15628 5870 15708 5880
rect 15958 5940 16038 5950
rect 15958 5880 15968 5940
rect 16028 5880 16038 5940
rect 15958 5870 16038 5880
rect 16388 5940 16468 5950
rect 16388 5880 16398 5940
rect 16458 5880 16468 5940
rect 16388 5870 16468 5880
rect 16778 5940 16858 5950
rect 16778 5880 16788 5940
rect 16848 5880 16858 5940
rect 16778 5870 16858 5880
rect 17168 5940 17248 5950
rect 17168 5880 17178 5940
rect 17238 5880 17248 5940
rect 17168 5870 17248 5880
rect 17688 5880 17768 6410
rect 17998 6390 18078 6400
rect 17998 6330 18008 6390
rect 18068 6330 18078 6390
rect 17998 6320 18078 6330
rect 18288 6390 18368 7210
rect 18288 6330 18298 6390
rect 18358 6330 18368 6390
rect 18288 6320 18368 6330
rect 18398 7160 18478 7170
rect 18398 7100 18408 7160
rect 18468 7100 18478 7160
rect 18398 6050 18478 7100
rect 18918 7040 18998 11190
rect 19028 8770 19108 11350
rect 19138 10030 19218 12730
rect 20318 12790 20398 12800
rect 20318 12730 20328 12790
rect 20388 12730 20398 12790
rect 19518 12660 19598 12680
rect 19518 12620 19538 12660
rect 19578 12620 19598 12660
rect 19518 12560 19598 12620
rect 19518 12520 19538 12560
rect 19578 12520 19598 12560
rect 19518 12460 19598 12520
rect 19518 12420 19538 12460
rect 19578 12420 19598 12460
rect 19518 12360 19598 12420
rect 19518 12320 19538 12360
rect 19578 12320 19598 12360
rect 19518 12260 19598 12320
rect 19518 12220 19538 12260
rect 19578 12220 19598 12260
rect 19518 12200 19598 12220
rect 19718 12660 19798 12680
rect 19718 12620 19738 12660
rect 19778 12620 19798 12660
rect 19718 12560 19798 12620
rect 19718 12520 19738 12560
rect 19778 12520 19798 12560
rect 19718 12460 19798 12520
rect 19718 12420 19738 12460
rect 19778 12420 19798 12460
rect 19718 12360 19798 12420
rect 19718 12320 19738 12360
rect 19778 12320 19798 12360
rect 19718 12260 19798 12320
rect 19718 12220 19738 12260
rect 19778 12220 19798 12260
rect 19518 12140 19598 12160
rect 19518 12100 19538 12140
rect 19578 12100 19598 12140
rect 19518 11990 19598 12100
rect 19518 11930 19528 11990
rect 19588 11930 19598 11990
rect 19518 11920 19598 11930
rect 19718 11990 19798 12220
rect 19718 11930 19728 11990
rect 19788 11930 19798 11990
rect 19718 11920 19798 11930
rect 19918 12660 19998 12680
rect 19918 12620 19938 12660
rect 19978 12620 19998 12660
rect 19918 12560 19998 12620
rect 19918 12520 19938 12560
rect 19978 12520 19998 12560
rect 19918 12460 19998 12520
rect 19918 12420 19938 12460
rect 19978 12420 19998 12460
rect 19918 12360 19998 12420
rect 19918 12320 19938 12360
rect 19978 12320 19998 12360
rect 19918 12260 19998 12320
rect 19918 12220 19938 12260
rect 19978 12220 19998 12260
rect 19918 12130 19998 12220
rect 19918 12070 19928 12130
rect 19988 12070 19998 12130
rect 19918 11880 19998 12070
rect 20118 12660 20198 12680
rect 20118 12620 20138 12660
rect 20178 12620 20198 12660
rect 20118 12560 20198 12620
rect 20118 12520 20138 12560
rect 20178 12520 20198 12560
rect 20118 12460 20198 12520
rect 20118 12420 20138 12460
rect 20178 12420 20198 12460
rect 20118 12360 20198 12420
rect 20118 12320 20138 12360
rect 20178 12320 20198 12360
rect 20118 12260 20198 12320
rect 20118 12220 20138 12260
rect 20178 12220 20198 12260
rect 20118 11990 20198 12220
rect 20318 12660 20398 12730
rect 20718 12790 20798 12800
rect 20718 12730 20728 12790
rect 20788 12730 20798 12790
rect 20318 12620 20338 12660
rect 20378 12620 20398 12660
rect 20318 12560 20398 12620
rect 20318 12520 20338 12560
rect 20378 12520 20398 12560
rect 20318 12460 20398 12520
rect 20318 12420 20338 12460
rect 20378 12420 20398 12460
rect 20318 12360 20398 12420
rect 20318 12320 20338 12360
rect 20378 12320 20398 12360
rect 20318 12260 20398 12320
rect 20318 12220 20338 12260
rect 20378 12220 20398 12260
rect 20318 12200 20398 12220
rect 20518 12660 20598 12680
rect 20518 12620 20538 12660
rect 20578 12620 20598 12660
rect 20518 12560 20598 12620
rect 20518 12520 20538 12560
rect 20578 12520 20598 12560
rect 20518 12460 20598 12520
rect 20518 12420 20538 12460
rect 20578 12420 20598 12460
rect 20518 12360 20598 12420
rect 20518 12320 20538 12360
rect 20578 12320 20598 12360
rect 20518 12260 20598 12320
rect 20518 12220 20538 12260
rect 20578 12220 20598 12260
rect 20118 11930 20128 11990
rect 20188 11930 20198 11990
rect 20118 11920 20198 11930
rect 20518 11990 20598 12220
rect 20718 12660 20798 12730
rect 23218 12733 23238 13130
rect 23276 12733 23298 13130
rect 23218 12720 23298 12733
rect 20718 12620 20738 12660
rect 20778 12620 20798 12660
rect 20718 12560 20798 12620
rect 20718 12520 20738 12560
rect 20778 12520 20798 12560
rect 20718 12460 20798 12520
rect 20718 12420 20738 12460
rect 20778 12420 20798 12460
rect 20718 12360 20798 12420
rect 20718 12320 20738 12360
rect 20778 12320 20798 12360
rect 20718 12260 20798 12320
rect 20718 12220 20738 12260
rect 20778 12220 20798 12260
rect 20718 12200 20798 12220
rect 20918 12660 20998 12680
rect 20918 12620 20938 12660
rect 20978 12620 20998 12660
rect 20918 12560 20998 12620
rect 20918 12520 20938 12560
rect 20978 12520 20998 12560
rect 20918 12460 20998 12520
rect 20918 12420 20938 12460
rect 20978 12420 20998 12460
rect 20918 12360 20998 12420
rect 20918 12320 20938 12360
rect 20978 12320 20998 12360
rect 20918 12260 20998 12320
rect 20918 12220 20938 12260
rect 20978 12220 20998 12260
rect 20518 11930 20528 11990
rect 20588 11930 20598 11990
rect 20518 11920 20598 11930
rect 20918 12000 20998 12220
rect 21118 12660 21198 12680
rect 21118 12620 21138 12660
rect 21178 12620 21198 12660
rect 21118 12560 21198 12620
rect 21118 12520 21138 12560
rect 21178 12520 21198 12560
rect 21118 12460 21198 12520
rect 21118 12420 21138 12460
rect 21178 12420 21198 12460
rect 21118 12360 21198 12420
rect 21118 12320 21138 12360
rect 21178 12320 21198 12360
rect 21118 12260 21198 12320
rect 21118 12220 21138 12260
rect 21178 12220 21198 12260
rect 21118 12130 21198 12220
rect 21118 12070 21128 12130
rect 21188 12070 21198 12130
rect 21118 12060 21198 12070
rect 21318 12660 21398 12680
rect 21318 12620 21338 12660
rect 21378 12620 21398 12660
rect 21318 12560 21398 12620
rect 21318 12520 21338 12560
rect 21378 12520 21398 12560
rect 21318 12460 21398 12520
rect 21318 12420 21338 12460
rect 21378 12420 21398 12460
rect 21318 12360 21398 12420
rect 21318 12320 21338 12360
rect 21378 12320 21398 12360
rect 21318 12260 21398 12320
rect 21318 12220 21338 12260
rect 21378 12220 21398 12260
rect 20918 11990 21078 12000
rect 20918 11930 20928 11990
rect 20988 11930 21008 11990
rect 21068 11930 21078 11990
rect 20918 11920 21078 11930
rect 21318 11990 21398 12220
rect 21318 11930 21328 11990
rect 21388 11930 21398 11990
rect 21318 11920 21398 11930
rect 21518 12660 21598 12680
rect 21518 12620 21538 12660
rect 21578 12620 21598 12660
rect 21518 12560 21598 12620
rect 21518 12520 21538 12560
rect 21578 12520 21598 12560
rect 21518 12460 21598 12520
rect 21518 12420 21538 12460
rect 21578 12420 21598 12460
rect 21518 12360 21598 12420
rect 21518 12320 21538 12360
rect 21578 12320 21598 12360
rect 21518 12260 21598 12320
rect 21518 12220 21538 12260
rect 21578 12220 21598 12260
rect 21518 12140 21598 12220
rect 21518 12100 21538 12140
rect 21578 12100 21598 12140
rect 21518 11990 21598 12100
rect 23218 12503 23298 12520
rect 23218 12106 23238 12503
rect 23276 12106 23298 12503
rect 21518 11930 21528 11990
rect 21588 11930 21598 11990
rect 21518 11920 21598 11930
rect 22118 11990 22198 12000
rect 22118 11930 22128 11990
rect 22188 11930 22198 11990
rect 22118 11920 22198 11930
rect 19918 11820 19928 11880
rect 19988 11820 19998 11880
rect 19918 11810 19998 11820
rect 19448 11710 19528 11730
rect 19448 11670 19468 11710
rect 19508 11670 19528 11710
rect 19448 11610 19528 11670
rect 19448 11570 19468 11610
rect 19508 11570 19528 11610
rect 19448 11550 19528 11570
rect 19578 11710 19658 11730
rect 19578 11670 19598 11710
rect 19638 11670 19658 11710
rect 19578 11610 19658 11670
rect 19578 11570 19598 11610
rect 19638 11570 19658 11610
rect 19578 11550 19658 11570
rect 19708 11710 19788 11730
rect 19708 11670 19728 11710
rect 19768 11670 19788 11710
rect 19708 11610 19788 11670
rect 19708 11570 19728 11610
rect 19768 11570 19788 11610
rect 19708 11550 19788 11570
rect 19838 11710 19918 11730
rect 19838 11670 19858 11710
rect 19898 11670 19918 11710
rect 19838 11610 19918 11670
rect 19838 11570 19858 11610
rect 19898 11570 19918 11610
rect 19838 11550 19918 11570
rect 19968 11710 20048 11730
rect 19968 11670 19988 11710
rect 20028 11670 20048 11710
rect 19968 11610 20048 11670
rect 19968 11570 19988 11610
rect 20028 11570 20048 11610
rect 19968 11550 20048 11570
rect 20098 11710 20178 11730
rect 20098 11670 20118 11710
rect 20158 11670 20178 11710
rect 20098 11610 20178 11670
rect 20098 11570 20118 11610
rect 20158 11570 20178 11610
rect 20098 11550 20178 11570
rect 20228 11710 20308 11730
rect 20228 11670 20248 11710
rect 20288 11670 20308 11710
rect 20228 11610 20308 11670
rect 20228 11570 20248 11610
rect 20288 11570 20308 11610
rect 20228 11550 20308 11570
rect 20588 11710 20668 11730
rect 20588 11670 20608 11710
rect 20648 11670 20668 11710
rect 20588 11610 20668 11670
rect 20588 11570 20608 11610
rect 20648 11570 20668 11610
rect 20588 11550 20668 11570
rect 20718 11710 20798 11730
rect 20718 11670 20738 11710
rect 20778 11670 20798 11710
rect 20718 11610 20798 11670
rect 20718 11570 20738 11610
rect 20778 11570 20798 11610
rect 20718 11550 20798 11570
rect 20848 11710 20928 11730
rect 20848 11670 20868 11710
rect 20908 11670 20928 11710
rect 20848 11610 20928 11670
rect 20848 11570 20868 11610
rect 20908 11570 20928 11610
rect 19618 11500 19698 11510
rect 19618 11440 19628 11500
rect 19688 11440 19698 11500
rect 19618 11430 19698 11440
rect 19728 11170 19768 11550
rect 19988 11330 20028 11550
rect 20058 11500 20138 11510
rect 20058 11440 20068 11500
rect 20128 11440 20138 11500
rect 20058 11430 20138 11440
rect 20848 11480 20928 11570
rect 20978 11710 21058 11730
rect 20978 11670 20998 11710
rect 21038 11670 21058 11710
rect 20978 11610 21058 11670
rect 20978 11570 20998 11610
rect 21038 11570 21058 11610
rect 20978 11550 21058 11570
rect 21108 11710 21188 11730
rect 21108 11670 21128 11710
rect 21168 11670 21188 11710
rect 21108 11610 21188 11670
rect 21108 11570 21128 11610
rect 21168 11570 21188 11610
rect 21108 11550 21188 11570
rect 21238 11710 21318 11730
rect 21238 11670 21258 11710
rect 21298 11670 21318 11710
rect 21238 11610 21318 11670
rect 21238 11570 21258 11610
rect 21298 11570 21318 11610
rect 21238 11550 21318 11570
rect 21368 11710 21448 11730
rect 21368 11670 21388 11710
rect 21428 11670 21448 11710
rect 21368 11610 21448 11670
rect 21368 11570 21388 11610
rect 21428 11570 21448 11610
rect 21368 11550 21448 11570
rect 20848 11440 20868 11480
rect 20908 11440 20928 11480
rect 19968 11270 19978 11330
rect 20038 11270 20048 11330
rect 19708 11150 19788 11170
rect 19708 11110 19728 11150
rect 19768 11110 19788 11150
rect 19448 11030 19528 11050
rect 19448 10990 19468 11030
rect 19508 10990 19528 11030
rect 19448 10970 19528 10990
rect 19578 11030 19658 11050
rect 19578 10990 19598 11030
rect 19638 10990 19658 11030
rect 19578 10970 19658 10990
rect 19708 11030 19788 11110
rect 19988 11090 20028 11270
rect 20078 11240 20118 11430
rect 20848 11420 20928 11440
rect 21128 11490 21168 11550
rect 21898 11500 21978 11510
rect 21128 11480 21208 11490
rect 21128 11420 21138 11480
rect 21198 11420 21208 11480
rect 21898 11440 21908 11500
rect 21968 11440 21978 11500
rect 21898 11430 21978 11440
rect 22738 11500 22818 11510
rect 22738 11440 22748 11500
rect 22808 11440 22818 11500
rect 22738 11430 22818 11440
rect 23218 11500 23298 12106
rect 23218 11440 23228 11500
rect 23288 11440 23298 11500
rect 23438 11580 23548 11600
rect 23438 11510 23458 11580
rect 23528 11510 23548 11580
rect 23438 11490 23548 11510
rect 23218 11430 23298 11440
rect 20718 11350 20728 11410
rect 20788 11350 20798 11410
rect 20058 11230 20138 11240
rect 20058 11170 20068 11230
rect 20128 11170 20138 11230
rect 20058 11160 20138 11170
rect 20758 11170 20798 11350
rect 20758 11160 20838 11170
rect 20758 11100 20768 11160
rect 20828 11100 20838 11160
rect 20758 11090 20838 11100
rect 19708 10990 19728 11030
rect 19768 10990 19788 11030
rect 19708 10970 19788 10990
rect 19838 11030 19918 11050
rect 19838 10990 19858 11030
rect 19898 10990 19918 11030
rect 19838 10970 19918 10990
rect 19968 11030 20048 11090
rect 20868 11050 20908 11420
rect 21128 11410 21208 11420
rect 21128 11050 21168 11410
rect 23608 11330 23688 11340
rect 21898 11280 21978 11290
rect 21898 11220 21908 11280
rect 21968 11220 21978 11280
rect 23608 11270 23618 11330
rect 23678 11270 23688 11330
rect 23608 11260 23688 11270
rect 25888 11330 25968 11340
rect 25888 11270 25898 11330
rect 25958 11270 25968 11330
rect 21898 11210 21978 11220
rect 21198 11160 21278 11170
rect 21198 11100 21208 11160
rect 21268 11100 21278 11160
rect 21198 11090 21278 11100
rect 22738 11160 22818 11170
rect 22738 11100 22748 11160
rect 22808 11100 22818 11160
rect 22738 11090 22818 11100
rect 23218 11160 23298 11170
rect 23218 11100 23228 11160
rect 23288 11100 23298 11160
rect 19968 10990 19988 11030
rect 20028 10990 20048 11030
rect 19968 10970 20048 10990
rect 20098 11030 20178 11050
rect 20098 10990 20118 11030
rect 20158 10990 20178 11030
rect 20098 10970 20178 10990
rect 20228 11030 20308 11050
rect 20228 10990 20248 11030
rect 20288 10990 20308 11030
rect 20228 10970 20308 10990
rect 20588 11030 20668 11050
rect 20588 10990 20608 11030
rect 20648 10990 20668 11030
rect 20588 10970 20668 10990
rect 20718 11030 20798 11050
rect 20718 10990 20738 11030
rect 20778 10990 20798 11030
rect 20718 10970 20798 10990
rect 20848 11030 20928 11050
rect 20848 10990 20868 11030
rect 20908 10990 20928 11030
rect 20848 10970 20928 10990
rect 20978 11030 21058 11050
rect 20978 10990 20998 11030
rect 21038 10990 21058 11030
rect 20978 10970 21058 10990
rect 21108 11030 21188 11050
rect 21108 10990 21128 11030
rect 21168 10990 21188 11030
rect 21108 10970 21188 10990
rect 21238 11030 21318 11050
rect 21238 10990 21258 11030
rect 21298 10990 21318 11030
rect 21238 10970 21318 10990
rect 21368 11030 21448 11050
rect 21368 10990 21388 11030
rect 21428 10990 21448 11030
rect 21368 10970 21448 10990
rect 20978 10880 21058 10890
rect 20978 10820 20988 10880
rect 21048 10820 21058 10880
rect 19398 10770 19478 10780
rect 19398 10710 19408 10770
rect 19468 10710 19478 10770
rect 19398 10610 19478 10710
rect 19398 10570 19418 10610
rect 19458 10570 19478 10610
rect 19398 10550 19478 10570
rect 19598 10770 19678 10780
rect 19598 10710 19608 10770
rect 19668 10710 19678 10770
rect 19598 10490 19678 10710
rect 19838 10770 19918 10780
rect 19838 10710 19848 10770
rect 19908 10710 19918 10770
rect 19838 10700 19918 10710
rect 19998 10770 20078 10780
rect 19998 10710 20008 10770
rect 20068 10710 20078 10770
rect 19598 10440 19618 10490
rect 19658 10440 19678 10490
rect 19598 10350 19678 10440
rect 19598 10300 19618 10350
rect 19658 10300 19678 10350
rect 19598 10280 19678 10300
rect 19998 10490 20078 10710
rect 19998 10440 20018 10490
rect 20058 10440 20078 10490
rect 19998 10350 20078 10440
rect 19998 10300 20018 10350
rect 20058 10300 20078 10350
rect 19998 10280 20078 10300
rect 20398 10770 20478 10780
rect 20398 10710 20408 10770
rect 20468 10710 20478 10770
rect 20398 10490 20478 10710
rect 20398 10440 20418 10490
rect 20458 10440 20478 10490
rect 20398 10350 20478 10440
rect 20398 10300 20418 10350
rect 20458 10300 20478 10350
rect 20398 10280 20478 10300
rect 20798 10770 20878 10780
rect 20798 10710 20808 10770
rect 20868 10710 20878 10770
rect 20798 10490 20878 10710
rect 20978 10660 21058 10820
rect 20978 10600 20988 10660
rect 21048 10600 21058 10660
rect 20978 10590 21058 10600
rect 21198 10770 21278 10780
rect 21198 10710 21208 10770
rect 21268 10710 21278 10770
rect 20798 10440 20818 10490
rect 20858 10440 20878 10490
rect 20798 10350 20878 10440
rect 20798 10300 20818 10350
rect 20858 10300 20878 10350
rect 20798 10280 20878 10300
rect 21198 10490 21278 10710
rect 21398 10770 21478 10780
rect 21398 10710 21408 10770
rect 21468 10710 21478 10770
rect 21398 10610 21478 10710
rect 22118 10770 22198 10780
rect 22118 10710 22128 10770
rect 22188 10710 22198 10770
rect 22118 10700 22198 10710
rect 21398 10570 21418 10610
rect 21458 10570 21478 10610
rect 21398 10550 21478 10570
rect 23218 10610 23298 11100
rect 23438 11070 23548 11090
rect 23438 11000 23458 11070
rect 23528 11000 23548 11070
rect 23438 10980 23548 11000
rect 21198 10440 21218 10490
rect 21258 10440 21278 10490
rect 21198 10350 21278 10440
rect 21198 10300 21218 10350
rect 21258 10300 21278 10350
rect 21198 10280 21278 10300
rect 23218 10213 23238 10610
rect 23276 10213 23298 10610
rect 23218 10200 23298 10213
rect 23232 10050 23282 10051
rect 19138 9990 19158 10030
rect 19198 9990 19218 10030
rect 19138 9970 19218 9990
rect 23218 10039 23298 10050
rect 23008 9650 23088 9660
rect 23008 9590 23018 9650
rect 23078 9590 23088 9650
rect 23008 9580 23088 9590
rect 23218 9642 23238 10039
rect 23276 9642 23298 10039
rect 23218 9150 23298 9642
rect 23208 9130 23308 9150
rect 23208 9070 23228 9130
rect 23288 9070 23308 9130
rect 23208 9050 23308 9070
rect 19028 8710 19038 8770
rect 19098 8710 19108 8770
rect 19028 8690 19108 8710
rect 19028 8630 19038 8690
rect 19098 8630 19108 8690
rect 19028 8610 19108 8630
rect 19028 8550 19038 8610
rect 19098 8550 19108 8610
rect 19028 8540 19108 8550
rect 19138 8500 19218 8510
rect 19138 8440 19148 8500
rect 19208 8440 19218 8500
rect 19138 7160 19218 8440
rect 25888 8500 25968 11270
rect 25888 8440 25898 8500
rect 25958 8440 25968 8500
rect 25888 8430 25968 8440
rect 25998 8770 26478 19420
rect 25998 8710 26008 8770
rect 26068 8710 26088 8770
rect 26148 8710 26168 8770
rect 26228 8710 26248 8770
rect 26308 8710 26328 8770
rect 26388 8710 26408 8770
rect 26468 8710 26478 8770
rect 25998 8690 26478 8710
rect 25998 8630 26008 8690
rect 26068 8630 26088 8690
rect 26148 8630 26168 8690
rect 26228 8630 26248 8690
rect 26308 8630 26328 8690
rect 26388 8630 26408 8690
rect 26468 8630 26478 8690
rect 25998 8610 26478 8630
rect 25998 8550 26008 8610
rect 26068 8550 26088 8610
rect 26148 8550 26168 8610
rect 26228 8550 26248 8610
rect 26308 8550 26328 8610
rect 26388 8550 26408 8610
rect 26468 8550 26478 8610
rect 23088 8380 23198 8400
rect 23088 8310 23108 8380
rect 23178 8310 23198 8380
rect 23088 8290 23198 8310
rect 19338 8230 19418 8240
rect 19338 8170 19348 8230
rect 19408 8170 19418 8230
rect 19338 8130 19418 8170
rect 19338 8090 19358 8130
rect 19398 8090 19418 8130
rect 19338 8010 19418 8090
rect 19338 7970 19358 8010
rect 19398 7970 19418 8010
rect 19338 7910 19418 7970
rect 19338 7870 19358 7910
rect 19398 7870 19418 7910
rect 19338 7810 19418 7870
rect 19338 7770 19358 7810
rect 19398 7770 19418 7810
rect 19338 7710 19418 7770
rect 19338 7670 19358 7710
rect 19398 7670 19418 7710
rect 19338 7650 19418 7670
rect 19558 8230 19638 8240
rect 19558 8170 19568 8230
rect 19628 8170 19638 8230
rect 19558 8010 19638 8170
rect 19998 8230 20078 8240
rect 19998 8170 20008 8230
rect 20068 8170 20078 8230
rect 19558 7970 19578 8010
rect 19618 7970 19638 8010
rect 19558 7910 19638 7970
rect 19558 7870 19578 7910
rect 19618 7870 19638 7910
rect 19558 7810 19638 7870
rect 19558 7770 19578 7810
rect 19618 7770 19638 7810
rect 19558 7710 19638 7770
rect 19558 7670 19578 7710
rect 19618 7670 19638 7710
rect 19558 7650 19638 7670
rect 19778 8010 19858 8030
rect 19778 7970 19798 8010
rect 19838 7970 19858 8010
rect 19778 7910 19858 7970
rect 19778 7870 19798 7910
rect 19838 7870 19858 7910
rect 19778 7810 19858 7870
rect 19778 7770 19798 7810
rect 19838 7770 19858 7810
rect 19778 7710 19858 7770
rect 19778 7670 19798 7710
rect 19838 7670 19858 7710
rect 19778 7650 19858 7670
rect 19998 8010 20078 8170
rect 20318 8230 20398 8240
rect 20318 8170 20328 8230
rect 20388 8170 20398 8230
rect 20318 8030 20398 8170
rect 20638 8230 20718 8240
rect 20638 8170 20648 8230
rect 20708 8170 20718 8230
rect 19998 7970 20018 8010
rect 20058 7970 20078 8010
rect 19998 7910 20078 7970
rect 19998 7870 20018 7910
rect 20058 7870 20078 7910
rect 19998 7810 20078 7870
rect 19998 7770 20018 7810
rect 20058 7770 20078 7810
rect 19998 7710 20078 7770
rect 19998 7670 20018 7710
rect 20058 7670 20078 7710
rect 19998 7650 20078 7670
rect 20218 8010 20498 8030
rect 20218 7970 20238 8010
rect 20278 7970 20338 8010
rect 20378 7970 20438 8010
rect 20478 7970 20498 8010
rect 20218 7910 20498 7970
rect 20218 7870 20238 7910
rect 20278 7870 20338 7910
rect 20378 7870 20438 7910
rect 20478 7870 20498 7910
rect 20218 7810 20498 7870
rect 20218 7770 20238 7810
rect 20278 7770 20338 7810
rect 20378 7770 20438 7810
rect 20478 7770 20498 7810
rect 20218 7710 20498 7770
rect 20218 7670 20238 7710
rect 20278 7670 20338 7710
rect 20378 7670 20438 7710
rect 20478 7670 20498 7710
rect 20218 7650 20498 7670
rect 20638 8010 20718 8170
rect 21078 8230 21158 8240
rect 21078 8170 21088 8230
rect 21148 8170 21158 8230
rect 20638 7970 20658 8010
rect 20698 7970 20718 8010
rect 20638 7910 20718 7970
rect 20638 7870 20658 7910
rect 20698 7870 20718 7910
rect 20638 7810 20718 7870
rect 20638 7770 20658 7810
rect 20698 7770 20718 7810
rect 20638 7710 20718 7770
rect 20638 7670 20658 7710
rect 20698 7670 20718 7710
rect 20638 7650 20718 7670
rect 20858 8010 20938 8030
rect 20858 7970 20878 8010
rect 20918 7970 20938 8010
rect 20858 7910 20938 7970
rect 20858 7870 20878 7910
rect 20918 7870 20938 7910
rect 20858 7810 20938 7870
rect 20858 7770 20878 7810
rect 20918 7770 20938 7810
rect 20858 7710 20938 7770
rect 20858 7670 20878 7710
rect 20918 7670 20938 7710
rect 19778 7600 19858 7620
rect 19778 7560 19798 7600
rect 19838 7560 19858 7600
rect 19778 7380 19858 7560
rect 19778 7320 19788 7380
rect 19848 7320 19858 7380
rect 19778 7310 19858 7320
rect 19138 7100 19148 7160
rect 19208 7100 19218 7160
rect 19138 7090 19218 7100
rect 20198 7160 20278 7170
rect 20198 7100 20208 7160
rect 20268 7100 20278 7160
rect 18918 6980 18928 7040
rect 18988 6980 18998 7040
rect 18918 6970 18998 6980
rect 19978 7040 20058 7050
rect 19978 6980 19988 7040
rect 20048 6980 20058 7040
rect 19538 6910 19618 6930
rect 19538 6870 19558 6910
rect 19598 6870 19618 6910
rect 19538 6810 19618 6870
rect 19538 6770 19558 6810
rect 19598 6770 19618 6810
rect 19538 6710 19618 6770
rect 19538 6670 19558 6710
rect 19598 6670 19618 6710
rect 19538 6610 19618 6670
rect 19538 6570 19558 6610
rect 19598 6570 19618 6610
rect 19538 6490 19618 6570
rect 19538 6450 19558 6490
rect 19598 6450 19618 6490
rect 19538 6390 19618 6450
rect 19538 6330 19548 6390
rect 19608 6330 19618 6390
rect 19538 6320 19618 6330
rect 19758 6910 19838 6930
rect 19758 6870 19778 6910
rect 19818 6870 19838 6910
rect 19758 6810 19838 6870
rect 19758 6770 19778 6810
rect 19818 6770 19838 6810
rect 19758 6710 19838 6770
rect 19758 6670 19778 6710
rect 19818 6670 19838 6710
rect 19758 6610 19838 6670
rect 19758 6570 19778 6610
rect 19818 6570 19838 6610
rect 19758 6390 19838 6570
rect 19978 6910 20058 6980
rect 20198 7030 20278 7100
rect 20198 6990 20218 7030
rect 20258 6990 20278 7030
rect 20198 6970 20278 6990
rect 20418 7040 20498 7050
rect 20418 6980 20428 7040
rect 20488 6980 20498 7040
rect 19978 6870 19998 6910
rect 20038 6870 20058 6910
rect 19978 6810 20058 6870
rect 19978 6770 19998 6810
rect 20038 6770 20058 6810
rect 19978 6710 20058 6770
rect 19978 6670 19998 6710
rect 20038 6670 20058 6710
rect 19978 6610 20058 6670
rect 19978 6570 19998 6610
rect 20038 6570 20058 6610
rect 19978 6550 20058 6570
rect 20198 6910 20278 6930
rect 20198 6870 20218 6910
rect 20258 6870 20278 6910
rect 20198 6810 20278 6870
rect 20198 6770 20218 6810
rect 20258 6770 20278 6810
rect 20198 6710 20278 6770
rect 20198 6670 20218 6710
rect 20258 6670 20278 6710
rect 20198 6610 20278 6670
rect 20198 6570 20218 6610
rect 20258 6570 20278 6610
rect 19758 6330 19768 6390
rect 19828 6330 19838 6390
rect 19758 6320 19838 6330
rect 20198 6390 20278 6570
rect 20418 6910 20498 6980
rect 20858 7040 20938 7670
rect 21078 8010 21158 8170
rect 21398 8230 21478 8240
rect 21398 8170 21408 8230
rect 21468 8170 21478 8230
rect 21398 8030 21478 8170
rect 21718 8230 21798 8240
rect 21718 8170 21728 8230
rect 21788 8170 21798 8230
rect 21078 7970 21098 8010
rect 21138 7970 21158 8010
rect 21078 7910 21158 7970
rect 21078 7870 21098 7910
rect 21138 7870 21158 7910
rect 21078 7810 21158 7870
rect 21078 7770 21098 7810
rect 21138 7770 21158 7810
rect 21078 7710 21158 7770
rect 21078 7670 21098 7710
rect 21138 7670 21158 7710
rect 21078 7650 21158 7670
rect 21298 8010 21578 8030
rect 21298 7970 21318 8010
rect 21358 7970 21418 8010
rect 21458 7970 21518 8010
rect 21558 7970 21578 8010
rect 21298 7910 21578 7970
rect 21298 7870 21318 7910
rect 21358 7870 21418 7910
rect 21458 7870 21518 7910
rect 21558 7870 21578 7910
rect 21298 7810 21578 7870
rect 21298 7770 21318 7810
rect 21358 7770 21418 7810
rect 21458 7770 21518 7810
rect 21558 7770 21578 7810
rect 21298 7710 21578 7770
rect 21298 7670 21318 7710
rect 21358 7670 21418 7710
rect 21458 7670 21518 7710
rect 21558 7670 21578 7710
rect 21298 7650 21578 7670
rect 21718 8010 21798 8170
rect 22158 8230 22238 8240
rect 22158 8170 22168 8230
rect 22228 8170 22238 8230
rect 21718 7970 21738 8010
rect 21778 7970 21798 8010
rect 21718 7910 21798 7970
rect 21718 7870 21738 7910
rect 21778 7870 21798 7910
rect 21718 7810 21798 7870
rect 21718 7770 21738 7810
rect 21778 7770 21798 7810
rect 21718 7710 21798 7770
rect 21718 7670 21738 7710
rect 21778 7670 21798 7710
rect 21718 7650 21798 7670
rect 21938 8010 22018 8030
rect 21938 7970 21958 8010
rect 21998 7970 22018 8010
rect 21938 7910 22018 7970
rect 21938 7870 21958 7910
rect 21998 7870 22018 7910
rect 21938 7810 22018 7870
rect 21938 7770 21958 7810
rect 21998 7770 22018 7810
rect 21938 7710 22018 7770
rect 21938 7670 21958 7710
rect 21998 7670 22018 7710
rect 21808 7570 21888 7580
rect 21808 7510 21818 7570
rect 21878 7510 21888 7570
rect 21808 7500 21888 7510
rect 21938 7320 22018 7670
rect 22158 8010 22238 8170
rect 22158 7970 22178 8010
rect 22218 7970 22238 8010
rect 22158 7910 22238 7970
rect 22158 7870 22178 7910
rect 22218 7870 22238 7910
rect 22158 7810 22238 7870
rect 22158 7770 22178 7810
rect 22218 7770 22238 7810
rect 22158 7710 22238 7770
rect 22158 7670 22178 7710
rect 22218 7670 22238 7710
rect 22158 7650 22238 7670
rect 22378 8230 22458 8240
rect 22378 8170 22388 8230
rect 22448 8170 22458 8230
rect 22378 8130 22458 8170
rect 22378 8090 22398 8130
rect 22438 8090 22458 8130
rect 22378 8010 22458 8090
rect 22378 7970 22398 8010
rect 22438 7970 22458 8010
rect 22378 7910 22458 7970
rect 22378 7870 22398 7910
rect 22438 7870 22458 7910
rect 22378 7810 22458 7870
rect 22378 7770 22398 7810
rect 22438 7770 22458 7810
rect 22378 7710 22458 7770
rect 22378 7670 22398 7710
rect 22438 7670 22458 7710
rect 22378 7650 22458 7670
rect 22738 7590 22848 7610
rect 22068 7570 22148 7580
rect 22068 7510 22078 7570
rect 22138 7510 22148 7570
rect 22068 7500 22148 7510
rect 22738 7520 22758 7590
rect 22828 7520 22848 7590
rect 22738 7500 22848 7520
rect 20858 6980 20868 7040
rect 20928 6980 20938 7040
rect 21368 7270 21448 7280
rect 21368 7210 21378 7270
rect 21438 7210 21448 7270
rect 21368 7070 21448 7210
rect 21368 7010 21378 7070
rect 21438 7010 21448 7070
rect 21938 7260 21948 7320
rect 22008 7260 22018 7320
rect 21368 7000 21448 7010
rect 21498 7040 21578 7050
rect 20858 6970 20938 6980
rect 21498 6980 21508 7040
rect 21568 6980 21578 7040
rect 20418 6870 20438 6910
rect 20478 6870 20498 6910
rect 20418 6810 20498 6870
rect 20418 6770 20438 6810
rect 20478 6770 20498 6810
rect 20418 6710 20498 6770
rect 20418 6670 20438 6710
rect 20478 6670 20498 6710
rect 20418 6610 20498 6670
rect 20418 6570 20438 6610
rect 20478 6570 20498 6610
rect 20418 6550 20498 6570
rect 20638 6910 20718 6930
rect 20638 6870 20658 6910
rect 20698 6870 20718 6910
rect 20638 6810 20718 6870
rect 20638 6770 20658 6810
rect 20698 6770 20718 6810
rect 20638 6710 20718 6770
rect 20638 6670 20658 6710
rect 20698 6670 20718 6710
rect 20638 6610 20718 6670
rect 20638 6570 20658 6610
rect 20698 6570 20718 6610
rect 20198 6330 20208 6390
rect 20268 6330 20278 6390
rect 20198 6320 20278 6330
rect 20638 6390 20718 6570
rect 20858 6910 21138 6930
rect 20858 6870 20878 6910
rect 20918 6870 20978 6910
rect 21018 6870 21078 6910
rect 21118 6870 21138 6910
rect 20858 6810 21138 6870
rect 20858 6770 20878 6810
rect 20918 6770 20978 6810
rect 21018 6770 21078 6810
rect 21118 6770 21138 6810
rect 20858 6710 21138 6770
rect 20858 6670 20878 6710
rect 20918 6670 20978 6710
rect 21018 6670 21078 6710
rect 21118 6670 21138 6710
rect 20858 6610 21138 6670
rect 20858 6570 20878 6610
rect 20918 6570 20978 6610
rect 21018 6570 21078 6610
rect 21118 6570 21138 6610
rect 20858 6550 21138 6570
rect 21278 6910 21358 6930
rect 21278 6870 21298 6910
rect 21338 6870 21358 6910
rect 21278 6810 21358 6870
rect 21278 6770 21298 6810
rect 21338 6770 21358 6810
rect 21278 6710 21358 6770
rect 21278 6670 21298 6710
rect 21338 6670 21358 6710
rect 21278 6610 21358 6670
rect 21278 6570 21298 6610
rect 21338 6570 21358 6610
rect 20638 6330 20648 6390
rect 20708 6330 20718 6390
rect 20638 6320 20718 6330
rect 20958 6390 21038 6550
rect 20958 6330 20968 6390
rect 21028 6330 21038 6390
rect 20958 6320 21038 6330
rect 21278 6390 21358 6570
rect 21498 6910 21578 6980
rect 21938 7040 22018 7260
rect 25998 7320 26478 8550
rect 25998 7260 26008 7320
rect 26068 7260 26088 7320
rect 26148 7260 26168 7320
rect 26228 7260 26248 7320
rect 26308 7260 26328 7320
rect 26388 7260 26408 7320
rect 26468 7260 26478 7320
rect 21938 6980 21948 7040
rect 22008 6980 22018 7040
rect 22068 7070 22148 7080
rect 22068 7010 22078 7070
rect 22138 7010 22148 7070
rect 22068 7000 22148 7010
rect 22738 7060 22848 7080
rect 21498 6870 21518 6910
rect 21558 6870 21578 6910
rect 21498 6810 21578 6870
rect 21498 6770 21518 6810
rect 21558 6770 21578 6810
rect 21498 6710 21578 6770
rect 21498 6670 21518 6710
rect 21558 6670 21578 6710
rect 21498 6610 21578 6670
rect 21498 6570 21518 6610
rect 21558 6570 21578 6610
rect 21498 6550 21578 6570
rect 21718 6910 21798 6930
rect 21718 6870 21738 6910
rect 21778 6870 21798 6910
rect 21718 6810 21798 6870
rect 21718 6770 21738 6810
rect 21778 6770 21798 6810
rect 21718 6710 21798 6770
rect 21718 6670 21738 6710
rect 21778 6670 21798 6710
rect 21718 6610 21798 6670
rect 21718 6570 21738 6610
rect 21778 6570 21798 6610
rect 21278 6330 21288 6390
rect 21348 6330 21358 6390
rect 21278 6320 21358 6330
rect 21718 6390 21798 6570
rect 21938 6910 22018 6980
rect 22738 6990 22758 7060
rect 22828 6990 22848 7060
rect 22738 6970 22848 6990
rect 21938 6870 21958 6910
rect 21998 6870 22018 6910
rect 21938 6810 22018 6870
rect 21938 6770 21958 6810
rect 21998 6770 22018 6810
rect 21938 6710 22018 6770
rect 21938 6670 21958 6710
rect 21998 6670 22018 6710
rect 21938 6610 22018 6670
rect 21938 6570 21958 6610
rect 21998 6570 22018 6610
rect 21938 6550 22018 6570
rect 22158 6910 22238 6930
rect 22158 6870 22178 6910
rect 22218 6870 22238 6910
rect 22158 6810 22238 6870
rect 22158 6770 22178 6810
rect 22218 6770 22238 6810
rect 22158 6710 22238 6770
rect 22158 6670 22178 6710
rect 22218 6670 22238 6710
rect 22158 6610 22238 6670
rect 22158 6570 22178 6610
rect 22218 6570 22238 6610
rect 21718 6330 21728 6390
rect 21788 6330 21798 6390
rect 21718 6320 21798 6330
rect 22158 6390 22238 6570
rect 22158 6330 22168 6390
rect 22228 6330 22238 6390
rect 22158 6320 22238 6330
rect 22378 6910 22458 6930
rect 22378 6870 22398 6910
rect 22438 6870 22458 6910
rect 22378 6810 22458 6870
rect 22378 6770 22398 6810
rect 22438 6770 22458 6810
rect 22378 6710 22458 6770
rect 22378 6670 22398 6710
rect 22438 6670 22458 6710
rect 22378 6610 22458 6670
rect 22378 6570 22398 6610
rect 22438 6570 22458 6610
rect 22378 6490 22458 6570
rect 22378 6450 22398 6490
rect 22438 6450 22458 6490
rect 22378 6390 22458 6450
rect 22378 6330 22388 6390
rect 22448 6330 22458 6390
rect 22378 6320 22458 6330
rect 18398 5990 18408 6050
rect 18468 5990 18478 6050
rect 18398 5980 18478 5990
rect 17688 5820 17698 5880
rect 17758 5820 17768 5880
rect 17688 5810 17768 5820
rect 22978 5880 23088 5900
rect 22978 5810 22998 5880
rect 23068 5810 23088 5880
rect 22978 5790 23088 5810
rect 23578 5640 23658 5650
rect 23578 5580 23588 5640
rect 23648 5580 23658 5640
rect 23578 5530 23658 5580
rect 23578 5490 23598 5530
rect 23638 5490 23658 5530
rect 23578 5470 23658 5490
rect 24098 5640 24178 5650
rect 24098 5580 24108 5640
rect 24168 5580 24178 5640
rect 24098 5530 24178 5580
rect 24098 5490 24118 5530
rect 24158 5490 24178 5530
rect 24098 5470 24178 5490
rect 24618 5640 24698 5650
rect 24618 5580 24628 5640
rect 24688 5580 24698 5640
rect 24618 5530 24698 5580
rect 24618 5490 24638 5530
rect 24678 5490 24698 5530
rect 24618 5470 24698 5490
rect 25138 5640 25218 5650
rect 25138 5580 25148 5640
rect 25208 5580 25218 5640
rect 25138 5530 25218 5580
rect 25138 5490 25158 5530
rect 25198 5490 25218 5530
rect 25138 5470 25218 5490
rect 23208 5400 23268 5420
rect 23208 5360 23218 5400
rect 23258 5360 23268 5400
rect 23208 5300 23268 5360
rect 23208 5260 23218 5300
rect 23258 5260 23268 5300
rect 23208 5200 23268 5260
rect 23208 5160 23218 5200
rect 23258 5160 23268 5200
rect 23208 5100 23268 5160
rect 23208 5060 23218 5100
rect 23258 5060 23268 5100
rect 23208 4710 23268 5060
rect 23588 5400 23648 5470
rect 23588 5360 23598 5400
rect 23638 5360 23648 5400
rect 23588 5300 23648 5360
rect 23588 5260 23598 5300
rect 23638 5260 23648 5300
rect 23588 5200 23648 5260
rect 23588 5160 23598 5200
rect 23638 5160 23648 5200
rect 23588 5100 23648 5160
rect 23588 5060 23598 5100
rect 23638 5060 23648 5100
rect 23388 4990 23468 5000
rect 23388 4930 23398 4990
rect 23458 4930 23468 4990
rect 23388 4920 23468 4930
rect 23588 4820 23648 5060
rect 23728 5400 23788 5420
rect 23728 5360 23738 5400
rect 23778 5360 23788 5400
rect 23728 5300 23788 5360
rect 23728 5260 23738 5300
rect 23778 5260 23788 5300
rect 23728 5200 23788 5260
rect 23728 5160 23738 5200
rect 23778 5160 23788 5200
rect 23728 5100 23788 5160
rect 23728 5060 23738 5100
rect 23778 5060 23788 5100
rect 23308 4810 23388 4820
rect 23308 4750 23318 4810
rect 23378 4750 23388 4810
rect 23308 4740 23388 4750
rect 23578 4810 23658 4820
rect 23578 4750 23588 4810
rect 23648 4750 23658 4810
rect 23578 4740 23658 4750
rect 23208 4670 23218 4710
rect 23258 4670 23268 4710
rect 23208 4610 23268 4670
rect 23208 4570 23218 4610
rect 23258 4570 23268 4610
rect 23208 4510 23268 4570
rect 23208 4470 23218 4510
rect 23258 4470 23268 4510
rect 23208 4410 23268 4470
rect 23208 4370 23218 4410
rect 23258 4370 23268 4410
rect 23208 4310 23268 4370
rect 23208 4270 23218 4310
rect 23258 4270 23268 4310
rect 23208 4210 23268 4270
rect 23208 4170 23218 4210
rect 23258 4170 23268 4210
rect 23208 4150 23268 4170
rect 23318 4710 23378 4740
rect 23318 4670 23328 4710
rect 23368 4670 23378 4710
rect 23318 4610 23378 4670
rect 23318 4570 23328 4610
rect 23368 4570 23378 4610
rect 23318 4510 23378 4570
rect 23318 4470 23328 4510
rect 23368 4470 23378 4510
rect 23318 4410 23378 4470
rect 23318 4370 23328 4410
rect 23368 4370 23378 4410
rect 23318 4310 23378 4370
rect 23318 4270 23328 4310
rect 23368 4270 23378 4310
rect 23318 4220 23378 4270
rect 23728 4710 23788 5060
rect 24108 5400 24168 5470
rect 24108 5360 24118 5400
rect 24158 5360 24168 5400
rect 24108 5300 24168 5360
rect 24108 5260 24118 5300
rect 24158 5260 24168 5300
rect 24108 5200 24168 5260
rect 24108 5160 24118 5200
rect 24158 5160 24168 5200
rect 24108 5100 24168 5160
rect 24108 5060 24118 5100
rect 24158 5060 24168 5100
rect 23908 4990 23988 5000
rect 23908 4930 23918 4990
rect 23978 4930 23988 4990
rect 23908 4920 23988 4930
rect 24108 4820 24168 5060
rect 24248 5400 24308 5420
rect 24248 5360 24258 5400
rect 24298 5360 24308 5400
rect 24248 5300 24308 5360
rect 24248 5260 24258 5300
rect 24298 5260 24308 5300
rect 24248 5200 24308 5260
rect 24248 5160 24258 5200
rect 24298 5160 24308 5200
rect 24248 5100 24308 5160
rect 24248 5060 24258 5100
rect 24298 5060 24308 5100
rect 23828 4810 23908 4820
rect 23828 4750 23838 4810
rect 23898 4750 23908 4810
rect 23828 4740 23908 4750
rect 24098 4810 24178 4820
rect 24098 4750 24108 4810
rect 24168 4750 24178 4810
rect 24098 4740 24178 4750
rect 23728 4670 23738 4710
rect 23778 4670 23788 4710
rect 23728 4610 23788 4670
rect 23728 4570 23738 4610
rect 23778 4570 23788 4610
rect 23728 4510 23788 4570
rect 23728 4470 23738 4510
rect 23778 4470 23788 4510
rect 23728 4410 23788 4470
rect 23728 4370 23738 4410
rect 23778 4370 23788 4410
rect 23728 4310 23788 4370
rect 23728 4270 23738 4310
rect 23778 4270 23788 4310
rect 23318 4150 23378 4160
rect 23408 4220 23488 4230
rect 23408 4160 23418 4220
rect 23478 4160 23488 4220
rect 23408 4150 23488 4160
rect 23208 3950 23248 4150
rect 23278 4100 23336 4110
rect 23278 4048 23282 4100
rect 23334 4048 23336 4100
rect 23278 4040 23336 4048
rect 23206 3930 23266 3950
rect 23206 3890 23216 3930
rect 23256 3890 23266 3930
rect 23206 3830 23266 3890
rect 23206 3790 23216 3830
rect 23256 3790 23266 3830
rect 12698 3740 12778 3750
rect 12698 3680 12708 3740
rect 12768 3680 12778 3740
rect 12698 3670 12778 3680
rect 13118 3740 13198 3750
rect 13118 3680 13128 3740
rect 13188 3680 13198 3740
rect 13118 3670 13198 3680
rect 13788 3740 13868 3750
rect 13788 3680 13798 3740
rect 13858 3680 13868 3740
rect 13788 3670 13868 3680
rect 14358 3740 14438 3750
rect 14358 3680 14368 3740
rect 14428 3680 14438 3740
rect 14358 3670 14438 3680
rect 15068 3740 15148 3750
rect 15068 3680 15078 3740
rect 15138 3680 15148 3740
rect 15068 3670 15148 3680
rect 15498 3740 15578 3750
rect 15498 3680 15508 3740
rect 15568 3680 15578 3740
rect 15498 3670 15578 3680
rect 15938 3740 16018 3750
rect 15938 3680 15948 3740
rect 16008 3680 16018 3740
rect 15938 3670 16018 3680
rect 16188 3740 16268 3750
rect 16188 3680 16198 3740
rect 16258 3680 16268 3740
rect 16188 3670 16268 3680
rect 16408 3740 16488 3750
rect 16408 3680 16418 3740
rect 16478 3680 16488 3740
rect 16408 3670 16488 3680
rect 16878 3740 16958 3750
rect 16878 3680 16888 3740
rect 16948 3680 16958 3740
rect 16878 3670 16958 3680
rect 17318 3740 17398 3750
rect 17318 3680 17328 3740
rect 17388 3680 17398 3740
rect 17318 3670 17398 3680
rect 17938 3740 18018 3750
rect 17938 3680 17948 3740
rect 18008 3680 18018 3740
rect 17938 3670 18018 3680
rect 18278 3740 18358 3750
rect 18278 3680 18288 3740
rect 18348 3680 18358 3740
rect 18278 3670 18358 3680
rect 18638 3740 18718 3750
rect 18638 3680 18648 3740
rect 18708 3680 18718 3740
rect 18638 3670 18718 3680
rect 19238 3740 19318 3750
rect 19238 3680 19248 3740
rect 19308 3680 19318 3740
rect 19238 3670 19318 3680
rect 19578 3740 19658 3750
rect 19578 3680 19588 3740
rect 19648 3680 19658 3740
rect 19578 3670 19658 3680
rect 19938 3740 20018 3750
rect 19938 3680 19948 3740
rect 20008 3680 20018 3740
rect 19938 3670 20018 3680
rect 20538 3740 20618 3750
rect 20538 3680 20548 3740
rect 20608 3680 20618 3740
rect 20538 3670 20618 3680
rect 20878 3740 20958 3750
rect 20878 3680 20888 3740
rect 20948 3680 20958 3740
rect 20878 3670 20958 3680
rect 21238 3740 21318 3750
rect 21238 3680 21248 3740
rect 21308 3680 21318 3740
rect 21238 3670 21318 3680
rect 21838 3740 21918 3750
rect 21838 3680 21848 3740
rect 21908 3680 21918 3740
rect 21838 3670 21918 3680
rect 22178 3740 22258 3750
rect 22178 3680 22188 3740
rect 22248 3680 22258 3740
rect 22178 3670 22258 3680
rect 22538 3740 22618 3750
rect 22538 3680 22548 3740
rect 22608 3680 22618 3740
rect 22538 3670 22618 3680
rect 23206 3730 23266 3790
rect 23206 3690 23216 3730
rect 23256 3690 23266 3730
rect 13018 3620 13098 3640
rect 13018 3580 13038 3620
rect 13078 3600 13098 3620
rect 13218 3620 13288 3640
rect 14138 3620 14218 3640
rect 13218 3600 13228 3620
rect 13078 3580 13228 3600
rect 13268 3580 13288 3620
rect 13018 3560 13288 3580
rect 13328 3600 13408 3620
rect 14138 3600 14158 3620
rect 13328 3560 13348 3600
rect 13388 3580 14158 3600
rect 14198 3580 14218 3620
rect 13388 3560 14218 3580
rect 14278 3620 14338 3640
rect 14278 3580 14288 3620
rect 14328 3600 14338 3620
rect 15398 3620 15478 3640
rect 14328 3580 14768 3600
rect 14278 3560 14768 3580
rect 15398 3580 15418 3620
rect 15458 3600 15478 3620
rect 15618 3620 15698 3640
rect 15618 3600 15638 3620
rect 15458 3580 15638 3600
rect 15678 3580 15698 3620
rect 15398 3560 15698 3580
rect 16748 3630 16828 3640
rect 16748 3590 16768 3630
rect 16808 3610 16828 3630
rect 17158 3630 17238 3640
rect 17158 3610 17178 3630
rect 16808 3590 17178 3610
rect 17218 3590 17238 3630
rect 16748 3570 17238 3590
rect 19108 3620 19188 3640
rect 19108 3580 19128 3620
rect 19168 3600 19188 3620
rect 19688 3620 19768 3640
rect 19688 3600 19708 3620
rect 19168 3580 19708 3600
rect 19748 3580 19768 3620
rect 19108 3560 19768 3580
rect 20408 3620 20488 3640
rect 20408 3580 20428 3620
rect 20468 3600 20488 3620
rect 20988 3620 21068 3640
rect 20988 3600 21008 3620
rect 20468 3580 21008 3600
rect 21048 3580 21068 3620
rect 20408 3560 21068 3580
rect 21708 3620 21788 3640
rect 21708 3580 21728 3620
rect 21768 3600 21788 3620
rect 22288 3620 22368 3640
rect 22288 3600 22308 3620
rect 21768 3580 22308 3600
rect 22348 3580 22368 3620
rect 21708 3560 22368 3580
rect 23206 3630 23266 3690
rect 23206 3590 23216 3630
rect 23256 3590 23266 3630
rect 23206 3570 23266 3590
rect 23318 3930 23378 3950
rect 23318 3890 23328 3930
rect 23368 3890 23378 3930
rect 23318 3830 23378 3890
rect 23318 3790 23328 3830
rect 23368 3790 23378 3830
rect 23318 3730 23378 3790
rect 23318 3690 23328 3730
rect 23368 3690 23378 3730
rect 23318 3630 23378 3690
rect 23318 3590 23328 3630
rect 23368 3590 23378 3630
rect 23318 3560 23378 3590
rect 13328 3540 13408 3560
rect 14728 3520 14768 3560
rect 19148 3520 19188 3560
rect 20448 3520 20488 3560
rect 21748 3520 21788 3560
rect 14728 3500 14808 3520
rect 14728 3460 14748 3500
rect 14788 3460 14808 3500
rect 23250 3512 23308 3530
rect 23250 3478 23262 3512
rect 23296 3478 23308 3512
rect 23250 3460 23308 3478
rect 14728 3440 14808 3460
rect 23258 3420 23308 3460
rect 22808 3410 23048 3420
rect 22808 3350 22818 3410
rect 22878 3350 22898 3410
rect 22958 3350 22978 3410
rect 23038 3350 23048 3410
rect 12108 3280 12118 3340
rect 12178 3280 12188 3340
rect 12108 3270 12188 3280
rect 12318 3340 12398 3350
rect 22808 3340 23048 3350
rect 12318 3280 12328 3340
rect 12388 3280 12398 3340
rect 22750 3330 23048 3340
rect 16228 3310 16308 3330
rect 12318 3270 12398 3280
rect 13988 3300 14588 3310
rect 13988 3260 14008 3300
rect 14048 3270 14528 3300
rect 14048 3260 14068 3270
rect 13988 3240 14068 3260
rect 14508 3260 14528 3270
rect 14568 3260 14588 3300
rect 14508 3240 14588 3260
rect 16228 3270 16248 3310
rect 16288 3270 16308 3310
rect 16228 3250 16308 3270
rect 22750 3278 22754 3330
rect 22806 3278 22818 3330
rect 22750 3270 22818 3278
rect 22878 3270 22898 3330
rect 22958 3270 22978 3330
rect 23038 3270 23048 3330
rect 22750 3260 23048 3270
rect 22808 3250 23048 3260
rect 13328 3080 13408 3100
rect 16228 3080 16268 3250
rect 22808 3190 22818 3250
rect 22878 3190 22898 3250
rect 22958 3190 22978 3250
rect 23038 3190 23048 3250
rect 12378 3060 12458 3080
rect 13328 3060 13348 3080
rect 12378 3020 12398 3060
rect 12438 3040 13348 3060
rect 13388 3040 13408 3080
rect 12438 3020 13408 3040
rect 13458 3070 13538 3080
rect 13458 3030 13478 3070
rect 13518 3050 13538 3070
rect 14398 3070 14478 3080
rect 14398 3050 14418 3070
rect 13518 3030 14418 3050
rect 14458 3050 14478 3070
rect 15958 3070 16038 3080
rect 15958 3050 15978 3070
rect 14458 3030 15978 3050
rect 16018 3030 16038 3070
rect 16228 3060 18638 3080
rect 16228 3040 18582 3060
rect 12378 3000 12458 3020
rect 13458 3010 16038 3030
rect 18572 3020 18582 3040
rect 18622 3020 18638 3060
rect 18572 3000 18638 3020
rect 12538 2960 12618 2970
rect 12538 2900 12548 2960
rect 12608 2900 12618 2960
rect 12538 2890 12618 2900
rect 12758 2960 12838 2970
rect 12758 2900 12768 2960
rect 12828 2900 12838 2960
rect 12758 2890 12838 2900
rect 13228 2960 13308 2970
rect 13228 2900 13238 2960
rect 13298 2900 13308 2960
rect 13228 2890 13308 2900
rect 13568 2960 13648 2970
rect 13568 2900 13578 2960
rect 13638 2900 13648 2960
rect 13568 2890 13648 2900
rect 13788 2960 13868 2970
rect 13788 2900 13798 2960
rect 13858 2900 13868 2960
rect 13788 2890 13868 2900
rect 14228 2960 14308 2970
rect 14228 2900 14238 2960
rect 14298 2900 14308 2960
rect 14228 2890 14308 2900
rect 14908 2960 14988 2970
rect 14908 2900 14918 2960
rect 14978 2900 14988 2960
rect 14908 2890 14988 2900
rect 15128 2960 15208 2970
rect 15128 2900 15138 2960
rect 15198 2900 15208 2960
rect 15128 2890 15208 2900
rect 15598 2960 15678 2970
rect 15598 2900 15608 2960
rect 15668 2900 15678 2960
rect 15598 2890 15678 2900
rect 16058 2960 16138 2970
rect 16058 2900 16068 2960
rect 16128 2900 16138 2960
rect 16058 2890 16138 2900
rect 16408 2960 16488 2970
rect 16408 2900 16418 2960
rect 16478 2900 16488 2960
rect 16408 2890 16488 2900
rect 16658 2960 16738 2970
rect 16658 2900 16668 2960
rect 16728 2900 16738 2960
rect 16658 2890 16738 2900
rect 16878 2960 16958 2970
rect 16878 2900 16888 2960
rect 16948 2900 16958 2960
rect 16878 2890 16958 2900
rect 17208 2960 17288 2970
rect 17208 2900 17218 2960
rect 17278 2900 17288 2960
rect 17208 2890 17288 2900
rect 17868 2960 17948 2970
rect 17868 2900 17878 2960
rect 17938 2900 17948 2960
rect 17868 2890 17948 2900
rect 18088 2960 18168 2970
rect 18088 2900 18098 2960
rect 18158 2900 18168 2960
rect 18088 2890 18168 2900
rect 18658 2960 18738 2970
rect 18658 2900 18668 2960
rect 18728 2900 18738 2960
rect 18658 2890 18738 2900
rect 18918 2960 18998 2970
rect 18918 2900 18928 2960
rect 18988 2900 18998 2960
rect 18918 2890 18998 2900
rect 19168 2960 19248 2970
rect 19168 2900 19178 2960
rect 19238 2900 19248 2960
rect 19168 2890 19248 2900
rect 19388 2960 19468 2970
rect 19388 2900 19398 2960
rect 19458 2900 19468 2960
rect 19388 2890 19468 2900
rect 19938 2960 20018 2970
rect 19938 2900 19948 2960
rect 20008 2900 20018 2960
rect 19938 2890 20018 2900
rect 20218 2960 20298 2970
rect 20218 2900 20228 2960
rect 20288 2900 20298 2960
rect 20218 2890 20298 2900
rect 20468 2960 20548 2970
rect 20468 2900 20478 2960
rect 20538 2900 20548 2960
rect 20468 2890 20548 2900
rect 20688 2960 20768 2970
rect 20688 2900 20698 2960
rect 20758 2900 20768 2960
rect 20688 2890 20768 2900
rect 21238 2960 21318 2970
rect 21238 2900 21248 2960
rect 21308 2900 21318 2960
rect 21238 2890 21318 2900
rect 21518 2960 21598 2970
rect 21518 2900 21528 2960
rect 21588 2900 21598 2960
rect 21518 2890 21598 2900
rect 21768 2960 21848 2970
rect 21768 2900 21778 2960
rect 21838 2900 21848 2960
rect 21768 2890 21848 2900
rect 21988 2960 22068 2970
rect 21988 2900 21998 2960
rect 22058 2900 22068 2960
rect 21988 2890 22068 2900
rect 22538 2960 22618 2970
rect 22538 2900 22548 2960
rect 22608 2900 22618 2960
rect 22538 2890 22618 2900
rect 22808 1830 23048 3190
rect 23248 3410 23308 3420
rect 23248 3330 23308 3350
rect 23248 3250 23308 3270
rect 23248 3180 23308 3190
rect 23258 3140 23308 3180
rect 23250 3122 23308 3140
rect 23250 3088 23262 3122
rect 23296 3088 23308 3122
rect 23250 3070 23308 3088
rect 23338 3420 23378 3560
rect 23338 3410 23398 3420
rect 23338 3330 23398 3350
rect 23338 3250 23398 3270
rect 23338 3180 23398 3190
rect 23338 3030 23378 3180
rect 23168 3010 23266 3030
rect 23168 2970 23216 3010
rect 23256 2970 23266 3010
rect 23168 2910 23266 2970
rect 23168 2870 23216 2910
rect 23256 2870 23266 2910
rect 23168 2850 23266 2870
rect 23318 3010 23378 3030
rect 23318 2970 23328 3010
rect 23368 2970 23378 3010
rect 23318 2910 23378 2970
rect 23318 2870 23328 2910
rect 23368 2870 23378 2910
rect 23318 2850 23378 2870
rect 23168 2800 23210 2850
rect 23168 2650 23208 2800
rect 23428 2770 23488 4150
rect 23728 4210 23788 4270
rect 23728 4170 23738 4210
rect 23778 4170 23788 4210
rect 23728 4150 23788 4170
rect 23838 4710 23898 4740
rect 23838 4670 23848 4710
rect 23888 4670 23898 4710
rect 23838 4610 23898 4670
rect 23838 4570 23848 4610
rect 23888 4570 23898 4610
rect 23838 4510 23898 4570
rect 23838 4470 23848 4510
rect 23888 4470 23898 4510
rect 23838 4410 23898 4470
rect 23838 4370 23848 4410
rect 23888 4370 23898 4410
rect 23838 4310 23898 4370
rect 23838 4270 23848 4310
rect 23888 4270 23898 4310
rect 23838 4220 23898 4270
rect 24248 4710 24308 5060
rect 24628 5400 24688 5470
rect 24628 5360 24638 5400
rect 24678 5360 24688 5400
rect 24628 5300 24688 5360
rect 24628 5260 24638 5300
rect 24678 5260 24688 5300
rect 24628 5200 24688 5260
rect 24628 5160 24638 5200
rect 24678 5160 24688 5200
rect 24628 5100 24688 5160
rect 24628 5060 24638 5100
rect 24678 5060 24688 5100
rect 24428 4990 24508 5000
rect 24428 4930 24438 4990
rect 24498 4930 24508 4990
rect 24428 4920 24508 4930
rect 24628 4820 24688 5060
rect 24768 5400 24828 5420
rect 24768 5360 24778 5400
rect 24818 5360 24828 5400
rect 24768 5300 24828 5360
rect 24768 5260 24778 5300
rect 24818 5260 24828 5300
rect 24768 5200 24828 5260
rect 24768 5160 24778 5200
rect 24818 5160 24828 5200
rect 24768 5100 24828 5160
rect 24768 5060 24778 5100
rect 24818 5060 24828 5100
rect 24768 4990 24828 5060
rect 25148 5400 25208 5470
rect 25148 5360 25158 5400
rect 25198 5360 25208 5400
rect 25148 5300 25208 5360
rect 25148 5260 25158 5300
rect 25198 5260 25208 5300
rect 25148 5200 25208 5260
rect 25148 5160 25158 5200
rect 25198 5160 25208 5200
rect 25148 5100 25208 5160
rect 25148 5060 25158 5100
rect 25198 5060 25208 5100
rect 25148 5040 25208 5060
rect 24768 4920 24828 4930
rect 24958 4990 25018 5000
rect 24348 4810 24428 4820
rect 24348 4750 24358 4810
rect 24418 4750 24428 4810
rect 24348 4740 24428 4750
rect 24618 4810 24698 4820
rect 24618 4750 24628 4810
rect 24688 4750 24698 4810
rect 24618 4740 24698 4750
rect 24248 4670 24258 4710
rect 24298 4670 24308 4710
rect 24248 4610 24308 4670
rect 24248 4570 24258 4610
rect 24298 4570 24308 4610
rect 24248 4510 24308 4570
rect 24248 4470 24258 4510
rect 24298 4470 24308 4510
rect 24248 4410 24308 4470
rect 24248 4370 24258 4410
rect 24298 4370 24308 4410
rect 24248 4310 24308 4370
rect 24248 4270 24258 4310
rect 24298 4270 24308 4310
rect 23838 4150 23898 4160
rect 23928 4220 24008 4230
rect 23928 4160 23938 4220
rect 23998 4160 24008 4220
rect 23928 4150 24008 4160
rect 23408 2760 23488 2770
rect 23278 2750 23336 2760
rect 23278 2698 23282 2750
rect 23334 2698 23336 2750
rect 23278 2690 23336 2698
rect 23408 2700 23418 2760
rect 23478 2700 23488 2760
rect 23408 2690 23488 2700
rect 23518 4100 23598 4110
rect 23518 4040 23528 4100
rect 23588 4040 23598 4100
rect 23168 2630 23268 2650
rect 23168 2590 23218 2630
rect 23258 2590 23268 2630
rect 23168 2530 23268 2590
rect 23168 2490 23218 2530
rect 23258 2490 23268 2530
rect 23168 2430 23268 2490
rect 23168 2390 23218 2430
rect 23258 2390 23268 2430
rect 23168 2370 23268 2390
rect 23318 2640 23418 2650
rect 23378 2580 23418 2640
rect 23318 2530 23418 2580
rect 23518 2640 23598 4040
rect 23728 3950 23768 4150
rect 23798 4100 23856 4110
rect 23798 4048 23802 4100
rect 23854 4048 23856 4100
rect 23798 4040 23856 4048
rect 23726 3930 23786 3950
rect 23726 3890 23736 3930
rect 23776 3890 23786 3930
rect 23726 3830 23786 3890
rect 23726 3790 23736 3830
rect 23776 3790 23786 3830
rect 23726 3730 23786 3790
rect 23726 3690 23736 3730
rect 23776 3690 23786 3730
rect 23726 3630 23786 3690
rect 23726 3590 23736 3630
rect 23776 3590 23786 3630
rect 23726 3570 23786 3590
rect 23838 3930 23898 3950
rect 23838 3890 23848 3930
rect 23888 3890 23898 3930
rect 23838 3830 23898 3890
rect 23838 3790 23848 3830
rect 23888 3790 23898 3830
rect 23838 3730 23898 3790
rect 23838 3690 23848 3730
rect 23888 3690 23898 3730
rect 23838 3630 23898 3690
rect 23838 3590 23848 3630
rect 23888 3590 23898 3630
rect 23838 3560 23898 3590
rect 23770 3512 23828 3530
rect 23770 3478 23782 3512
rect 23816 3478 23828 3512
rect 23770 3460 23828 3478
rect 23778 3420 23828 3460
rect 23768 3410 23828 3420
rect 23768 3330 23828 3350
rect 23768 3250 23828 3270
rect 23768 3180 23828 3190
rect 23778 3140 23828 3180
rect 23770 3122 23828 3140
rect 23770 3088 23782 3122
rect 23816 3088 23828 3122
rect 23770 3070 23828 3088
rect 23858 3420 23898 3560
rect 23858 3410 23918 3420
rect 23858 3330 23918 3350
rect 23858 3250 23918 3270
rect 23858 3180 23918 3190
rect 23858 3030 23898 3180
rect 23518 2580 23528 2640
rect 23588 2580 23598 2640
rect 23518 2570 23598 2580
rect 23688 3010 23786 3030
rect 23688 2970 23736 3010
rect 23776 2970 23786 3010
rect 23688 2910 23786 2970
rect 23688 2870 23736 2910
rect 23776 2870 23786 2910
rect 23688 2850 23786 2870
rect 23838 3010 23898 3030
rect 23838 2970 23848 3010
rect 23888 2970 23898 3010
rect 23838 2910 23898 2970
rect 23838 2870 23848 2910
rect 23888 2870 23898 2910
rect 23838 2850 23898 2870
rect 23688 2800 23730 2850
rect 23688 2650 23728 2800
rect 23948 2770 24008 4150
rect 24248 4210 24308 4270
rect 24248 4170 24258 4210
rect 24298 4170 24308 4210
rect 24248 4150 24308 4170
rect 24358 4710 24418 4740
rect 24358 4670 24368 4710
rect 24408 4670 24418 4710
rect 24358 4610 24418 4670
rect 24358 4570 24368 4610
rect 24408 4570 24418 4610
rect 24358 4510 24418 4570
rect 24358 4470 24368 4510
rect 24408 4470 24418 4510
rect 24358 4410 24418 4470
rect 24358 4370 24368 4410
rect 24408 4370 24418 4410
rect 24358 4310 24418 4370
rect 24358 4270 24368 4310
rect 24408 4270 24418 4310
rect 24358 4220 24418 4270
rect 24358 4150 24418 4160
rect 24448 4220 24528 4230
rect 24448 4160 24458 4220
rect 24518 4160 24528 4220
rect 24448 4150 24528 4160
rect 23928 2760 24008 2770
rect 23798 2750 23856 2760
rect 23798 2698 23802 2750
rect 23854 2698 23856 2750
rect 23798 2690 23856 2698
rect 23928 2700 23938 2760
rect 23998 2700 24008 2760
rect 23928 2690 24008 2700
rect 24038 4100 24118 4110
rect 24038 4040 24048 4100
rect 24108 4040 24118 4100
rect 23688 2630 23788 2650
rect 23688 2590 23738 2630
rect 23778 2590 23788 2630
rect 23318 2490 23328 2530
rect 23368 2490 23418 2530
rect 23318 2430 23418 2490
rect 23318 2390 23328 2430
rect 23368 2390 23418 2430
rect 23318 2370 23418 2390
rect 23168 2170 23208 2370
rect 23264 2270 23322 2280
rect 23264 2218 23268 2270
rect 23320 2218 23322 2270
rect 23264 2210 23322 2218
rect 23378 2170 23418 2370
rect 23168 2150 23268 2170
rect 23168 2110 23218 2150
rect 23258 2110 23268 2150
rect 23168 2050 23268 2110
rect 23168 2010 23218 2050
rect 23258 2010 23268 2050
rect 23168 1990 23268 2010
rect 23318 2150 23418 2170
rect 23318 2110 23328 2150
rect 23368 2110 23418 2150
rect 23318 2050 23418 2110
rect 23318 2010 23328 2050
rect 23368 2010 23418 2050
rect 23318 1990 23418 2010
rect 23688 2530 23788 2590
rect 23688 2490 23738 2530
rect 23778 2490 23788 2530
rect 23688 2430 23788 2490
rect 23688 2390 23738 2430
rect 23778 2390 23788 2430
rect 23688 2370 23788 2390
rect 23838 2640 23938 2650
rect 23898 2580 23938 2640
rect 23838 2530 23938 2580
rect 24038 2640 24118 4040
rect 24248 3950 24288 4150
rect 24318 4100 24376 4110
rect 24318 4048 24322 4100
rect 24374 4048 24376 4100
rect 24318 4040 24376 4048
rect 24246 3930 24306 3950
rect 24246 3890 24256 3930
rect 24296 3890 24306 3930
rect 24246 3830 24306 3890
rect 24246 3790 24256 3830
rect 24296 3790 24306 3830
rect 24246 3730 24306 3790
rect 24246 3690 24256 3730
rect 24296 3690 24306 3730
rect 24246 3630 24306 3690
rect 24246 3590 24256 3630
rect 24296 3590 24306 3630
rect 24246 3570 24306 3590
rect 24358 3930 24418 3950
rect 24358 3890 24368 3930
rect 24408 3890 24418 3930
rect 24358 3830 24418 3890
rect 24358 3790 24368 3830
rect 24408 3790 24418 3830
rect 24358 3730 24418 3790
rect 24358 3690 24368 3730
rect 24408 3690 24418 3730
rect 24358 3630 24418 3690
rect 24358 3590 24368 3630
rect 24408 3590 24418 3630
rect 24358 3560 24418 3590
rect 24290 3512 24348 3530
rect 24290 3478 24302 3512
rect 24336 3478 24348 3512
rect 24290 3460 24348 3478
rect 24298 3420 24348 3460
rect 24288 3410 24348 3420
rect 24288 3330 24348 3350
rect 24288 3250 24348 3270
rect 24288 3180 24348 3190
rect 24298 3140 24348 3180
rect 24290 3122 24348 3140
rect 24290 3088 24302 3122
rect 24336 3088 24348 3122
rect 24290 3070 24348 3088
rect 24378 3420 24418 3560
rect 24378 3410 24438 3420
rect 24378 3330 24438 3350
rect 24378 3250 24438 3270
rect 24378 3180 24438 3190
rect 24378 3030 24418 3180
rect 24038 2580 24048 2640
rect 24108 2580 24118 2640
rect 24038 2570 24118 2580
rect 24208 3010 24306 3030
rect 24208 2970 24256 3010
rect 24296 2970 24306 3010
rect 24208 2910 24306 2970
rect 24208 2870 24256 2910
rect 24296 2870 24306 2910
rect 24208 2850 24306 2870
rect 24358 3010 24418 3030
rect 24358 2970 24368 3010
rect 24408 2970 24418 3010
rect 24358 2910 24418 2970
rect 24358 2870 24368 2910
rect 24408 2870 24418 2910
rect 24358 2850 24418 2870
rect 24208 2800 24250 2850
rect 24208 2650 24248 2800
rect 24468 2770 24528 4150
rect 24448 2760 24528 2770
rect 24318 2750 24376 2760
rect 24318 2698 24322 2750
rect 24374 2698 24376 2750
rect 24318 2690 24376 2698
rect 24448 2700 24458 2760
rect 24518 2700 24528 2760
rect 24448 2690 24528 2700
rect 24558 4100 24638 4110
rect 24558 4040 24568 4100
rect 24628 4040 24638 4100
rect 24208 2630 24308 2650
rect 24208 2590 24258 2630
rect 24298 2590 24308 2630
rect 23838 2490 23848 2530
rect 23888 2490 23938 2530
rect 23838 2430 23938 2490
rect 23838 2390 23848 2430
rect 23888 2390 23938 2430
rect 23838 2370 23938 2390
rect 23688 2170 23728 2370
rect 23784 2270 23842 2280
rect 23784 2218 23788 2270
rect 23840 2218 23842 2270
rect 23784 2210 23842 2218
rect 23898 2170 23938 2370
rect 23688 2150 23788 2170
rect 23688 2110 23738 2150
rect 23778 2110 23788 2150
rect 23688 2050 23788 2110
rect 23688 2010 23738 2050
rect 23778 2010 23788 2050
rect 23688 1990 23788 2010
rect 23838 2150 23938 2170
rect 23838 2110 23848 2150
rect 23888 2110 23938 2150
rect 23838 2050 23938 2110
rect 23838 2010 23848 2050
rect 23888 2010 23938 2050
rect 23838 1990 23938 2010
rect 24208 2530 24308 2590
rect 24208 2490 24258 2530
rect 24298 2490 24308 2530
rect 24208 2430 24308 2490
rect 24208 2390 24258 2430
rect 24298 2390 24308 2430
rect 24208 2370 24308 2390
rect 24358 2640 24458 2650
rect 24418 2580 24458 2640
rect 24358 2530 24458 2580
rect 24558 2640 24638 4040
rect 24558 2580 24568 2640
rect 24628 2580 24638 2640
rect 24558 2570 24638 2580
rect 24358 2490 24368 2530
rect 24408 2490 24458 2530
rect 24358 2430 24458 2490
rect 24358 2390 24368 2430
rect 24408 2390 24458 2430
rect 24358 2370 24458 2390
rect 24208 2170 24248 2370
rect 24304 2270 24362 2280
rect 24304 2218 24308 2270
rect 24360 2218 24362 2270
rect 24304 2210 24362 2218
rect 24418 2170 24458 2370
rect 24872 2270 24930 2280
rect 24872 2218 24874 2270
rect 24926 2218 24930 2270
rect 24872 2210 24930 2218
rect 24208 2150 24308 2170
rect 24208 2110 24258 2150
rect 24298 2110 24308 2150
rect 24208 2050 24308 2110
rect 24208 2010 24258 2050
rect 24298 2010 24308 2050
rect 24208 1990 24308 2010
rect 24358 2150 24458 2170
rect 24358 2110 24368 2150
rect 24408 2110 24458 2150
rect 24358 2050 24458 2110
rect 24358 2010 24368 2050
rect 24408 2010 24458 2050
rect 24358 1990 24458 2010
rect 24848 2150 24908 2170
rect 24848 2110 24858 2150
rect 24898 2110 24908 2150
rect 24848 2050 24908 2110
rect 24848 2010 24858 2050
rect 24898 2010 24908 2050
rect 23318 1940 23378 1990
rect 23838 1940 23898 1990
rect 24358 1940 24418 1990
rect 24848 1940 24908 2010
rect 24958 2150 25018 4930
rect 24958 2110 24968 2150
rect 25008 2110 25018 2150
rect 24958 2050 25018 2110
rect 24958 2010 24968 2050
rect 25008 2010 25018 2050
rect 24958 1990 25018 2010
rect 25168 3410 25408 3420
rect 25168 3350 25178 3410
rect 25238 3350 25258 3410
rect 25318 3350 25338 3410
rect 25398 3350 25408 3410
rect 25168 3330 25408 3350
rect 25168 3270 25178 3330
rect 25238 3270 25258 3330
rect 25318 3270 25338 3330
rect 25398 3270 25408 3330
rect 25168 3250 25408 3270
rect 25168 3190 25178 3250
rect 25238 3190 25258 3250
rect 25318 3190 25338 3250
rect 25398 3190 25408 3250
rect 22808 1770 22818 1830
rect 22878 1770 22898 1830
rect 22958 1770 22978 1830
rect 23038 1770 23048 1830
rect 22808 1750 23048 1770
rect 22808 1690 22818 1750
rect 22878 1690 22898 1750
rect 22958 1690 22978 1750
rect 23038 1690 23048 1750
rect 22808 1670 23048 1690
rect 22808 1610 22818 1670
rect 22878 1610 22898 1670
rect 22958 1610 22978 1670
rect 23038 1610 23048 1670
rect 22808 1600 23048 1610
rect 23308 1920 23388 1940
rect 23308 1880 23328 1920
rect 23368 1880 23388 1920
rect 23308 1560 23388 1880
rect 23308 1500 23318 1560
rect 23378 1500 23388 1560
rect 23308 1490 23388 1500
rect 23828 1920 23908 1940
rect 23828 1880 23848 1920
rect 23888 1880 23908 1920
rect 23828 1560 23908 1880
rect 23828 1500 23838 1560
rect 23898 1500 23908 1560
rect 23828 1490 23908 1500
rect 24348 1920 24428 1940
rect 24348 1880 24368 1920
rect 24408 1880 24428 1920
rect 24348 1560 24428 1880
rect 24348 1500 24358 1560
rect 24418 1500 24428 1560
rect 24348 1490 24428 1500
rect 24838 1920 24918 1940
rect 24838 1880 24858 1920
rect 24898 1880 24918 1920
rect 24838 1560 24918 1880
rect 25168 1830 25408 3190
rect 25998 2280 26478 7260
rect 25998 2220 26008 2280
rect 26068 2220 26088 2280
rect 26148 2220 26168 2280
rect 26228 2220 26248 2280
rect 26308 2220 26328 2280
rect 26388 2220 26408 2280
rect 26468 2220 26478 2280
rect 25998 2210 26478 2220
rect 25168 1770 25178 1830
rect 25238 1770 25258 1830
rect 25318 1770 25338 1830
rect 25398 1770 25408 1830
rect 25168 1750 25408 1770
rect 25168 1690 25178 1750
rect 25238 1690 25258 1750
rect 25318 1690 25338 1750
rect 25398 1690 25408 1750
rect 25168 1670 25408 1690
rect 25168 1610 25178 1670
rect 25238 1610 25258 1670
rect 25318 1610 25338 1670
rect 25398 1610 25408 1670
rect 25168 1600 25408 1610
rect 24838 1500 24848 1560
rect 24908 1500 24918 1560
rect 24838 1490 24918 1500
rect 11938 1270 11948 1330
rect 12008 1270 12018 1330
rect 11938 1260 12018 1270
<< via1 >>
rect 16128 19680 16188 19690
rect 16128 19640 16138 19680
rect 16138 19640 16178 19680
rect 16178 19640 16188 19680
rect 16128 19630 16188 19640
rect 14998 19490 15408 19500
rect 14998 19452 15008 19490
rect 15008 19452 15405 19490
rect 15405 19452 15408 19490
rect 14998 19440 15408 19452
rect 16908 19490 17318 19500
rect 16908 19452 16911 19490
rect 16911 19452 17308 19490
rect 17308 19452 17318 19490
rect 16908 19440 17318 19452
rect 26008 19440 26068 19500
rect 26098 19440 26158 19500
rect 26198 19440 26258 19500
rect 26308 19440 26368 19500
rect 26408 19440 26468 19500
rect 8878 19130 8938 19190
rect 8458 19020 8518 19080
rect 8458 18940 8518 19000
rect 8458 18860 8518 18920
rect 8458 18043 8468 18440
rect 8468 18043 8506 18440
rect 8506 18043 8518 18440
rect 8458 18040 8518 18043
rect 8878 18390 8938 18450
rect 8878 18310 8938 18370
rect 8878 18220 8938 18280
rect 8878 18130 8938 18190
rect 8878 18050 8938 18110
rect 9248 19020 9308 19080
rect 9248 18940 9308 19000
rect 9248 18860 9308 18920
rect 10688 19020 10748 19080
rect 10688 18940 10748 19000
rect 10688 18860 10748 18920
rect 8458 11520 8518 11580
rect 9468 14150 9528 14210
rect 10358 14660 10418 14720
rect 9578 12460 9638 12520
rect 9578 11140 9638 11200
rect 9688 14430 9748 14490
rect 9688 12690 9748 12750
rect 9468 11030 9528 11090
rect 8458 9700 8518 9760
rect 10628 14320 10688 14380
rect 18198 19130 18258 19190
rect 13248 19070 13308 19080
rect 13248 19030 13258 19070
rect 13258 19030 13298 19070
rect 13298 19030 13308 19070
rect 13248 19020 13308 19030
rect 13248 18990 13308 19000
rect 13248 18950 13258 18990
rect 13258 18950 13298 18990
rect 13298 18950 13308 18990
rect 13248 18940 13308 18950
rect 13248 18910 13308 18920
rect 13248 18870 13258 18910
rect 13258 18870 13298 18910
rect 13298 18870 13308 18910
rect 13248 18860 13308 18870
rect 15678 19020 15738 19080
rect 15678 18940 15738 19000
rect 15678 18860 15738 18920
rect 16788 19020 16848 19080
rect 16788 18940 16848 19000
rect 16788 18860 16848 18920
rect 17578 19020 17638 19080
rect 17578 18940 17638 19000
rect 17578 18860 17638 18920
rect 18198 18790 18258 18850
rect 17578 18043 17588 18440
rect 17588 18043 17626 18440
rect 17626 18043 17638 18440
rect 17578 18040 17638 18043
rect 17958 18390 18018 18450
rect 17958 18310 18018 18370
rect 17958 18220 18018 18280
rect 17958 18130 18018 18190
rect 17958 18050 18018 18110
rect 18658 18090 18718 18150
rect 11148 16750 11208 16810
rect 11578 16750 11638 16810
rect 13248 16754 13308 16810
rect 13248 16750 13252 16754
rect 13252 16750 13308 16754
rect 15348 16750 15408 16810
rect 15348 14740 15408 14800
rect 16358 15290 16418 15350
rect 16438 15290 16498 15350
rect 16518 15290 16578 15350
rect 16008 14740 16068 14800
rect 16248 14740 16308 14800
rect 13958 14660 14018 14720
rect 11148 14550 11208 14610
rect 12550 14600 12620 14610
rect 12550 14550 12560 14600
rect 12560 14550 12610 14600
rect 12610 14550 12620 14600
rect 12550 14540 12620 14550
rect 13948 14600 14018 14610
rect 13948 14550 13958 14600
rect 13958 14550 14008 14600
rect 14008 14550 14018 14600
rect 13948 14540 14018 14550
rect 16158 14540 16218 14600
rect 11038 14320 11098 14380
rect 11088 14200 11148 14210
rect 11088 14160 11098 14200
rect 11098 14160 11138 14200
rect 11138 14160 11148 14200
rect 11088 14150 11148 14160
rect 15478 14240 15538 14250
rect 15478 14200 15488 14240
rect 15488 14200 15528 14240
rect 15528 14200 15538 14240
rect 15478 14190 15538 14200
rect 15478 14160 15538 14170
rect 15478 14120 15488 14160
rect 15488 14120 15528 14160
rect 15528 14120 15538 14160
rect 15478 14110 15538 14120
rect 11168 14030 11228 14040
rect 11168 13990 11178 14030
rect 11178 13990 11218 14030
rect 11218 13990 11228 14030
rect 11168 13980 11228 13990
rect 11328 14030 11388 14040
rect 11328 13990 11338 14030
rect 11338 13990 11378 14030
rect 11378 13990 11388 14030
rect 11328 13980 11388 13990
rect 11488 14030 11548 14040
rect 11488 13990 11498 14030
rect 11498 13990 11538 14030
rect 11538 13990 11548 14030
rect 11488 13980 11548 13990
rect 11648 14030 11708 14040
rect 11648 13990 11658 14030
rect 11658 13990 11698 14030
rect 11698 13990 11708 14030
rect 11648 13980 11708 13990
rect 11808 14030 11868 14040
rect 11808 13990 11818 14030
rect 11818 13990 11858 14030
rect 11858 13990 11868 14030
rect 11808 13980 11868 13990
rect 11968 14030 12028 14040
rect 11968 13990 11978 14030
rect 11978 13990 12018 14030
rect 12018 13990 12028 14030
rect 11968 13980 12028 13990
rect 12128 14030 12188 14040
rect 12128 13990 12138 14030
rect 12138 13990 12178 14030
rect 12178 13990 12188 14030
rect 12128 13980 12188 13990
rect 12288 14030 12348 14040
rect 12288 13990 12298 14030
rect 12298 13990 12338 14030
rect 12338 13990 12348 14030
rect 12288 13980 12348 13990
rect 12448 14030 12508 14040
rect 12448 13990 12458 14030
rect 12458 13990 12498 14030
rect 12498 13990 12508 14030
rect 12448 13980 12508 13990
rect 12608 14030 12668 14040
rect 12608 13990 12618 14030
rect 12618 13990 12658 14030
rect 12658 13990 12668 14030
rect 12608 13980 12668 13990
rect 12768 14030 12828 14040
rect 12768 13990 12778 14030
rect 12778 13990 12818 14030
rect 12818 13990 12828 14030
rect 12768 13980 12828 13990
rect 12928 14030 12988 14040
rect 12928 13990 12938 14030
rect 12938 13990 12978 14030
rect 12978 13990 12988 14030
rect 12928 13980 12988 13990
rect 13088 14030 13148 14040
rect 13088 13990 13098 14030
rect 13098 13990 13138 14030
rect 13138 13990 13148 14030
rect 13088 13980 13148 13990
rect 13248 14030 13308 14040
rect 13248 13990 13258 14030
rect 13258 13990 13298 14030
rect 13298 13990 13308 14030
rect 13248 13980 13308 13990
rect 13408 14030 13468 14040
rect 13408 13990 13418 14030
rect 13418 13990 13458 14030
rect 13458 13990 13468 14030
rect 13408 13980 13468 13990
rect 13568 14030 13628 14040
rect 13568 13990 13578 14030
rect 13578 13990 13618 14030
rect 13618 13990 13628 14030
rect 13568 13980 13628 13990
rect 13728 14030 13788 14040
rect 13728 13990 13738 14030
rect 13738 13990 13778 14030
rect 13778 13990 13788 14030
rect 13728 13980 13788 13990
rect 13888 14030 13948 14040
rect 13888 13990 13898 14030
rect 13898 13990 13938 14030
rect 13938 13990 13948 14030
rect 13888 13980 13948 13990
rect 14048 14030 14108 14040
rect 14048 13990 14058 14030
rect 14058 13990 14098 14030
rect 14098 13990 14108 14030
rect 14048 13980 14108 13990
rect 14208 14030 14268 14040
rect 14208 13990 14218 14030
rect 14218 13990 14258 14030
rect 14258 13990 14268 14030
rect 14208 13980 14268 13990
rect 14368 14030 14428 14040
rect 14368 13990 14378 14030
rect 14378 13990 14418 14030
rect 14418 13990 14428 14030
rect 14368 13980 14428 13990
rect 14528 14030 14588 14040
rect 14528 13990 14538 14030
rect 14538 13990 14578 14030
rect 14578 13990 14588 14030
rect 14528 13980 14588 13990
rect 14688 14030 14748 14040
rect 14688 13990 14698 14030
rect 14698 13990 14738 14030
rect 14738 13990 14748 14030
rect 14688 13980 14748 13990
rect 14848 14030 14908 14040
rect 14848 13990 14858 14030
rect 14858 13990 14898 14030
rect 14898 13990 14908 14030
rect 14848 13980 14908 13990
rect 15008 14030 15068 14040
rect 15008 13990 15018 14030
rect 15018 13990 15058 14030
rect 15058 13990 15068 14030
rect 15008 13980 15068 13990
rect 15168 14030 15228 14040
rect 15168 13990 15178 14030
rect 15178 13990 15218 14030
rect 15218 13990 15228 14030
rect 15168 13980 15228 13990
rect 11908 13870 11968 13930
rect 11908 13790 11968 13850
rect 11908 13760 11968 13770
rect 11908 13720 11918 13760
rect 11918 13720 11958 13760
rect 11958 13720 11968 13760
rect 11908 13710 11968 13720
rect 13168 13870 13228 13930
rect 13248 13870 13308 13930
rect 13328 13870 13388 13930
rect 13168 13790 13228 13850
rect 13248 13790 13308 13850
rect 13328 13790 13388 13850
rect 13168 13710 13228 13770
rect 13248 13710 13308 13770
rect 13328 13710 13388 13770
rect 10928 13120 10988 13130
rect 10928 13080 10938 13120
rect 10938 13080 10978 13120
rect 10978 13080 10988 13120
rect 10928 13070 10988 13080
rect 10928 12990 10988 13050
rect 10928 12910 10988 12970
rect 11168 13120 11228 13130
rect 11168 13080 11178 13120
rect 11178 13080 11218 13120
rect 11218 13080 11228 13120
rect 11168 13070 11228 13080
rect 11168 12990 11228 13050
rect 11168 12910 11228 12970
rect 11408 13120 11468 13130
rect 11408 13080 11418 13120
rect 11418 13080 11458 13120
rect 11458 13080 11468 13120
rect 11408 13070 11468 13080
rect 11408 12990 11468 13050
rect 11408 12910 11468 12970
rect 11648 13120 11708 13130
rect 11648 13080 11658 13120
rect 11658 13080 11698 13120
rect 11698 13080 11708 13120
rect 11648 13070 11708 13080
rect 11648 12990 11708 13050
rect 11648 12910 11708 12970
rect 12288 13120 12348 13130
rect 12288 13080 12298 13120
rect 12298 13080 12338 13120
rect 12338 13080 12348 13120
rect 12288 13070 12348 13080
rect 12288 12990 12348 13050
rect 12288 12910 12348 12970
rect 12528 13120 12588 13130
rect 12528 13080 12538 13120
rect 12538 13080 12578 13120
rect 12578 13080 12588 13120
rect 12528 13070 12588 13080
rect 12528 12990 12588 13050
rect 12528 12910 12588 12970
rect 12768 13120 12828 13130
rect 12768 13080 12778 13120
rect 12778 13080 12818 13120
rect 12818 13080 12828 13120
rect 12768 13070 12828 13080
rect 12768 12990 12828 13050
rect 12768 12910 12828 12970
rect 10748 12800 10808 12860
rect 11498 12800 11558 12860
rect 11718 12800 11778 12860
rect 11978 12800 12038 12860
rect 12198 12800 12258 12860
rect 12458 12800 12518 12860
rect 11431 12742 11483 12750
rect 11431 12708 11441 12742
rect 11441 12708 11475 12742
rect 11475 12708 11483 12742
rect 11431 12698 11483 12708
rect 11791 12742 11843 12750
rect 11791 12708 11801 12742
rect 11801 12708 11835 12742
rect 11835 12708 11843 12742
rect 11791 12698 11843 12708
rect 11911 12742 11963 12750
rect 11911 12708 11921 12742
rect 11921 12708 11955 12742
rect 11955 12708 11963 12742
rect 11911 12698 11963 12708
rect 12271 12742 12323 12750
rect 12271 12708 12281 12742
rect 12281 12708 12315 12742
rect 12315 12708 12323 12742
rect 12271 12698 12323 12708
rect 12391 12742 12443 12750
rect 12391 12708 12401 12742
rect 12401 12708 12435 12742
rect 12435 12708 12443 12742
rect 12391 12698 12443 12708
rect 12808 12720 12868 12730
rect 12808 12680 12818 12720
rect 12818 12680 12858 12720
rect 12858 12680 12868 12720
rect 12808 12670 12868 12680
rect 12808 12640 12868 12650
rect 12808 12600 12818 12640
rect 12818 12600 12858 12640
rect 12858 12600 12868 12640
rect 12808 12590 12868 12600
rect 11534 12512 11586 12522
rect 11534 12478 11542 12512
rect 11542 12478 11576 12512
rect 11576 12478 11586 12512
rect 11534 12470 11586 12478
rect 11692 12512 11744 12522
rect 11692 12478 11700 12512
rect 11700 12478 11734 12512
rect 11734 12478 11744 12512
rect 11692 12470 11744 12478
rect 11608 12360 11668 12420
rect 11368 12250 11428 12310
rect 10628 11980 10688 12040
rect 10708 11980 10768 12040
rect 11128 11980 11188 12040
rect 11368 11980 11428 12040
rect 10888 11910 10948 11920
rect 10888 11870 10898 11910
rect 10898 11870 10938 11910
rect 10938 11870 10948 11910
rect 10888 11860 10948 11870
rect 10648 11520 10708 11580
rect 12016 12512 12068 12522
rect 12016 12478 12024 12512
rect 12024 12478 12058 12512
rect 12058 12478 12068 12512
rect 12016 12470 12068 12478
rect 12170 12512 12222 12522
rect 12170 12478 12178 12512
rect 12178 12478 12212 12512
rect 12212 12478 12222 12512
rect 12170 12470 12222 12478
rect 12088 12360 12148 12420
rect 12494 12512 12546 12522
rect 12494 12478 12502 12512
rect 12502 12478 12536 12512
rect 12536 12478 12546 12512
rect 12494 12470 12546 12478
rect 12808 12560 12868 12570
rect 12808 12520 12818 12560
rect 12818 12520 12858 12560
rect 12858 12520 12868 12560
rect 12808 12510 12868 12520
rect 12568 12360 12628 12420
rect 11848 12250 11908 12310
rect 12328 12250 12388 12310
rect 11848 11980 11908 12040
rect 12088 11980 12148 12040
rect 12568 11980 12628 12040
rect 12748 11980 12808 12040
rect 11608 11910 11668 11920
rect 11608 11870 11618 11910
rect 11618 11870 11658 11910
rect 11658 11870 11668 11910
rect 11608 11860 11668 11870
rect 11368 11520 11428 11580
rect 12328 11910 12388 11920
rect 12328 11870 12338 11910
rect 12338 11870 12378 11910
rect 12378 11870 12388 11910
rect 12328 11860 12388 11870
rect 12088 11520 12148 11580
rect 12808 11520 12868 11580
rect 14588 13870 14648 13930
rect 14588 13790 14648 13850
rect 14588 13760 14648 13770
rect 14588 13720 14598 13760
rect 14598 13720 14638 13760
rect 14638 13720 14648 13760
rect 14588 13710 14648 13720
rect 13168 12670 13228 12730
rect 13248 12670 13308 12730
rect 13328 12670 13388 12730
rect 13168 12590 13228 12650
rect 13248 12590 13308 12650
rect 13328 12590 13388 12650
rect 13168 12510 13228 12570
rect 13248 12510 13308 12570
rect 13328 12510 13388 12570
rect 13728 13120 13788 13130
rect 13728 13080 13738 13120
rect 13738 13080 13778 13120
rect 13778 13080 13788 13120
rect 13728 13070 13788 13080
rect 13728 12990 13788 13050
rect 13728 12910 13788 12970
rect 13968 13120 14028 13130
rect 13968 13080 13978 13120
rect 13978 13080 14018 13120
rect 14018 13080 14028 13120
rect 13968 13070 14028 13080
rect 13968 12990 14028 13050
rect 13968 12910 14028 12970
rect 14208 13120 14268 13130
rect 14208 13080 14218 13120
rect 14218 13080 14258 13120
rect 14258 13080 14268 13120
rect 14208 13070 14268 13080
rect 14208 12990 14268 13050
rect 14208 12910 14268 12970
rect 14848 13120 14908 13130
rect 14848 13080 14858 13120
rect 14858 13080 14898 13120
rect 14898 13080 14908 13120
rect 14848 13070 14908 13080
rect 14848 12990 14908 13050
rect 14848 12910 14908 12970
rect 15088 13120 15148 13130
rect 15088 13080 15098 13120
rect 15098 13080 15138 13120
rect 15138 13080 15148 13120
rect 15088 13070 15148 13080
rect 15088 12990 15148 13050
rect 15088 12910 15148 12970
rect 15328 13120 15388 13130
rect 15328 13080 15338 13120
rect 15338 13080 15378 13120
rect 15378 13080 15388 13120
rect 15328 13070 15388 13080
rect 15328 12990 15388 13050
rect 15328 12910 15388 12970
rect 15568 13120 15628 13130
rect 15568 13080 15578 13120
rect 15578 13080 15618 13120
rect 15618 13080 15628 13120
rect 15568 13070 15628 13080
rect 15568 12990 15628 13050
rect 15568 12910 15628 12970
rect 14038 12800 14098 12860
rect 14298 12800 14358 12860
rect 14518 12800 14578 12860
rect 14778 12800 14838 12860
rect 14998 12800 15058 12860
rect 15748 12800 15808 12860
rect 13688 12720 13748 12730
rect 13688 12680 13698 12720
rect 13698 12680 13738 12720
rect 13738 12680 13748 12720
rect 13688 12670 13748 12680
rect 14113 12742 14165 12750
rect 14113 12708 14121 12742
rect 14121 12708 14155 12742
rect 14155 12708 14165 12742
rect 14113 12698 14165 12708
rect 14233 12742 14285 12750
rect 14233 12708 14241 12742
rect 14241 12708 14275 12742
rect 14275 12708 14285 12742
rect 14233 12698 14285 12708
rect 14593 12742 14645 12750
rect 14593 12708 14601 12742
rect 14601 12708 14635 12742
rect 14635 12708 14645 12742
rect 14593 12698 14645 12708
rect 14713 12742 14765 12750
rect 14713 12708 14721 12742
rect 14721 12708 14755 12742
rect 14755 12708 14765 12742
rect 14713 12698 14765 12708
rect 15073 12742 15125 12750
rect 15073 12708 15081 12742
rect 15081 12708 15115 12742
rect 15115 12708 15125 12742
rect 15073 12698 15125 12708
rect 16158 12690 16218 12750
rect 13688 12640 13748 12650
rect 13688 12600 13698 12640
rect 13698 12600 13738 12640
rect 13738 12600 13748 12640
rect 13688 12590 13748 12600
rect 13688 12560 13748 12570
rect 13688 12520 13698 12560
rect 13698 12520 13738 12560
rect 13738 12520 13748 12560
rect 13688 12510 13748 12520
rect 14010 12512 14062 12522
rect 14010 12478 14020 12512
rect 14020 12478 14054 12512
rect 14054 12478 14062 12512
rect 14010 12470 14062 12478
rect 13928 12360 13988 12420
rect 14334 12512 14386 12522
rect 14334 12478 14344 12512
rect 14344 12478 14378 12512
rect 14378 12478 14386 12512
rect 14334 12470 14386 12478
rect 14488 12512 14540 12522
rect 14488 12478 14498 12512
rect 14498 12478 14532 12512
rect 14532 12478 14540 12512
rect 14488 12470 14540 12478
rect 14408 12360 14468 12420
rect 14812 12512 14864 12522
rect 14812 12478 14822 12512
rect 14822 12478 14856 12512
rect 14856 12478 14864 12512
rect 14812 12470 14864 12478
rect 14970 12512 15022 12522
rect 14970 12478 14980 12512
rect 14980 12478 15014 12512
rect 15014 12478 15022 12512
rect 14970 12470 15022 12478
rect 14888 12360 14948 12420
rect 14168 12250 14228 12310
rect 14648 12250 14708 12310
rect 13748 12140 13808 12200
rect 13748 12060 13808 12120
rect 13748 11980 13808 12040
rect 13928 12140 13988 12200
rect 13928 12060 13988 12120
rect 13928 11980 13988 12040
rect 14168 12140 14228 12200
rect 14168 12060 14228 12120
rect 14168 11980 14228 12040
rect 14408 12140 14468 12200
rect 14408 12060 14468 12120
rect 14408 11980 14468 12040
rect 14648 12140 14708 12200
rect 14648 12060 14708 12120
rect 14648 11980 14708 12040
rect 13068 11520 13128 11580
rect 13428 11520 13488 11580
rect 10528 11410 10588 11470
rect 10528 11330 10588 11390
rect 10528 11250 10588 11310
rect 10768 11410 10828 11470
rect 10768 11330 10828 11390
rect 10768 11250 10828 11310
rect 11008 11410 11068 11470
rect 11008 11330 11068 11390
rect 11008 11250 11068 11310
rect 11248 11410 11308 11470
rect 11248 11330 11308 11390
rect 11248 11250 11308 11310
rect 11488 11410 11548 11470
rect 11488 11330 11548 11390
rect 11488 11250 11548 11310
rect 11728 11410 11788 11470
rect 11728 11330 11788 11390
rect 11728 11250 11788 11310
rect 11968 11410 12028 11470
rect 11968 11330 12028 11390
rect 11968 11250 12028 11310
rect 12208 11410 12268 11470
rect 12208 11330 12268 11390
rect 12208 11250 12268 11310
rect 12448 11410 12508 11470
rect 12448 11330 12508 11390
rect 12448 11250 12508 11310
rect 12688 11410 12748 11470
rect 12688 11330 12748 11390
rect 12688 11250 12748 11310
rect 12928 11410 12988 11470
rect 12928 11330 12988 11390
rect 12928 11250 12988 11310
rect 11808 11140 11868 11200
rect 13248 11140 13308 11200
rect 12168 11030 12228 11090
rect 11898 10750 11958 10760
rect 11898 10710 11908 10750
rect 11908 10710 11948 10750
rect 11948 10710 11958 10750
rect 11898 10700 11958 10710
rect 12078 10750 12138 10760
rect 12078 10710 12088 10750
rect 12088 10710 12128 10750
rect 12128 10710 12138 10750
rect 12078 10700 12138 10710
rect 12528 10920 12588 10980
rect 12258 10750 12318 10760
rect 12258 10710 12268 10750
rect 12268 10710 12308 10750
rect 12308 10710 12318 10750
rect 12258 10700 12318 10710
rect 12438 10750 12498 10760
rect 12438 10710 12448 10750
rect 12448 10710 12488 10750
rect 12488 10710 12498 10750
rect 12438 10700 12498 10710
rect 12888 10810 12948 10870
rect 12618 10750 12678 10760
rect 12618 10710 12628 10750
rect 12628 10710 12668 10750
rect 12668 10710 12678 10750
rect 12618 10700 12678 10710
rect 12798 10750 12858 10760
rect 12798 10710 12808 10750
rect 12808 10710 12848 10750
rect 12848 10710 12858 10750
rect 12798 10700 12858 10710
rect 12978 10750 13038 10760
rect 12978 10710 12988 10750
rect 12988 10710 13028 10750
rect 13028 10710 13038 10750
rect 12978 10700 13038 10710
rect 13158 10750 13218 10760
rect 13158 10710 13168 10750
rect 13168 10710 13208 10750
rect 13208 10710 13218 10750
rect 13158 10700 13218 10710
rect 13688 11520 13748 11580
rect 14168 11910 14228 11920
rect 14168 11870 14178 11910
rect 14178 11870 14218 11910
rect 14218 11870 14228 11910
rect 14168 11860 14228 11870
rect 14408 11520 14468 11580
rect 15128 12250 15188 12310
rect 15128 12140 15188 12200
rect 15128 12060 15188 12120
rect 15128 11980 15188 12040
rect 15368 12140 15428 12200
rect 15368 12060 15428 12120
rect 15368 11980 15428 12040
rect 15788 12140 15848 12200
rect 15788 12060 15848 12120
rect 15788 11980 15848 12040
rect 14888 11910 14948 11920
rect 14888 11870 14898 11910
rect 14898 11870 14938 11910
rect 14938 11870 14948 11910
rect 14888 11860 14948 11870
rect 15128 11520 15188 11580
rect 15608 11910 15668 11920
rect 15608 11870 15618 11910
rect 15618 11870 15658 11910
rect 15658 11870 15668 11910
rect 15608 11860 15668 11870
rect 15848 11520 15908 11580
rect 13568 11410 13628 11470
rect 13568 11330 13628 11390
rect 13568 11250 13628 11310
rect 13808 11410 13868 11470
rect 13808 11330 13868 11390
rect 13808 11250 13868 11310
rect 14048 11410 14108 11470
rect 14048 11330 14108 11390
rect 14048 11250 14108 11310
rect 14288 11410 14348 11470
rect 14288 11330 14348 11390
rect 14288 11250 14348 11310
rect 14528 11410 14588 11470
rect 14528 11330 14588 11390
rect 14528 11250 14588 11310
rect 14768 11410 14828 11470
rect 14768 11330 14828 11390
rect 14768 11250 14828 11310
rect 15008 11410 15068 11470
rect 15008 11330 15068 11390
rect 15008 11250 15068 11310
rect 15248 11410 15308 11470
rect 15248 11330 15308 11390
rect 15248 11250 15308 11310
rect 15488 11410 15548 11470
rect 15488 11330 15548 11390
rect 15488 11250 15548 11310
rect 15728 11410 15788 11470
rect 15728 11330 15788 11390
rect 15728 11250 15788 11310
rect 14688 11140 14748 11200
rect 14328 11030 14388 11090
rect 13968 10920 14028 10980
rect 13608 10810 13668 10870
rect 13338 10750 13398 10760
rect 13338 10710 13348 10750
rect 13348 10710 13388 10750
rect 13388 10710 13398 10750
rect 13338 10700 13398 10710
rect 13428 10700 13488 10760
rect 13518 10750 13578 10760
rect 13518 10710 13528 10750
rect 13528 10710 13568 10750
rect 13568 10710 13578 10750
rect 13518 10700 13578 10710
rect 13698 10750 13758 10760
rect 13698 10710 13708 10750
rect 13708 10710 13748 10750
rect 13748 10710 13758 10750
rect 13698 10700 13758 10710
rect 13878 10750 13938 10760
rect 13878 10710 13888 10750
rect 13888 10710 13928 10750
rect 13928 10710 13938 10750
rect 13878 10700 13938 10710
rect 14058 10750 14118 10760
rect 14058 10710 14068 10750
rect 14068 10710 14108 10750
rect 14108 10710 14118 10750
rect 14058 10700 14118 10710
rect 14238 10750 14298 10760
rect 14238 10710 14248 10750
rect 14248 10710 14288 10750
rect 14288 10710 14298 10750
rect 14238 10700 14298 10710
rect 14418 10750 14478 10760
rect 14418 10710 14428 10750
rect 14428 10710 14468 10750
rect 14468 10710 14478 10750
rect 14418 10700 14478 10710
rect 14598 10750 14658 10760
rect 14598 10710 14608 10750
rect 14608 10710 14648 10750
rect 14648 10710 14658 10750
rect 14598 10700 14658 10710
rect 15718 11030 15778 11090
rect 15248 10920 15308 10980
rect 15598 10550 15658 10560
rect 15598 10510 15608 10550
rect 15608 10510 15648 10550
rect 15648 10510 15658 10550
rect 15598 10500 15658 10510
rect 15968 11410 16028 11470
rect 15968 11330 16028 11390
rect 15968 11250 16028 11310
rect 16248 12460 16308 12520
rect 16788 14430 16848 14490
rect 17578 16690 17638 16750
rect 16358 12140 16418 12200
rect 16438 12140 16498 12200
rect 16518 12140 16578 12200
rect 16358 12060 16418 12120
rect 16438 12060 16498 12120
rect 16518 12060 16578 12120
rect 16358 11980 16418 12040
rect 16438 11980 16498 12040
rect 16518 11980 16578 12040
rect 17958 15990 18018 16050
rect 18128 17390 18188 17450
rect 18798 16690 18858 16750
rect 18798 15290 18858 15350
rect 18658 14320 18718 14380
rect 23228 13450 23288 13510
rect 18078 13360 18138 13420
rect 18178 13360 18238 13420
rect 23018 13170 23078 13180
rect 23018 13130 23028 13170
rect 23028 13130 23068 13170
rect 23068 13130 23078 13170
rect 23018 13120 23078 13130
rect 17578 11520 17638 11580
rect 19148 12730 19208 12790
rect 19038 11350 19098 11410
rect 18928 11190 18988 11250
rect 16248 10920 16308 10980
rect 16158 10810 16218 10870
rect 15838 10550 15898 10560
rect 15838 10510 15848 10550
rect 15848 10510 15888 10550
rect 15888 10510 15898 10550
rect 15838 10500 15898 10510
rect 15248 10160 15308 10220
rect 15718 10210 15778 10220
rect 15718 10170 15728 10210
rect 15728 10170 15768 10210
rect 15768 10170 15778 10210
rect 15718 10160 15778 10170
rect 11628 10010 11688 10020
rect 11628 9970 11638 10010
rect 11638 9970 11678 10010
rect 11678 9970 11688 10010
rect 11628 9960 11688 9970
rect 11628 9880 11688 9940
rect 11628 9800 11688 9860
rect 11988 10010 12048 10020
rect 11988 9970 11998 10010
rect 11998 9970 12038 10010
rect 12038 9970 12048 10010
rect 11988 9960 12048 9970
rect 11988 9880 12048 9940
rect 11988 9800 12048 9860
rect 12348 10010 12408 10020
rect 12348 9970 12358 10010
rect 12358 9970 12398 10010
rect 12398 9970 12408 10010
rect 12348 9960 12408 9970
rect 12348 9880 12408 9940
rect 12348 9800 12408 9860
rect 12708 10010 12768 10020
rect 12708 9970 12718 10010
rect 12718 9970 12758 10010
rect 12758 9970 12768 10010
rect 12708 9960 12768 9970
rect 12708 9880 12768 9940
rect 12708 9800 12768 9860
rect 13068 10010 13128 10020
rect 13068 9970 13078 10010
rect 13078 9970 13118 10010
rect 13118 9970 13128 10010
rect 13068 9960 13128 9970
rect 13068 9880 13128 9940
rect 13068 9800 13128 9860
rect 13428 10010 13488 10020
rect 13428 9970 13438 10010
rect 13438 9970 13478 10010
rect 13478 9970 13488 10010
rect 13428 9960 13488 9970
rect 13428 9880 13488 9940
rect 13428 9800 13488 9860
rect 13788 10010 13848 10020
rect 13788 9970 13798 10010
rect 13798 9970 13838 10010
rect 13838 9970 13848 10010
rect 13788 9960 13848 9970
rect 13788 9880 13848 9940
rect 13788 9800 13848 9860
rect 14148 10010 14208 10020
rect 14148 9970 14158 10010
rect 14158 9970 14198 10010
rect 14198 9970 14208 10010
rect 14148 9960 14208 9970
rect 14148 9880 14208 9940
rect 14148 9800 14208 9860
rect 14508 10010 14568 10020
rect 14508 9970 14518 10010
rect 14518 9970 14558 10010
rect 14558 9970 14568 10010
rect 14508 9960 14568 9970
rect 14508 9880 14568 9940
rect 14508 9800 14568 9860
rect 14868 10010 14928 10020
rect 14868 9970 14878 10010
rect 14878 9970 14918 10010
rect 14918 9970 14928 10010
rect 14868 9960 14928 9970
rect 14868 9880 14928 9940
rect 14868 9800 14928 9860
rect 15498 9960 15558 10020
rect 15498 9880 15558 9940
rect 15498 9800 15558 9860
rect 15938 9960 15998 10020
rect 15938 9880 15998 9940
rect 15938 9800 15998 9860
rect 11806 9742 11858 9750
rect 11806 9708 11816 9742
rect 11816 9708 11850 9742
rect 11850 9708 11858 9742
rect 11806 9698 11858 9708
rect 11916 9742 11968 9750
rect 11916 9708 11926 9742
rect 11926 9708 11960 9742
rect 11960 9708 11968 9742
rect 11916 9698 11968 9708
rect 12026 9742 12078 9750
rect 12026 9708 12036 9742
rect 12036 9708 12070 9742
rect 12070 9708 12078 9742
rect 12026 9698 12078 9708
rect 12136 9742 12188 9750
rect 12136 9708 12146 9742
rect 12146 9708 12180 9742
rect 12180 9708 12188 9742
rect 12136 9698 12188 9708
rect 12246 9742 12298 9750
rect 12246 9708 12256 9742
rect 12256 9708 12290 9742
rect 12290 9708 12298 9742
rect 12246 9698 12298 9708
rect 12356 9742 12408 9750
rect 12356 9708 12366 9742
rect 12366 9708 12400 9742
rect 12400 9708 12408 9742
rect 12356 9698 12408 9708
rect 12466 9742 12518 9750
rect 12466 9708 12476 9742
rect 12476 9708 12510 9742
rect 12510 9708 12518 9742
rect 12466 9698 12518 9708
rect 12576 9742 12628 9750
rect 12576 9708 12586 9742
rect 12586 9708 12620 9742
rect 12620 9708 12628 9742
rect 12576 9698 12628 9708
rect 12686 9742 12738 9750
rect 12686 9708 12696 9742
rect 12696 9708 12730 9742
rect 12730 9708 12738 9742
rect 12686 9698 12738 9708
rect 12796 9742 12848 9750
rect 12796 9708 12806 9742
rect 12806 9708 12840 9742
rect 12840 9708 12848 9742
rect 12796 9698 12848 9708
rect 13706 9742 13758 9750
rect 13706 9708 13716 9742
rect 13716 9708 13750 9742
rect 13750 9708 13758 9742
rect 13706 9698 13758 9708
rect 13816 9742 13868 9750
rect 13816 9708 13826 9742
rect 13826 9708 13860 9742
rect 13860 9708 13868 9742
rect 13816 9698 13868 9708
rect 13926 9742 13978 9750
rect 13926 9708 13936 9742
rect 13936 9708 13970 9742
rect 13970 9708 13978 9742
rect 13926 9698 13978 9708
rect 14036 9742 14088 9750
rect 14036 9708 14046 9742
rect 14046 9708 14080 9742
rect 14080 9708 14088 9742
rect 14036 9698 14088 9708
rect 14146 9742 14198 9750
rect 14146 9708 14156 9742
rect 14156 9708 14190 9742
rect 14190 9708 14198 9742
rect 14146 9698 14198 9708
rect 14256 9742 14308 9750
rect 14256 9708 14266 9742
rect 14266 9708 14300 9742
rect 14300 9708 14308 9742
rect 14256 9698 14308 9708
rect 14366 9742 14418 9750
rect 14366 9708 14376 9742
rect 14376 9708 14410 9742
rect 14410 9708 14418 9742
rect 14366 9698 14418 9708
rect 14476 9742 14528 9750
rect 14476 9708 14486 9742
rect 14486 9708 14520 9742
rect 14520 9708 14528 9742
rect 14476 9698 14528 9708
rect 14586 9742 14638 9750
rect 14586 9708 14596 9742
rect 14596 9708 14630 9742
rect 14630 9708 14638 9742
rect 14586 9698 14638 9708
rect 14696 9742 14748 9750
rect 14696 9708 14706 9742
rect 14706 9708 14740 9742
rect 14740 9708 14748 9742
rect 14696 9698 14748 9708
rect 11638 9410 11698 9420
rect 11638 9370 11648 9410
rect 11648 9370 11688 9410
rect 11688 9370 11698 9410
rect 11638 9360 11698 9370
rect 11858 9360 11918 9420
rect 12078 9360 12138 9420
rect 12298 9360 12358 9420
rect 12518 9360 12578 9420
rect 12738 9360 12798 9420
rect 12958 9410 13018 9420
rect 12958 9370 12968 9410
rect 12968 9370 13008 9410
rect 13008 9370 13018 9410
rect 12958 9360 13018 9370
rect 13538 9410 13598 9420
rect 13538 9370 13548 9410
rect 13548 9370 13588 9410
rect 13588 9370 13598 9410
rect 13538 9360 13598 9370
rect 9688 9250 9748 9310
rect 11748 9250 11808 9310
rect 11968 9250 12028 9310
rect 12188 9250 12248 9310
rect 12408 9250 12468 9310
rect 12628 9250 12688 9310
rect 13758 9360 13818 9420
rect 13978 9360 14038 9420
rect 14198 9360 14258 9420
rect 14418 9360 14478 9420
rect 14638 9360 14698 9420
rect 14858 9410 14918 9420
rect 14858 9370 14868 9410
rect 14868 9370 14908 9410
rect 14908 9370 14918 9410
rect 14858 9360 14918 9370
rect 12848 9250 12908 9310
rect 13648 9240 13708 9300
rect 13648 9160 13708 9220
rect 13648 9080 13708 9140
rect 13868 9240 13928 9300
rect 13868 9160 13928 9220
rect 13868 9080 13928 9140
rect 14088 9240 14148 9300
rect 14088 9160 14148 9220
rect 14088 9080 14148 9140
rect 14308 9240 14368 9300
rect 14308 9160 14368 9220
rect 14308 9080 14368 9140
rect 14528 9240 14588 9300
rect 14528 9160 14588 9220
rect 14528 9080 14588 9140
rect 14748 9240 14808 9300
rect 14748 9160 14808 9220
rect 14748 9080 14808 9140
rect 18658 9240 18718 9300
rect 18738 9240 18798 9300
rect 18818 9240 18878 9300
rect 18658 9160 18718 9220
rect 18738 9160 18798 9220
rect 18818 9160 18878 9220
rect 18658 9080 18718 9140
rect 18738 9080 18798 9140
rect 18818 9080 18878 9140
rect 18108 8310 18168 8370
rect 13258 8290 13318 8300
rect 13258 8250 13268 8290
rect 13268 8250 13308 8290
rect 13308 8250 13318 8290
rect 13258 8240 13318 8250
rect 13478 8290 13538 8300
rect 13478 8250 13488 8290
rect 13488 8250 13528 8290
rect 13528 8250 13538 8290
rect 13478 8240 13538 8250
rect 13778 8290 13838 8300
rect 13778 8250 13788 8290
rect 13788 8250 13828 8290
rect 13828 8250 13838 8290
rect 13778 8240 13838 8250
rect 14008 8290 14068 8300
rect 14008 8250 14018 8290
rect 14018 8250 14058 8290
rect 14058 8250 14068 8290
rect 14008 8240 14068 8250
rect 14158 8290 14218 8300
rect 14158 8250 14168 8290
rect 14168 8250 14208 8290
rect 14208 8250 14218 8290
rect 14158 8240 14218 8250
rect 14378 8290 14438 8300
rect 14378 8250 14388 8290
rect 14388 8250 14428 8290
rect 14428 8250 14438 8290
rect 14378 8240 14438 8250
rect 14678 8290 14738 8300
rect 14678 8250 14688 8290
rect 14688 8250 14728 8290
rect 14728 8250 14738 8290
rect 14678 8240 14738 8250
rect 14898 8290 14958 8300
rect 14898 8250 14908 8290
rect 14908 8250 14948 8290
rect 14948 8250 14958 8290
rect 14898 8240 14958 8250
rect 15298 8290 15358 8300
rect 15298 8250 15308 8290
rect 15308 8250 15348 8290
rect 15348 8250 15358 8290
rect 15298 8240 15358 8250
rect 15628 8290 15688 8300
rect 15628 8250 15638 8290
rect 15638 8250 15678 8290
rect 15678 8250 15688 8290
rect 15628 8240 15688 8250
rect 15958 8290 16018 8300
rect 15958 8250 15968 8290
rect 15968 8250 16008 8290
rect 16008 8250 16018 8290
rect 15958 8240 16018 8250
rect 16398 8290 16458 8300
rect 16398 8250 16408 8290
rect 16408 8250 16448 8290
rect 16448 8250 16458 8290
rect 16398 8240 16458 8250
rect 16658 8240 16718 8300
rect 17178 8290 17238 8300
rect 17178 8250 17188 8290
rect 17188 8250 17228 8290
rect 17228 8250 17238 8290
rect 17178 8240 17238 8250
rect 17858 8290 17918 8300
rect 17858 8250 17868 8290
rect 17868 8250 17908 8290
rect 17908 8250 17918 8290
rect 17858 8240 17918 8250
rect 12118 7750 12178 7810
rect 11948 6370 12008 6430
rect 13138 7800 13198 7810
rect 13138 7760 13148 7800
rect 13148 7760 13188 7800
rect 13188 7760 13198 7800
rect 13138 7750 13198 7760
rect 15058 7790 15118 7800
rect 15058 7750 15068 7790
rect 15068 7750 15108 7790
rect 15108 7750 15118 7790
rect 15058 7740 15118 7750
rect 16088 7790 16148 7800
rect 16088 7750 16098 7790
rect 16098 7750 16138 7790
rect 16138 7750 16148 7790
rect 16088 7740 16148 7750
rect 13708 7220 13768 7230
rect 13708 7180 13718 7220
rect 13718 7180 13758 7220
rect 13758 7180 13768 7220
rect 13708 7170 13768 7180
rect 13258 7110 13318 7120
rect 13258 7070 13268 7110
rect 13268 7070 13308 7110
rect 13308 7070 13318 7110
rect 13258 7060 13318 7070
rect 13998 7110 14058 7120
rect 13998 7070 14008 7110
rect 14008 7070 14048 7110
rect 14048 7070 14058 7110
rect 13998 7060 14058 7070
rect 14158 7110 14218 7120
rect 14158 7070 14168 7110
rect 14168 7070 14208 7110
rect 14208 7070 14218 7110
rect 14158 7060 14218 7070
rect 14898 7110 14958 7120
rect 14898 7070 14908 7110
rect 14908 7070 14948 7110
rect 14948 7070 14958 7110
rect 14898 7060 14958 7070
rect 13138 6420 13198 6430
rect 13138 6380 13148 6420
rect 13148 6380 13188 6420
rect 13188 6380 13198 6420
rect 13138 6370 13198 6380
rect 15238 7170 15298 7230
rect 15148 7110 15208 7120
rect 15148 7070 15158 7110
rect 15158 7070 15198 7110
rect 15198 7070 15208 7110
rect 15148 7060 15208 7070
rect 15338 7110 15398 7120
rect 15338 7070 15348 7110
rect 15348 7070 15388 7110
rect 15388 7070 15398 7110
rect 15338 7060 15398 7070
rect 15418 7110 15478 7120
rect 15418 7070 15428 7110
rect 15428 7070 15468 7110
rect 15468 7070 15478 7110
rect 15418 7060 15478 7070
rect 15628 7110 15688 7120
rect 15628 7070 15638 7110
rect 15638 7070 15678 7110
rect 15678 7070 15688 7110
rect 15628 7060 15688 7070
rect 15958 7110 16018 7120
rect 15958 7070 15968 7110
rect 15968 7070 16008 7110
rect 16008 7070 16018 7110
rect 15958 7060 16018 7070
rect 15258 7000 15318 7010
rect 15258 6960 15268 7000
rect 15268 6960 15308 7000
rect 15308 6960 15318 7000
rect 15258 6950 15318 6960
rect 16238 7180 16298 7240
rect 16908 8180 16968 8190
rect 16908 8140 16918 8180
rect 16918 8140 16958 8180
rect 16958 8140 16968 8180
rect 16908 8130 16968 8140
rect 17538 8180 17598 8190
rect 17538 8140 17548 8180
rect 17548 8140 17588 8180
rect 17588 8140 17598 8180
rect 17538 8130 17598 8140
rect 18108 8130 18168 8190
rect 16658 7170 16718 7230
rect 16828 7220 16888 7230
rect 16828 7180 16838 7220
rect 16838 7180 16878 7220
rect 16878 7180 16888 7220
rect 16828 7170 16888 7180
rect 18008 7840 18068 7850
rect 18008 7800 18018 7840
rect 18018 7800 18058 7840
rect 18058 7800 18068 7840
rect 18008 7790 18068 7800
rect 18188 7790 18248 7850
rect 18188 7430 18248 7490
rect 18188 7320 18248 7380
rect 17468 7220 17528 7230
rect 17468 7180 17478 7220
rect 17478 7180 17518 7220
rect 17518 7180 17528 7220
rect 17468 7170 17528 7180
rect 18658 7320 18718 7380
rect 18738 7320 18798 7380
rect 18818 7320 18878 7380
rect 18188 7170 18248 7230
rect 18298 7210 18358 7270
rect 16398 7110 16458 7120
rect 16398 7070 16408 7110
rect 16408 7070 16448 7110
rect 16448 7070 16458 7110
rect 16398 7060 16458 7070
rect 16788 7110 16848 7120
rect 16788 7070 16798 7110
rect 16798 7070 16838 7110
rect 16838 7070 16848 7110
rect 16788 7060 16848 7070
rect 16998 7060 17058 7120
rect 17178 7110 17238 7120
rect 17178 7070 17188 7110
rect 17188 7070 17228 7110
rect 17228 7070 17238 7110
rect 17178 7060 17238 7070
rect 17858 7110 17918 7120
rect 17858 7070 17868 7110
rect 17868 7070 17908 7110
rect 17908 7070 17918 7110
rect 17858 7060 17918 7070
rect 15038 6390 15098 6400
rect 15038 6350 15048 6390
rect 15048 6350 15088 6390
rect 15088 6350 15098 6390
rect 15038 6340 15098 6350
rect 16128 6430 16188 6440
rect 16128 6390 16138 6430
rect 16138 6390 16178 6430
rect 16178 6390 16188 6430
rect 16128 6380 16188 6390
rect 17698 6460 17758 6470
rect 17698 6420 17708 6460
rect 17708 6420 17748 6460
rect 17748 6420 17758 6460
rect 17698 6410 17758 6420
rect 13668 6040 13728 6050
rect 13668 6000 13678 6040
rect 13678 6000 13718 6040
rect 13718 6000 13728 6040
rect 13668 5990 13728 6000
rect 15388 6040 15448 6050
rect 15388 6000 15398 6040
rect 15398 6000 15438 6040
rect 15438 6000 15448 6040
rect 15388 5990 15448 6000
rect 16238 6010 16298 6070
rect 17468 6040 17528 6050
rect 17468 6000 17478 6040
rect 17478 6000 17518 6040
rect 17518 6000 17528 6040
rect 17468 5990 17528 6000
rect 13258 5930 13318 5940
rect 13258 5890 13268 5930
rect 13268 5890 13308 5930
rect 13308 5890 13318 5930
rect 13258 5880 13318 5890
rect 13478 5930 13538 5940
rect 13478 5890 13488 5930
rect 13488 5890 13528 5930
rect 13528 5890 13538 5930
rect 13478 5880 13538 5890
rect 13778 5930 13838 5940
rect 13778 5890 13788 5930
rect 13788 5890 13828 5930
rect 13828 5890 13838 5930
rect 13778 5880 13838 5890
rect 13998 5930 14058 5940
rect 13998 5890 14008 5930
rect 14008 5890 14048 5930
rect 14048 5890 14058 5930
rect 13998 5880 14058 5890
rect 14158 5930 14218 5940
rect 14158 5890 14168 5930
rect 14168 5890 14208 5930
rect 14208 5890 14218 5930
rect 14158 5880 14218 5890
rect 14378 5930 14438 5940
rect 14378 5890 14388 5930
rect 14388 5890 14428 5930
rect 14428 5890 14438 5930
rect 14378 5880 14438 5890
rect 14678 5930 14738 5940
rect 14678 5890 14688 5930
rect 14688 5890 14728 5930
rect 14728 5890 14738 5930
rect 14678 5880 14738 5890
rect 14898 5930 14958 5940
rect 14898 5890 14908 5930
rect 14908 5890 14948 5930
rect 14948 5890 14958 5930
rect 14898 5880 14958 5890
rect 15198 5930 15258 5940
rect 15198 5890 15208 5930
rect 15208 5890 15248 5930
rect 15248 5890 15258 5930
rect 15198 5880 15258 5890
rect 15638 5930 15698 5940
rect 15638 5890 15648 5930
rect 15648 5890 15688 5930
rect 15688 5890 15698 5930
rect 15638 5880 15698 5890
rect 15968 5930 16028 5940
rect 15968 5890 15978 5930
rect 15978 5890 16018 5930
rect 16018 5890 16028 5930
rect 15968 5880 16028 5890
rect 16398 5930 16458 5940
rect 16398 5890 16408 5930
rect 16408 5890 16448 5930
rect 16448 5890 16458 5930
rect 16398 5880 16458 5890
rect 16788 5930 16848 5940
rect 16788 5890 16798 5930
rect 16798 5890 16838 5930
rect 16838 5890 16848 5930
rect 16788 5880 16848 5890
rect 17178 5930 17238 5940
rect 17178 5890 17188 5930
rect 17188 5890 17228 5930
rect 17228 5890 17238 5930
rect 17178 5880 17238 5890
rect 18008 6380 18068 6390
rect 18008 6340 18018 6380
rect 18018 6340 18058 6380
rect 18058 6340 18068 6380
rect 18008 6330 18068 6340
rect 18298 6330 18358 6390
rect 18408 7100 18468 7160
rect 20328 12780 20388 12790
rect 20328 12740 20338 12780
rect 20338 12740 20378 12780
rect 20378 12740 20388 12780
rect 20328 12730 20388 12740
rect 19528 11930 19588 11990
rect 19728 11930 19788 11990
rect 19928 12070 19988 12130
rect 20728 12780 20788 12790
rect 20728 12740 20738 12780
rect 20738 12740 20778 12780
rect 20778 12740 20788 12780
rect 20728 12730 20788 12740
rect 20128 11930 20188 11990
rect 20528 11930 20588 11990
rect 21128 12070 21188 12130
rect 20928 11930 20988 11990
rect 21008 11980 21068 11990
rect 21008 11940 21018 11980
rect 21018 11940 21058 11980
rect 21058 11940 21068 11980
rect 21008 11930 21068 11940
rect 21328 11930 21388 11990
rect 21528 11930 21588 11990
rect 22128 11980 22188 11990
rect 22128 11940 22138 11980
rect 22138 11940 22178 11980
rect 22178 11940 22188 11980
rect 22128 11930 22188 11940
rect 19928 11870 19988 11880
rect 19928 11830 19938 11870
rect 19938 11830 19978 11870
rect 19978 11830 19988 11870
rect 19928 11820 19988 11830
rect 19628 11490 19688 11500
rect 19628 11450 19638 11490
rect 19638 11450 19678 11490
rect 19678 11450 19688 11490
rect 19628 11440 19688 11450
rect 20068 11490 20128 11500
rect 20068 11450 20078 11490
rect 20078 11450 20118 11490
rect 20118 11450 20128 11490
rect 20068 11440 20128 11450
rect 19978 11270 20038 11330
rect 21138 11420 21198 11480
rect 21908 11490 21968 11500
rect 21908 11450 21918 11490
rect 21918 11450 21958 11490
rect 21958 11450 21968 11490
rect 21908 11440 21968 11450
rect 22748 11490 22808 11500
rect 22748 11450 22758 11490
rect 22758 11450 22798 11490
rect 22798 11450 22808 11490
rect 22748 11440 22808 11450
rect 23228 11440 23288 11500
rect 23458 11510 23528 11580
rect 20728 11350 20788 11410
rect 20068 11170 20128 11230
rect 20768 11150 20828 11160
rect 20768 11110 20778 11150
rect 20778 11110 20818 11150
rect 20818 11110 20828 11150
rect 20768 11100 20828 11110
rect 21908 11270 21968 11280
rect 21908 11230 21918 11270
rect 21918 11230 21958 11270
rect 21958 11230 21968 11270
rect 21908 11220 21968 11230
rect 23618 11320 23678 11330
rect 23618 11280 23628 11320
rect 23628 11280 23668 11320
rect 23668 11280 23678 11320
rect 23618 11270 23678 11280
rect 25898 11270 25958 11330
rect 21208 11150 21268 11160
rect 21208 11110 21218 11150
rect 21218 11110 21258 11150
rect 21258 11110 21268 11150
rect 21208 11100 21268 11110
rect 22748 11150 22808 11160
rect 22748 11110 22758 11150
rect 22758 11110 22798 11150
rect 22798 11110 22808 11150
rect 22748 11100 22808 11110
rect 23228 11100 23288 11160
rect 20988 10870 21048 10880
rect 20988 10830 20998 10870
rect 20998 10830 21038 10870
rect 21038 10830 21048 10870
rect 20988 10820 21048 10830
rect 19408 10710 19468 10770
rect 19608 10710 19668 10770
rect 19848 10760 19908 10770
rect 19848 10720 19858 10760
rect 19858 10720 19898 10760
rect 19898 10720 19908 10760
rect 19848 10710 19908 10720
rect 20008 10710 20068 10770
rect 20408 10710 20468 10770
rect 20808 10710 20868 10770
rect 20988 10650 21048 10660
rect 20988 10610 20998 10650
rect 20998 10610 21038 10650
rect 21038 10610 21048 10650
rect 20988 10600 21048 10610
rect 21208 10710 21268 10770
rect 21408 10710 21468 10770
rect 22128 10760 22188 10770
rect 22128 10720 22138 10760
rect 22138 10720 22178 10760
rect 22178 10720 22188 10760
rect 22128 10710 22188 10720
rect 23458 11000 23528 11070
rect 23018 9640 23078 9650
rect 23018 9600 23028 9640
rect 23028 9600 23068 9640
rect 23068 9600 23078 9640
rect 23018 9590 23078 9600
rect 23228 9070 23288 9130
rect 19038 8710 19098 8770
rect 19038 8630 19098 8690
rect 19038 8550 19098 8610
rect 19148 8440 19208 8500
rect 25898 8440 25958 8500
rect 26008 8710 26068 8770
rect 26088 8710 26148 8770
rect 26168 8710 26228 8770
rect 26248 8710 26308 8770
rect 26328 8710 26388 8770
rect 26408 8710 26468 8770
rect 26008 8630 26068 8690
rect 26088 8630 26148 8690
rect 26168 8630 26228 8690
rect 26248 8630 26308 8690
rect 26328 8630 26388 8690
rect 26408 8630 26468 8690
rect 26008 8550 26068 8610
rect 26088 8550 26148 8610
rect 26168 8550 26228 8610
rect 26248 8550 26308 8610
rect 26328 8550 26388 8610
rect 26408 8550 26468 8610
rect 23108 8310 23178 8380
rect 19348 8170 19408 8230
rect 19568 8170 19628 8230
rect 20008 8170 20068 8230
rect 20328 8170 20388 8230
rect 20648 8170 20708 8230
rect 21088 8170 21148 8230
rect 19788 7320 19848 7380
rect 19148 7100 19208 7160
rect 20208 7100 20268 7160
rect 18928 6980 18988 7040
rect 19988 6980 20048 7040
rect 19548 6330 19608 6390
rect 20428 6980 20488 7040
rect 19768 6330 19828 6390
rect 21408 8170 21468 8230
rect 21728 8170 21788 8230
rect 22168 8170 22228 8230
rect 21818 7560 21878 7570
rect 21818 7520 21828 7560
rect 21828 7520 21868 7560
rect 21868 7520 21878 7560
rect 21818 7510 21878 7520
rect 22388 8170 22448 8230
rect 22078 7560 22138 7570
rect 22078 7520 22088 7560
rect 22088 7520 22128 7560
rect 22128 7520 22138 7560
rect 22078 7510 22138 7520
rect 22758 7520 22828 7590
rect 20868 6980 20928 7040
rect 21378 7210 21438 7270
rect 21378 7060 21438 7070
rect 21378 7020 21388 7060
rect 21388 7020 21428 7060
rect 21428 7020 21438 7060
rect 21378 7010 21438 7020
rect 21948 7260 22008 7320
rect 21508 6980 21568 7040
rect 20208 6330 20268 6390
rect 20648 6330 20708 6390
rect 20968 6330 21028 6390
rect 26008 7260 26068 7320
rect 26088 7260 26148 7320
rect 26168 7260 26228 7320
rect 26248 7260 26308 7320
rect 26328 7260 26388 7320
rect 26408 7260 26468 7320
rect 21948 6980 22008 7040
rect 22078 7060 22138 7070
rect 22078 7020 22088 7060
rect 22088 7020 22128 7060
rect 22128 7020 22138 7060
rect 22078 7010 22138 7020
rect 21288 6330 21348 6390
rect 22758 6990 22828 7060
rect 21728 6330 21788 6390
rect 22168 6330 22228 6390
rect 22388 6330 22448 6390
rect 18408 5990 18468 6050
rect 17698 5820 17758 5880
rect 22998 5810 23068 5880
rect 23588 5580 23648 5640
rect 24108 5580 24168 5640
rect 24628 5580 24688 5640
rect 25148 5580 25208 5640
rect 23398 4980 23458 4990
rect 23398 4940 23408 4980
rect 23408 4940 23448 4980
rect 23448 4940 23458 4980
rect 23398 4930 23458 4940
rect 23318 4750 23378 4810
rect 23588 4750 23648 4810
rect 23918 4980 23978 4990
rect 23918 4940 23928 4980
rect 23928 4940 23968 4980
rect 23968 4940 23978 4980
rect 23918 4930 23978 4940
rect 23838 4750 23898 4810
rect 24108 4750 24168 4810
rect 23318 4210 23378 4220
rect 23318 4170 23328 4210
rect 23328 4170 23368 4210
rect 23368 4170 23378 4210
rect 23318 4160 23378 4170
rect 23418 4160 23478 4220
rect 23282 4092 23334 4100
rect 23282 4058 23290 4092
rect 23290 4058 23324 4092
rect 23324 4058 23334 4092
rect 23282 4048 23334 4058
rect 12708 3730 12768 3740
rect 12708 3690 12718 3730
rect 12718 3690 12758 3730
rect 12758 3690 12768 3730
rect 12708 3680 12768 3690
rect 13128 3730 13188 3740
rect 13128 3690 13138 3730
rect 13138 3690 13178 3730
rect 13178 3690 13188 3730
rect 13128 3680 13188 3690
rect 13798 3730 13858 3740
rect 13798 3690 13808 3730
rect 13808 3690 13848 3730
rect 13848 3690 13858 3730
rect 13798 3680 13858 3690
rect 14368 3730 14428 3740
rect 14368 3690 14378 3730
rect 14378 3690 14418 3730
rect 14418 3690 14428 3730
rect 14368 3680 14428 3690
rect 15078 3730 15138 3740
rect 15078 3690 15088 3730
rect 15088 3690 15128 3730
rect 15128 3690 15138 3730
rect 15078 3680 15138 3690
rect 15508 3730 15568 3740
rect 15508 3690 15518 3730
rect 15518 3690 15558 3730
rect 15558 3690 15568 3730
rect 15508 3680 15568 3690
rect 15948 3730 16008 3740
rect 15948 3690 15958 3730
rect 15958 3690 15998 3730
rect 15998 3690 16008 3730
rect 15948 3680 16008 3690
rect 16198 3730 16258 3740
rect 16198 3690 16208 3730
rect 16208 3690 16248 3730
rect 16248 3690 16258 3730
rect 16198 3680 16258 3690
rect 16418 3730 16478 3740
rect 16418 3690 16428 3730
rect 16428 3690 16468 3730
rect 16468 3690 16478 3730
rect 16418 3680 16478 3690
rect 16888 3730 16948 3740
rect 16888 3690 16898 3730
rect 16898 3690 16938 3730
rect 16938 3690 16948 3730
rect 16888 3680 16948 3690
rect 17328 3730 17388 3740
rect 17328 3690 17338 3730
rect 17338 3690 17378 3730
rect 17378 3690 17388 3730
rect 17328 3680 17388 3690
rect 17948 3730 18008 3740
rect 17948 3690 17958 3730
rect 17958 3690 17998 3730
rect 17998 3690 18008 3730
rect 17948 3680 18008 3690
rect 18288 3730 18348 3740
rect 18288 3690 18298 3730
rect 18298 3690 18338 3730
rect 18338 3690 18348 3730
rect 18288 3680 18348 3690
rect 18648 3730 18708 3740
rect 18648 3690 18658 3730
rect 18658 3690 18698 3730
rect 18698 3690 18708 3730
rect 18648 3680 18708 3690
rect 19248 3730 19308 3740
rect 19248 3690 19258 3730
rect 19258 3690 19298 3730
rect 19298 3690 19308 3730
rect 19248 3680 19308 3690
rect 19588 3730 19648 3740
rect 19588 3690 19598 3730
rect 19598 3690 19638 3730
rect 19638 3690 19648 3730
rect 19588 3680 19648 3690
rect 19948 3730 20008 3740
rect 19948 3690 19958 3730
rect 19958 3690 19998 3730
rect 19998 3690 20008 3730
rect 19948 3680 20008 3690
rect 20548 3730 20608 3740
rect 20548 3690 20558 3730
rect 20558 3690 20598 3730
rect 20598 3690 20608 3730
rect 20548 3680 20608 3690
rect 20888 3730 20948 3740
rect 20888 3690 20898 3730
rect 20898 3690 20938 3730
rect 20938 3690 20948 3730
rect 20888 3680 20948 3690
rect 21248 3730 21308 3740
rect 21248 3690 21258 3730
rect 21258 3690 21298 3730
rect 21298 3690 21308 3730
rect 21248 3680 21308 3690
rect 21848 3730 21908 3740
rect 21848 3690 21858 3730
rect 21858 3690 21898 3730
rect 21898 3690 21908 3730
rect 21848 3680 21908 3690
rect 22188 3730 22248 3740
rect 22188 3690 22198 3730
rect 22198 3690 22238 3730
rect 22238 3690 22248 3730
rect 22188 3680 22248 3690
rect 22548 3730 22608 3740
rect 22548 3690 22558 3730
rect 22558 3690 22598 3730
rect 22598 3690 22608 3730
rect 22548 3680 22608 3690
rect 22818 3350 22878 3410
rect 22898 3350 22958 3410
rect 22978 3350 23038 3410
rect 12118 3280 12178 3340
rect 12328 3330 12388 3340
rect 12328 3290 12338 3330
rect 12338 3290 12378 3330
rect 12378 3290 12388 3330
rect 12328 3280 12388 3290
rect 22754 3322 22806 3330
rect 22754 3288 22762 3322
rect 22762 3288 22796 3322
rect 22796 3288 22806 3322
rect 22754 3278 22806 3288
rect 22818 3270 22878 3330
rect 22898 3270 22958 3330
rect 22978 3270 23038 3330
rect 22818 3190 22878 3250
rect 22898 3190 22958 3250
rect 22978 3190 23038 3250
rect 12548 2950 12608 2960
rect 12548 2910 12558 2950
rect 12558 2910 12598 2950
rect 12598 2910 12608 2950
rect 12548 2900 12608 2910
rect 12768 2950 12828 2960
rect 12768 2910 12778 2950
rect 12778 2910 12818 2950
rect 12818 2910 12828 2950
rect 12768 2900 12828 2910
rect 13238 2950 13298 2960
rect 13238 2910 13248 2950
rect 13248 2910 13288 2950
rect 13288 2910 13298 2950
rect 13238 2900 13298 2910
rect 13578 2950 13638 2960
rect 13578 2910 13588 2950
rect 13588 2910 13628 2950
rect 13628 2910 13638 2950
rect 13578 2900 13638 2910
rect 13798 2950 13858 2960
rect 13798 2910 13808 2950
rect 13808 2910 13848 2950
rect 13848 2910 13858 2950
rect 13798 2900 13858 2910
rect 14238 2950 14298 2960
rect 14238 2910 14248 2950
rect 14248 2910 14288 2950
rect 14288 2910 14298 2950
rect 14238 2900 14298 2910
rect 14918 2950 14978 2960
rect 14918 2910 14928 2950
rect 14928 2910 14968 2950
rect 14968 2910 14978 2950
rect 14918 2900 14978 2910
rect 15138 2950 15198 2960
rect 15138 2910 15148 2950
rect 15148 2910 15188 2950
rect 15188 2910 15198 2950
rect 15138 2900 15198 2910
rect 15608 2950 15668 2960
rect 15608 2910 15618 2950
rect 15618 2910 15658 2950
rect 15658 2910 15668 2950
rect 15608 2900 15668 2910
rect 16068 2950 16128 2960
rect 16068 2910 16078 2950
rect 16078 2910 16118 2950
rect 16118 2910 16128 2950
rect 16068 2900 16128 2910
rect 16418 2950 16478 2960
rect 16418 2910 16428 2950
rect 16428 2910 16468 2950
rect 16468 2910 16478 2950
rect 16418 2900 16478 2910
rect 16668 2950 16728 2960
rect 16668 2910 16678 2950
rect 16678 2910 16718 2950
rect 16718 2910 16728 2950
rect 16668 2900 16728 2910
rect 16888 2950 16948 2960
rect 16888 2910 16898 2950
rect 16898 2910 16938 2950
rect 16938 2910 16948 2950
rect 16888 2900 16948 2910
rect 17218 2950 17278 2960
rect 17218 2910 17228 2950
rect 17228 2910 17268 2950
rect 17268 2910 17278 2950
rect 17218 2900 17278 2910
rect 17878 2950 17938 2960
rect 17878 2910 17888 2950
rect 17888 2910 17928 2950
rect 17928 2910 17938 2950
rect 17878 2900 17938 2910
rect 18098 2950 18158 2960
rect 18098 2910 18108 2950
rect 18108 2910 18148 2950
rect 18148 2910 18158 2950
rect 18098 2900 18158 2910
rect 18668 2950 18728 2960
rect 18668 2910 18678 2950
rect 18678 2910 18718 2950
rect 18718 2910 18728 2950
rect 18668 2900 18728 2910
rect 18928 2950 18988 2960
rect 18928 2910 18938 2950
rect 18938 2910 18978 2950
rect 18978 2910 18988 2950
rect 18928 2900 18988 2910
rect 19178 2950 19238 2960
rect 19178 2910 19188 2950
rect 19188 2910 19228 2950
rect 19228 2910 19238 2950
rect 19178 2900 19238 2910
rect 19398 2950 19458 2960
rect 19398 2910 19408 2950
rect 19408 2910 19448 2950
rect 19448 2910 19458 2950
rect 19398 2900 19458 2910
rect 19948 2950 20008 2960
rect 19948 2910 19958 2950
rect 19958 2910 19998 2950
rect 19998 2910 20008 2950
rect 19948 2900 20008 2910
rect 20228 2950 20288 2960
rect 20228 2910 20238 2950
rect 20238 2910 20278 2950
rect 20278 2910 20288 2950
rect 20228 2900 20288 2910
rect 20478 2950 20538 2960
rect 20478 2910 20488 2950
rect 20488 2910 20528 2950
rect 20528 2910 20538 2950
rect 20478 2900 20538 2910
rect 20698 2950 20758 2960
rect 20698 2910 20708 2950
rect 20708 2910 20748 2950
rect 20748 2910 20758 2950
rect 20698 2900 20758 2910
rect 21248 2950 21308 2960
rect 21248 2910 21258 2950
rect 21258 2910 21298 2950
rect 21298 2910 21308 2950
rect 21248 2900 21308 2910
rect 21528 2950 21588 2960
rect 21528 2910 21538 2950
rect 21538 2910 21578 2950
rect 21578 2910 21588 2950
rect 21528 2900 21588 2910
rect 21778 2950 21838 2960
rect 21778 2910 21788 2950
rect 21788 2910 21828 2950
rect 21828 2910 21838 2950
rect 21778 2900 21838 2910
rect 21998 2950 22058 2960
rect 21998 2910 22008 2950
rect 22008 2910 22048 2950
rect 22048 2910 22058 2950
rect 21998 2900 22058 2910
rect 22548 2950 22608 2960
rect 22548 2910 22558 2950
rect 22558 2910 22598 2950
rect 22598 2910 22608 2950
rect 22548 2900 22608 2910
rect 23248 3350 23308 3410
rect 23248 3270 23308 3330
rect 23248 3190 23308 3250
rect 23338 3350 23398 3410
rect 23338 3270 23398 3330
rect 23338 3190 23398 3250
rect 24438 4980 24498 4990
rect 24438 4940 24448 4980
rect 24448 4940 24488 4980
rect 24488 4940 24498 4980
rect 24438 4930 24498 4940
rect 24768 4930 24828 4990
rect 24958 4980 25018 4990
rect 24958 4940 24968 4980
rect 24968 4940 25008 4980
rect 25008 4940 25018 4980
rect 24958 4930 25018 4940
rect 24358 4750 24418 4810
rect 24628 4750 24688 4810
rect 23838 4210 23898 4220
rect 23838 4170 23848 4210
rect 23848 4170 23888 4210
rect 23888 4170 23898 4210
rect 23838 4160 23898 4170
rect 23938 4160 23998 4220
rect 23282 2742 23334 2750
rect 23282 2708 23290 2742
rect 23290 2708 23324 2742
rect 23324 2708 23334 2742
rect 23282 2698 23334 2708
rect 23418 2700 23478 2760
rect 23528 4040 23588 4100
rect 23318 2630 23378 2640
rect 23318 2590 23328 2630
rect 23328 2590 23368 2630
rect 23368 2590 23378 2630
rect 23318 2580 23378 2590
rect 23802 4092 23854 4100
rect 23802 4058 23810 4092
rect 23810 4058 23844 4092
rect 23844 4058 23854 4092
rect 23802 4048 23854 4058
rect 23768 3350 23828 3410
rect 23768 3270 23828 3330
rect 23768 3190 23828 3250
rect 23858 3350 23918 3410
rect 23858 3270 23918 3330
rect 23858 3190 23918 3250
rect 23528 2580 23588 2640
rect 24358 4210 24418 4220
rect 24358 4170 24368 4210
rect 24368 4170 24408 4210
rect 24408 4170 24418 4210
rect 24358 4160 24418 4170
rect 24458 4160 24518 4220
rect 23802 2742 23854 2750
rect 23802 2708 23810 2742
rect 23810 2708 23844 2742
rect 23844 2708 23854 2742
rect 23802 2698 23854 2708
rect 23938 2700 23998 2760
rect 24048 4040 24108 4100
rect 23268 2262 23320 2270
rect 23268 2228 23276 2262
rect 23276 2228 23310 2262
rect 23310 2228 23320 2262
rect 23268 2218 23320 2228
rect 23838 2630 23898 2640
rect 23838 2590 23848 2630
rect 23848 2590 23888 2630
rect 23888 2590 23898 2630
rect 23838 2580 23898 2590
rect 24322 4092 24374 4100
rect 24322 4058 24330 4092
rect 24330 4058 24364 4092
rect 24364 4058 24374 4092
rect 24322 4048 24374 4058
rect 24288 3350 24348 3410
rect 24288 3270 24348 3330
rect 24288 3190 24348 3250
rect 24378 3350 24438 3410
rect 24378 3270 24438 3330
rect 24378 3190 24438 3250
rect 24048 2580 24108 2640
rect 24322 2742 24374 2750
rect 24322 2708 24330 2742
rect 24330 2708 24364 2742
rect 24364 2708 24374 2742
rect 24322 2698 24374 2708
rect 24458 2700 24518 2760
rect 24568 4040 24628 4100
rect 23788 2262 23840 2270
rect 23788 2228 23796 2262
rect 23796 2228 23830 2262
rect 23830 2228 23840 2262
rect 23788 2218 23840 2228
rect 24358 2630 24418 2640
rect 24358 2590 24368 2630
rect 24368 2590 24408 2630
rect 24408 2590 24418 2630
rect 24358 2580 24418 2590
rect 24568 2580 24628 2640
rect 24308 2262 24360 2270
rect 24308 2228 24316 2262
rect 24316 2228 24350 2262
rect 24350 2228 24360 2262
rect 24308 2218 24360 2228
rect 24874 2262 24926 2270
rect 24874 2228 24884 2262
rect 24884 2228 24918 2262
rect 24918 2228 24926 2262
rect 24874 2218 24926 2228
rect 25178 3350 25238 3410
rect 25258 3350 25318 3410
rect 25338 3350 25398 3410
rect 25178 3270 25238 3330
rect 25258 3270 25318 3330
rect 25338 3270 25398 3330
rect 25178 3190 25238 3250
rect 25258 3190 25318 3250
rect 25338 3190 25398 3250
rect 22818 1770 22878 1830
rect 22898 1770 22958 1830
rect 22978 1770 23038 1830
rect 22818 1690 22878 1750
rect 22898 1690 22958 1750
rect 22978 1690 23038 1750
rect 22818 1610 22878 1670
rect 22898 1610 22958 1670
rect 22978 1610 23038 1670
rect 23318 1500 23378 1560
rect 23838 1500 23898 1560
rect 24358 1500 24418 1560
rect 26008 2220 26068 2280
rect 26088 2220 26148 2280
rect 26168 2220 26228 2280
rect 26248 2220 26308 2280
rect 26328 2220 26388 2280
rect 26408 2220 26468 2280
rect 25178 1770 25238 1830
rect 25258 1770 25318 1830
rect 25338 1770 25398 1830
rect 25178 1690 25238 1750
rect 25258 1690 25318 1750
rect 25338 1690 25398 1750
rect 25178 1610 25238 1670
rect 25258 1610 25318 1670
rect 25338 1610 25398 1670
rect 24848 1500 24908 1560
rect 11948 1270 12008 1330
<< metal2 >>
rect 7458 19880 7718 19890
rect 7458 19820 7468 19880
rect 7528 19820 7558 19880
rect 7618 19820 7648 19880
rect 7708 19820 7718 19880
rect 7458 19810 7718 19820
rect 7458 19790 23408 19810
rect 7458 19730 7468 19790
rect 7528 19730 7558 19790
rect 7618 19730 7648 19790
rect 7708 19730 22818 19790
rect 7458 19720 22818 19730
rect 22888 19720 23318 19790
rect 23388 19720 23408 19790
rect 7458 19700 23408 19720
rect 7458 19640 7468 19700
rect 7528 19640 7558 19700
rect 7618 19640 7648 19700
rect 7708 19640 7718 19700
rect 7458 19630 7718 19640
rect 16118 19690 16198 19700
rect 16118 19630 16128 19690
rect 16188 19630 16198 19690
rect 16118 19620 16198 19630
rect 8918 19510 9018 19520
rect 25988 19510 26088 19520
rect 8918 19500 15418 19510
rect 8918 19440 8938 19500
rect 8998 19440 14998 19500
rect 15408 19440 15418 19500
rect 8918 19430 15418 19440
rect 16898 19500 26478 19510
rect 16898 19440 16908 19500
rect 17318 19440 26008 19500
rect 26068 19440 26098 19500
rect 26158 19440 26198 19500
rect 26258 19440 26308 19500
rect 26368 19440 26408 19500
rect 26468 19440 26478 19500
rect 16898 19430 26478 19440
rect 8918 19420 9018 19430
rect 25988 19420 26088 19430
rect 8868 19190 18268 19200
rect 8868 19130 8878 19190
rect 8938 19130 18198 19190
rect 18258 19130 18268 19190
rect 8868 19120 18268 19130
rect 7458 19080 17648 19090
rect 7458 19050 8458 19080
rect 7458 18990 7468 19050
rect 7528 18990 7558 19050
rect 7618 18990 7648 19050
rect 7708 19020 8458 19050
rect 8518 19020 9248 19080
rect 9308 19020 10688 19080
rect 10748 19020 13248 19080
rect 13308 19020 15678 19080
rect 15738 19020 16788 19080
rect 16848 19020 17578 19080
rect 17638 19020 17648 19080
rect 7708 19000 17648 19020
rect 7708 18990 8458 19000
rect 7458 18950 8458 18990
rect 7458 18890 7468 18950
rect 7528 18890 7558 18950
rect 7618 18890 7648 18950
rect 7708 18940 8458 18950
rect 8518 18940 9248 19000
rect 9308 18940 10688 19000
rect 10748 18940 13248 19000
rect 13308 18940 15678 19000
rect 15738 18940 16788 19000
rect 16848 18940 17578 19000
rect 17638 18940 17648 19000
rect 7708 18920 17648 18940
rect 7708 18890 8458 18920
rect 7458 18860 8458 18890
rect 8518 18860 9248 18920
rect 9308 18860 10688 18920
rect 10748 18860 13248 18920
rect 13308 18860 15678 18920
rect 15738 18860 16788 18920
rect 16848 18860 17578 18920
rect 17638 18860 17648 18920
rect 7458 18850 17648 18860
rect 18188 18850 18268 18860
rect 18188 18790 18198 18850
rect 18258 18790 18268 18850
rect 18188 18780 18268 18790
rect 8448 18450 8948 18460
rect 8448 18440 8878 18450
rect 8448 18040 8458 18440
rect 8518 18390 8878 18440
rect 8938 18390 8948 18450
rect 8518 18370 8948 18390
rect 8518 18310 8878 18370
rect 8938 18310 8948 18370
rect 8518 18280 8948 18310
rect 8518 18220 8878 18280
rect 8938 18220 8948 18280
rect 8518 18190 8948 18220
rect 8518 18130 8878 18190
rect 8938 18130 8948 18190
rect 8518 18110 8948 18130
rect 8518 18050 8878 18110
rect 8938 18050 8948 18110
rect 8518 18040 8948 18050
rect 8448 18030 8948 18040
rect 17568 18450 18028 18460
rect 17568 18440 17958 18450
rect 17568 18040 17578 18440
rect 17638 18390 17958 18440
rect 18018 18390 18028 18450
rect 17638 18370 18028 18390
rect 17638 18310 17958 18370
rect 18018 18310 18028 18370
rect 17638 18280 18028 18310
rect 17638 18220 17958 18280
rect 18018 18220 18028 18280
rect 17638 18190 18028 18220
rect 17638 18130 17958 18190
rect 18018 18130 18028 18190
rect 17638 18110 18028 18130
rect 17638 18050 17958 18110
rect 18018 18050 18028 18110
rect 18638 18150 18738 18170
rect 18638 18090 18658 18150
rect 18718 18090 18738 18150
rect 18638 18070 18738 18090
rect 17638 18040 18028 18050
rect 17568 18030 18028 18040
rect 18118 17450 18198 17460
rect 18118 17390 18128 17450
rect 18188 17390 18198 17450
rect 18118 17380 18198 17390
rect 11138 16810 11648 16820
rect 11138 16750 11148 16810
rect 11208 16750 11578 16810
rect 11638 16750 11648 16810
rect 11138 16740 11648 16750
rect 13238 16810 15418 16820
rect 13238 16750 13248 16810
rect 13308 16750 15348 16810
rect 15408 16750 15418 16810
rect 13238 16740 15418 16750
rect 17568 16750 18878 16770
rect 17568 16690 17578 16750
rect 17638 16690 18798 16750
rect 18858 16690 18878 16750
rect 17568 16670 18878 16690
rect 17948 16050 19068 16060
rect 17948 15990 17958 16050
rect 18018 15990 18998 16050
rect 19058 15990 19068 16050
rect 17948 15980 19068 15990
rect 16348 15350 18878 15370
rect 16348 15290 16358 15350
rect 16418 15290 16438 15350
rect 16498 15290 16518 15350
rect 16578 15290 18798 15350
rect 18858 15290 18878 15350
rect 16348 15270 18878 15290
rect 15338 14800 16318 14810
rect 15338 14740 15348 14800
rect 15408 14740 16008 14800
rect 16068 14740 16248 14800
rect 16308 14740 16318 14800
rect 15338 14730 16318 14740
rect 10348 14720 14028 14730
rect 10348 14660 10358 14720
rect 10418 14660 13958 14720
rect 14018 14660 14028 14720
rect 10348 14650 14028 14660
rect 11138 14610 12548 14620
rect 11138 14550 11148 14610
rect 11208 14550 12550 14610
rect 11138 14540 12550 14550
rect 12620 14540 12630 14610
rect 13938 14540 13948 14610
rect 14018 14590 14028 14610
rect 16148 14600 16228 14610
rect 16148 14590 16158 14600
rect 14018 14550 16158 14590
rect 14018 14540 14028 14550
rect 16148 14540 16158 14550
rect 16218 14540 16228 14600
rect 16148 14530 16228 14540
rect 9678 14490 16858 14500
rect 9678 14430 9688 14490
rect 9748 14430 16788 14490
rect 16848 14430 16858 14490
rect 9678 14420 16858 14430
rect 10618 14380 18728 14390
rect 10618 14320 10628 14380
rect 10688 14320 11038 14380
rect 11098 14320 18658 14380
rect 18718 14320 18728 14380
rect 10618 14310 18728 14320
rect 15468 14250 18578 14260
rect 9458 14210 11158 14220
rect 9458 14150 9468 14210
rect 9528 14150 11088 14210
rect 11148 14150 11158 14210
rect 9458 14140 11158 14150
rect 15468 14190 15478 14250
rect 15538 14210 18578 14250
rect 15538 14190 18378 14210
rect 15468 14170 18378 14190
rect 15468 14110 15478 14170
rect 15538 14150 18378 14170
rect 18438 14150 18478 14210
rect 18538 14150 18578 14210
rect 15538 14110 18578 14150
rect 15468 14100 18578 14110
rect 11158 14040 11238 14050
rect 11158 13980 11168 14040
rect 11228 14030 11238 14040
rect 11318 14040 11398 14050
rect 11318 14030 11328 14040
rect 11228 13990 11328 14030
rect 11228 13980 11238 13990
rect 11158 13970 11238 13980
rect 11318 13980 11328 13990
rect 11388 14030 11398 14040
rect 11478 14040 11558 14050
rect 11478 14030 11488 14040
rect 11388 13990 11488 14030
rect 11388 13980 11398 13990
rect 11318 13970 11398 13980
rect 11478 13980 11488 13990
rect 11548 14030 11558 14040
rect 11638 14040 11718 14050
rect 11638 14030 11648 14040
rect 11548 13990 11648 14030
rect 11548 13980 11558 13990
rect 11478 13970 11558 13980
rect 11638 13980 11648 13990
rect 11708 14030 11718 14040
rect 11798 14040 11878 14050
rect 11798 14030 11808 14040
rect 11708 13990 11808 14030
rect 11708 13980 11718 13990
rect 11638 13970 11718 13980
rect 11798 13980 11808 13990
rect 11868 14030 11878 14040
rect 11958 14040 12038 14050
rect 11958 14030 11968 14040
rect 11868 13990 11968 14030
rect 11868 13980 11878 13990
rect 11798 13970 11878 13980
rect 11958 13980 11968 13990
rect 12028 14030 12038 14040
rect 12118 14040 12198 14050
rect 12118 14030 12128 14040
rect 12028 13990 12128 14030
rect 12028 13980 12038 13990
rect 11958 13970 12038 13980
rect 12118 13980 12128 13990
rect 12188 14030 12198 14040
rect 12278 14040 12358 14050
rect 12278 14030 12288 14040
rect 12188 13990 12288 14030
rect 12188 13980 12198 13990
rect 12118 13970 12198 13980
rect 12278 13980 12288 13990
rect 12348 14030 12358 14040
rect 12438 14040 12518 14050
rect 12438 14030 12448 14040
rect 12348 13990 12448 14030
rect 12348 13980 12358 13990
rect 12278 13970 12358 13980
rect 12438 13980 12448 13990
rect 12508 14030 12518 14040
rect 12598 14040 12678 14050
rect 12598 14030 12608 14040
rect 12508 13990 12608 14030
rect 12508 13980 12518 13990
rect 12438 13970 12518 13980
rect 12598 13980 12608 13990
rect 12668 14030 12678 14040
rect 12758 14040 12838 14050
rect 12758 14030 12768 14040
rect 12668 13990 12768 14030
rect 12668 13980 12678 13990
rect 12598 13970 12678 13980
rect 12758 13980 12768 13990
rect 12828 14030 12838 14040
rect 12918 14040 12998 14050
rect 12918 14030 12928 14040
rect 12828 13990 12928 14030
rect 12828 13980 12838 13990
rect 12758 13970 12838 13980
rect 12918 13980 12928 13990
rect 12988 14030 12998 14040
rect 13078 14040 13158 14050
rect 13078 14030 13088 14040
rect 12988 13990 13088 14030
rect 12988 13980 12998 13990
rect 12918 13970 12998 13980
rect 13078 13980 13088 13990
rect 13148 13980 13158 14040
rect 13078 13970 13158 13980
rect 13238 14040 13318 14050
rect 13238 13980 13248 14040
rect 13308 14030 13318 14040
rect 13398 14040 13478 14050
rect 13398 14030 13408 14040
rect 13308 13990 13408 14030
rect 13308 13980 13318 13990
rect 13238 13970 13318 13980
rect 13398 13980 13408 13990
rect 13468 14030 13478 14040
rect 13558 14040 13638 14050
rect 13558 14030 13568 14040
rect 13468 13990 13568 14030
rect 13468 13980 13478 13990
rect 13398 13970 13478 13980
rect 13558 13980 13568 13990
rect 13628 14030 13638 14040
rect 13718 14040 13798 14050
rect 13718 14030 13728 14040
rect 13628 13990 13728 14030
rect 13628 13980 13638 13990
rect 13558 13970 13638 13980
rect 13718 13980 13728 13990
rect 13788 14030 13798 14040
rect 13878 14040 13958 14050
rect 13878 14030 13888 14040
rect 13788 13990 13888 14030
rect 13788 13980 13798 13990
rect 13718 13970 13798 13980
rect 13878 13980 13888 13990
rect 13948 14030 13958 14040
rect 14038 14040 14118 14050
rect 14038 14030 14048 14040
rect 13948 13990 14048 14030
rect 13948 13980 13958 13990
rect 13878 13970 13958 13980
rect 14038 13980 14048 13990
rect 14108 14030 14118 14040
rect 14198 14040 14278 14050
rect 14198 14030 14208 14040
rect 14108 13990 14208 14030
rect 14108 13980 14118 13990
rect 14038 13970 14118 13980
rect 14198 13980 14208 13990
rect 14268 14030 14278 14040
rect 14358 14040 14438 14050
rect 14358 14030 14368 14040
rect 14268 13990 14368 14030
rect 14268 13980 14278 13990
rect 14198 13970 14278 13980
rect 14358 13980 14368 13990
rect 14428 14030 14438 14040
rect 14518 14040 14598 14050
rect 14518 14030 14528 14040
rect 14428 13990 14528 14030
rect 14428 13980 14438 13990
rect 14358 13970 14438 13980
rect 14518 13980 14528 13990
rect 14588 14030 14598 14040
rect 14678 14040 14758 14050
rect 14678 14030 14688 14040
rect 14588 13990 14688 14030
rect 14588 13980 14598 13990
rect 14518 13970 14598 13980
rect 14678 13980 14688 13990
rect 14748 14030 14758 14040
rect 14838 14040 14918 14050
rect 14838 14030 14848 14040
rect 14748 13990 14848 14030
rect 14748 13980 14758 13990
rect 14678 13970 14758 13980
rect 14838 13980 14848 13990
rect 14908 14030 14918 14040
rect 14998 14040 15078 14050
rect 14998 14030 15008 14040
rect 14908 13990 15008 14030
rect 14908 13980 14918 13990
rect 14838 13970 14918 13980
rect 14998 13980 15008 13990
rect 15068 14030 15078 14040
rect 15158 14040 15238 14050
rect 15158 14030 15168 14040
rect 15068 13990 15168 14030
rect 15068 13980 15078 13990
rect 14998 13970 15078 13980
rect 15158 13980 15168 13990
rect 15228 13980 15238 14040
rect 15158 13970 15238 13980
rect 11898 13930 18578 13940
rect 11898 13870 11908 13930
rect 11968 13870 13168 13930
rect 13228 13870 13248 13930
rect 13308 13870 13328 13930
rect 13388 13870 14588 13930
rect 14648 13900 18578 13930
rect 14648 13870 18378 13900
rect 11898 13850 18378 13870
rect 11898 13790 11908 13850
rect 11968 13790 13168 13850
rect 13228 13790 13248 13850
rect 13308 13790 13328 13850
rect 13388 13790 14588 13850
rect 14648 13840 18378 13850
rect 18438 13840 18478 13900
rect 18538 13840 18578 13900
rect 14648 13800 18578 13840
rect 14648 13790 18378 13800
rect 11898 13770 18378 13790
rect 11898 13710 11908 13770
rect 11968 13710 13168 13770
rect 13228 13710 13248 13770
rect 13308 13710 13328 13770
rect 13388 13710 14588 13770
rect 14648 13740 18378 13770
rect 18438 13740 18478 13800
rect 18538 13740 18578 13800
rect 14648 13710 18578 13740
rect 11898 13700 18578 13710
rect 23208 13510 23308 13530
rect 23208 13450 23228 13510
rect 23288 13450 23308 13510
rect 18038 13420 18278 13440
rect 23208 13430 23308 13450
rect 18038 13360 18078 13420
rect 18138 13360 18178 13420
rect 18238 13360 18278 13420
rect 18038 13340 18278 13360
rect 18338 13180 23088 13190
rect 10918 13130 18278 13140
rect 10918 13070 10928 13130
rect 10988 13070 11168 13130
rect 11228 13070 11408 13130
rect 11468 13070 11648 13130
rect 11708 13070 12288 13130
rect 12348 13070 12528 13130
rect 12588 13070 12768 13130
rect 12828 13070 13728 13130
rect 13788 13070 13968 13130
rect 14028 13070 14208 13130
rect 14268 13070 14848 13130
rect 14908 13070 15088 13130
rect 15148 13070 15328 13130
rect 15388 13070 15568 13130
rect 15628 13100 18278 13130
rect 18338 13120 18378 13180
rect 18438 13120 18478 13180
rect 18538 13120 23018 13180
rect 23078 13120 23088 13180
rect 18338 13110 23088 13120
rect 15628 13070 18078 13100
rect 10918 13050 18078 13070
rect 10918 12990 10928 13050
rect 10988 12990 11168 13050
rect 11228 12990 11408 13050
rect 11468 12990 11648 13050
rect 11708 12990 12288 13050
rect 12348 12990 12528 13050
rect 12588 12990 12768 13050
rect 12828 12990 13728 13050
rect 13788 12990 13968 13050
rect 14028 12990 14208 13050
rect 14268 12990 14848 13050
rect 14908 12990 15088 13050
rect 15148 12990 15328 13050
rect 15388 12990 15568 13050
rect 15628 13040 18078 13050
rect 18138 13040 18178 13100
rect 18238 13040 18278 13100
rect 15628 13000 18278 13040
rect 15628 12990 18078 13000
rect 10918 12970 18078 12990
rect 10918 12910 10928 12970
rect 10988 12910 11168 12970
rect 11228 12910 11408 12970
rect 11468 12910 11648 12970
rect 11708 12910 12288 12970
rect 12348 12910 12528 12970
rect 12588 12910 12768 12970
rect 12828 12910 13728 12970
rect 13788 12910 13968 12970
rect 14028 12910 14208 12970
rect 14268 12910 14848 12970
rect 14908 12910 15088 12970
rect 15148 12910 15328 12970
rect 15388 12910 15568 12970
rect 15628 12940 18078 12970
rect 18138 12940 18178 13000
rect 18238 12940 18278 13000
rect 15628 12910 18278 12940
rect 10918 12900 18278 12910
rect 10738 12860 12528 12870
rect 10738 12800 10748 12860
rect 10808 12800 11498 12860
rect 11558 12800 11718 12860
rect 11778 12800 11978 12860
rect 12038 12800 12198 12860
rect 12258 12800 12458 12860
rect 12518 12800 12528 12860
rect 10738 12790 12528 12800
rect 14028 12860 15818 12870
rect 14028 12800 14038 12860
rect 14098 12800 14298 12860
rect 14358 12800 14518 12860
rect 14578 12800 14778 12860
rect 14838 12800 14998 12860
rect 15058 12800 15748 12860
rect 15808 12800 15818 12860
rect 14028 12790 15818 12800
rect 19138 12790 20798 12800
rect 9678 12750 12447 12760
rect 9678 12690 9688 12750
rect 9748 12698 11431 12750
rect 11483 12698 11791 12750
rect 11843 12698 11911 12750
rect 11963 12698 12271 12750
rect 12323 12698 12391 12750
rect 12443 12698 12447 12750
rect 14109 12750 16228 12760
rect 9748 12690 12447 12698
rect 12798 12730 13758 12740
rect 9678 12680 9758 12690
rect 12798 12670 12808 12730
rect 12868 12670 13168 12730
rect 13228 12670 13248 12730
rect 13308 12670 13328 12730
rect 13388 12670 13688 12730
rect 13748 12670 13758 12730
rect 14109 12698 14113 12750
rect 14165 12698 14233 12750
rect 14285 12698 14593 12750
rect 14645 12698 14713 12750
rect 14765 12698 15073 12750
rect 15125 12698 16158 12750
rect 14109 12690 16158 12698
rect 16218 12690 16228 12750
rect 19138 12730 19148 12790
rect 19208 12730 20328 12790
rect 20388 12730 20728 12790
rect 20788 12730 20798 12790
rect 19138 12720 20798 12730
rect 16148 12680 16228 12690
rect 12798 12650 13758 12670
rect 12798 12590 12808 12650
rect 12868 12590 13168 12650
rect 13228 12590 13248 12650
rect 13308 12590 13328 12650
rect 13388 12590 13688 12650
rect 13748 12590 13758 12650
rect 12798 12570 13758 12590
rect 9568 12522 12548 12530
rect 9568 12520 11534 12522
rect 9568 12460 9578 12520
rect 9638 12470 11534 12520
rect 11586 12470 11692 12522
rect 11744 12470 12016 12522
rect 12068 12470 12170 12522
rect 12222 12470 12494 12522
rect 12546 12470 12548 12522
rect 12798 12510 12808 12570
rect 12868 12510 13168 12570
rect 13228 12510 13248 12570
rect 13308 12510 13328 12570
rect 13388 12510 13688 12570
rect 13748 12510 13758 12570
rect 12798 12500 13758 12510
rect 14008 12522 16318 12530
rect 9638 12460 12548 12470
rect 14008 12470 14010 12522
rect 14062 12470 14334 12522
rect 14386 12470 14488 12522
rect 14540 12470 14812 12522
rect 14864 12470 14970 12522
rect 15022 12520 16318 12522
rect 15022 12470 16248 12520
rect 14008 12460 16248 12470
rect 16308 12460 16318 12520
rect 9568 12450 9648 12460
rect 16238 12450 16318 12460
rect 11598 12420 12638 12430
rect 11598 12360 11608 12420
rect 11668 12360 12088 12420
rect 12148 12360 12568 12420
rect 12628 12360 12638 12420
rect 11598 12350 12638 12360
rect 13918 12420 14958 12430
rect 13918 12360 13928 12420
rect 13988 12360 14408 12420
rect 14468 12360 14888 12420
rect 14948 12360 14958 12420
rect 13918 12350 14958 12360
rect 11358 12310 12398 12320
rect 11358 12250 11368 12310
rect 11428 12250 11848 12310
rect 11908 12250 12328 12310
rect 12388 12250 12398 12310
rect 11358 12240 12398 12250
rect 14158 12310 15198 12320
rect 14158 12250 14168 12310
rect 14228 12250 14648 12310
rect 14708 12250 15128 12310
rect 15188 12250 15198 12310
rect 14158 12240 15198 12250
rect 13738 12200 16588 12210
rect 13738 12140 13748 12200
rect 13808 12140 13928 12200
rect 13988 12140 14168 12200
rect 14228 12140 14408 12200
rect 14468 12140 14648 12200
rect 14708 12140 15128 12200
rect 15188 12140 15368 12200
rect 15428 12140 15788 12200
rect 15848 12140 16358 12200
rect 16418 12140 16438 12200
rect 16498 12140 16518 12200
rect 16578 12140 16588 12200
rect 13738 12120 16588 12140
rect 13738 12060 13748 12120
rect 13808 12060 13928 12120
rect 13988 12060 14168 12120
rect 14228 12060 14408 12120
rect 14468 12060 14648 12120
rect 14708 12060 15128 12120
rect 15188 12060 15368 12120
rect 15428 12060 15788 12120
rect 15848 12060 16358 12120
rect 16418 12060 16438 12120
rect 16498 12060 16518 12120
rect 16578 12060 16588 12120
rect 19918 12130 21198 12140
rect 19918 12070 19928 12130
rect 19988 12070 21128 12130
rect 21188 12070 21198 12130
rect 19918 12060 21198 12070
rect 10618 12040 12818 12050
rect 10618 11980 10628 12040
rect 10688 11980 10708 12040
rect 10768 11980 11128 12040
rect 11188 11980 11368 12040
rect 11428 11980 11848 12040
rect 11908 11980 12088 12040
rect 12148 11980 12568 12040
rect 12628 11980 12748 12040
rect 12808 11980 12818 12040
rect 10618 11970 12818 11980
rect 13738 12040 16588 12060
rect 13738 11980 13748 12040
rect 13808 11980 13928 12040
rect 13988 11980 14168 12040
rect 14228 11980 14408 12040
rect 14468 11980 14648 12040
rect 14708 11980 15128 12040
rect 15188 11980 15368 12040
rect 15428 11980 15788 12040
rect 15848 11980 16358 12040
rect 16418 11980 16438 12040
rect 16498 11980 16518 12040
rect 16578 11980 16588 12040
rect 13738 11970 16588 11980
rect 18038 12000 18278 12010
rect 18038 11990 22198 12000
rect 18038 11930 18078 11990
rect 18138 11930 18178 11990
rect 18238 11930 19528 11990
rect 19588 11930 19728 11990
rect 19788 11930 20128 11990
rect 20188 11930 20528 11990
rect 20588 11930 20928 11990
rect 20988 11930 21008 11990
rect 21068 11930 21328 11990
rect 21388 11930 21528 11990
rect 21588 11930 22128 11990
rect 22188 11930 22198 11990
rect 10878 11920 10958 11930
rect 10878 11860 10888 11920
rect 10948 11910 10958 11920
rect 11598 11920 11678 11930
rect 11598 11910 11608 11920
rect 10948 11870 11608 11910
rect 10948 11860 10958 11870
rect 10878 11850 10958 11860
rect 11598 11860 11608 11870
rect 11668 11910 11678 11920
rect 12318 11920 12398 11930
rect 12318 11910 12328 11920
rect 11668 11870 12328 11910
rect 11668 11860 11678 11870
rect 11598 11850 11678 11860
rect 12318 11860 12328 11870
rect 12388 11860 12398 11920
rect 12318 11850 12398 11860
rect 14158 11920 14238 11930
rect 14158 11860 14168 11920
rect 14228 11910 14238 11920
rect 14878 11920 14958 11930
rect 14878 11910 14888 11920
rect 14228 11870 14888 11910
rect 14228 11860 14238 11870
rect 14158 11850 14238 11860
rect 14878 11860 14888 11870
rect 14948 11910 14958 11920
rect 15598 11920 15678 11930
rect 15598 11910 15608 11920
rect 14948 11870 15608 11910
rect 14948 11860 14958 11870
rect 14878 11850 14958 11860
rect 15598 11860 15608 11870
rect 15668 11860 15678 11920
rect 18038 11920 22198 11930
rect 18038 11910 18278 11920
rect 15598 11850 15678 11860
rect 19918 11880 19998 11890
rect 19918 11820 19928 11880
rect 19988 11820 19998 11880
rect 19918 11810 19998 11820
rect 11368 11590 11428 11620
rect 15128 11590 15188 11630
rect 8448 11580 13138 11590
rect 8448 11520 8458 11580
rect 8518 11520 10648 11580
rect 10708 11520 11368 11580
rect 11428 11520 12088 11580
rect 12148 11520 12808 11580
rect 12868 11520 13068 11580
rect 13128 11520 13138 11580
rect 8448 11510 13138 11520
rect 13418 11580 17648 11590
rect 13418 11520 13428 11580
rect 13488 11520 13688 11580
rect 13748 11520 14408 11580
rect 14468 11520 15128 11580
rect 15188 11520 15848 11580
rect 15908 11520 17578 11580
rect 17638 11520 17648 11580
rect 13418 11510 17648 11520
rect 23438 11580 23548 11600
rect 23438 11510 23458 11580
rect 23528 11510 23548 11580
rect 19618 11500 19698 11510
rect 10518 11470 18278 11480
rect 10518 11410 10528 11470
rect 10588 11410 10768 11470
rect 10828 11410 11008 11470
rect 11068 11410 11248 11470
rect 11308 11410 11488 11470
rect 11548 11410 11728 11470
rect 11788 11410 11968 11470
rect 12028 11410 12208 11470
rect 12268 11410 12448 11470
rect 12508 11410 12688 11470
rect 12748 11410 12928 11470
rect 12988 11410 13568 11470
rect 13628 11410 13808 11470
rect 13868 11410 14048 11470
rect 14108 11410 14288 11470
rect 14348 11410 14528 11470
rect 14588 11410 14768 11470
rect 14828 11410 15008 11470
rect 15068 11410 15248 11470
rect 15308 11410 15488 11470
rect 15548 11410 15728 11470
rect 15788 11410 15968 11470
rect 16028 11440 18278 11470
rect 16028 11410 18078 11440
rect 10518 11390 18078 11410
rect 10518 11330 10528 11390
rect 10588 11330 10768 11390
rect 10828 11330 11008 11390
rect 11068 11330 11248 11390
rect 11308 11330 11488 11390
rect 11548 11330 11728 11390
rect 11788 11330 11968 11390
rect 12028 11330 12208 11390
rect 12268 11330 12448 11390
rect 12508 11330 12688 11390
rect 12748 11330 12928 11390
rect 12988 11330 13568 11390
rect 13628 11330 13808 11390
rect 13868 11330 14048 11390
rect 14108 11330 14288 11390
rect 14348 11330 14528 11390
rect 14588 11330 14768 11390
rect 14828 11330 15008 11390
rect 15068 11330 15248 11390
rect 15308 11330 15488 11390
rect 15548 11330 15728 11390
rect 15788 11330 15968 11390
rect 16028 11380 18078 11390
rect 18138 11380 18178 11440
rect 18238 11380 18278 11440
rect 19618 11440 19628 11500
rect 19688 11440 19698 11500
rect 16028 11340 18278 11380
rect 19028 11410 19108 11420
rect 19028 11350 19038 11410
rect 19098 11400 19108 11410
rect 19618 11400 19698 11440
rect 20058 11500 20138 11510
rect 20058 11440 20068 11500
rect 20128 11440 20138 11500
rect 21898 11500 21978 11510
rect 20058 11430 20138 11440
rect 21128 11480 21208 11490
rect 21128 11420 21138 11480
rect 21198 11470 21208 11480
rect 21898 11470 21908 11500
rect 21198 11440 21908 11470
rect 21968 11440 21978 11500
rect 21198 11430 21978 11440
rect 22738 11500 23298 11510
rect 22738 11440 22748 11500
rect 22808 11440 23228 11500
rect 23288 11440 23298 11500
rect 23438 11490 23548 11510
rect 22738 11430 23298 11440
rect 21198 11420 21208 11430
rect 21128 11410 21208 11420
rect 20718 11400 20728 11410
rect 19098 11360 20728 11400
rect 19098 11350 19108 11360
rect 20718 11350 20728 11360
rect 20788 11350 20798 11410
rect 19028 11340 19108 11350
rect 16028 11330 18078 11340
rect 10518 11310 18078 11330
rect 10518 11250 10528 11310
rect 10588 11250 10768 11310
rect 10828 11250 11008 11310
rect 11068 11250 11248 11310
rect 11308 11250 11488 11310
rect 11548 11250 11728 11310
rect 11788 11250 11968 11310
rect 12028 11250 12208 11310
rect 12268 11250 12448 11310
rect 12508 11250 12688 11310
rect 12748 11250 12928 11310
rect 12988 11250 13568 11310
rect 13628 11250 13808 11310
rect 13868 11250 14048 11310
rect 14108 11250 14288 11310
rect 14348 11250 14528 11310
rect 14588 11250 14768 11310
rect 14828 11250 15008 11310
rect 15068 11250 15248 11310
rect 15308 11250 15488 11310
rect 15548 11250 15728 11310
rect 15788 11250 15968 11310
rect 16028 11280 18078 11310
rect 18138 11280 18178 11340
rect 18238 11280 18278 11340
rect 23608 11330 25968 11340
rect 16028 11250 18278 11280
rect 19968 11270 19978 11330
rect 20038 11320 20048 11330
rect 20038 11280 21978 11320
rect 20038 11270 20048 11280
rect 10518 11240 18278 11250
rect 18918 11250 18998 11260
rect 9568 11200 14758 11210
rect 9568 11140 9578 11200
rect 9638 11140 11808 11200
rect 11868 11140 13248 11200
rect 13308 11140 14688 11200
rect 14748 11140 14758 11200
rect 18918 11190 18928 11250
rect 18988 11240 18998 11250
rect 18988 11230 21278 11240
rect 18988 11200 20068 11230
rect 18988 11190 18998 11200
rect 18918 11180 18998 11190
rect 20058 11170 20068 11200
rect 20128 11200 21278 11230
rect 21898 11220 21908 11280
rect 21968 11220 21978 11280
rect 23608 11270 23618 11330
rect 23678 11270 25898 11330
rect 25958 11270 25968 11330
rect 23608 11260 25968 11270
rect 21898 11210 21978 11220
rect 20128 11170 20138 11200
rect 20058 11160 20138 11170
rect 20758 11160 20838 11170
rect 9568 11130 14758 11140
rect 20758 11100 20768 11160
rect 20828 11100 20838 11160
rect 9458 11090 15788 11100
rect 20758 11090 20838 11100
rect 21198 11160 21278 11200
rect 21198 11100 21208 11160
rect 21268 11100 21278 11160
rect 21198 11090 21278 11100
rect 22738 11160 23298 11170
rect 22738 11100 22748 11160
rect 22808 11100 23228 11160
rect 23288 11100 23298 11160
rect 22738 11090 23298 11100
rect 9458 11030 9468 11090
rect 9528 11030 12168 11090
rect 12228 11030 14328 11090
rect 14388 11030 15718 11090
rect 15778 11030 15788 11090
rect 9458 11020 15788 11030
rect 23438 11070 23548 11090
rect 23438 11000 23458 11070
rect 23528 11000 23548 11070
rect 12518 10980 16318 10990
rect 23438 10980 23548 11000
rect 12518 10920 12528 10980
rect 12588 10920 13968 10980
rect 14028 10920 15248 10980
rect 15308 10920 16248 10980
rect 16308 10920 16318 10980
rect 12518 10910 16318 10920
rect 20978 10880 21058 10890
rect 12878 10870 16228 10880
rect 12878 10810 12888 10870
rect 12948 10810 13608 10870
rect 13668 10810 16158 10870
rect 16218 10810 16228 10870
rect 20978 10820 20988 10880
rect 21048 10820 21058 10880
rect 20978 10810 21058 10820
rect 12878 10800 16228 10810
rect 18338 10780 18578 10790
rect 18338 10770 22198 10780
rect 11898 10760 14658 10770
rect 11958 10700 12078 10760
rect 12138 10700 12258 10760
rect 12318 10700 12438 10760
rect 12498 10700 12618 10760
rect 12678 10700 12798 10760
rect 12858 10700 12978 10760
rect 13038 10700 13158 10760
rect 13218 10700 13338 10760
rect 13398 10700 13428 10760
rect 13488 10700 13518 10760
rect 13578 10700 13698 10760
rect 13758 10700 13878 10760
rect 13938 10700 14058 10760
rect 14118 10700 14238 10760
rect 14298 10700 14418 10760
rect 14478 10700 14598 10760
rect 11898 10690 14658 10700
rect 18338 10710 18378 10770
rect 18438 10710 18478 10770
rect 18538 10710 19408 10770
rect 19468 10710 19608 10770
rect 19668 10710 19848 10770
rect 19908 10710 20008 10770
rect 20068 10710 20408 10770
rect 20468 10710 20808 10770
rect 20868 10710 21208 10770
rect 21268 10710 21408 10770
rect 21468 10710 22128 10770
rect 22188 10710 22198 10770
rect 18338 10700 22198 10710
rect 18338 10690 18578 10700
rect 20978 10660 21058 10670
rect 20978 10600 20988 10660
rect 21048 10600 21058 10660
rect 20978 10590 21058 10600
rect 15588 10560 15908 10570
rect 15588 10500 15598 10560
rect 15658 10500 15838 10560
rect 15898 10500 15908 10560
rect 15588 10490 15908 10500
rect 15238 10220 15318 10230
rect 15238 10160 15248 10220
rect 15308 10210 15318 10220
rect 15708 10220 15788 10230
rect 15708 10210 15718 10220
rect 15308 10170 15718 10210
rect 15308 10160 15318 10170
rect 15238 10150 15318 10160
rect 15708 10160 15718 10170
rect 15778 10160 15788 10220
rect 15708 10150 15788 10160
rect 11618 10020 18278 10030
rect 11618 9960 11628 10020
rect 11688 9960 11988 10020
rect 12048 9960 12348 10020
rect 12408 9960 12708 10020
rect 12768 9960 13068 10020
rect 13128 9960 13428 10020
rect 13488 9960 13788 10020
rect 13848 9960 14148 10020
rect 14208 9960 14508 10020
rect 14568 9960 14868 10020
rect 14928 9960 15498 10020
rect 15558 9960 15938 10020
rect 15998 9990 18278 10020
rect 15998 9960 18078 9990
rect 11618 9940 18078 9960
rect 11618 9880 11628 9940
rect 11688 9880 11988 9940
rect 12048 9880 12348 9940
rect 12408 9880 12708 9940
rect 12768 9880 13068 9940
rect 13128 9880 13428 9940
rect 13488 9880 13788 9940
rect 13848 9880 14148 9940
rect 14208 9880 14508 9940
rect 14568 9880 14868 9940
rect 14928 9880 15498 9940
rect 15558 9880 15938 9940
rect 15998 9930 18078 9940
rect 18138 9930 18178 9990
rect 18238 9930 18278 9990
rect 15998 9890 18278 9930
rect 15998 9880 18078 9890
rect 11618 9860 18078 9880
rect 11618 9800 11628 9860
rect 11688 9800 11988 9860
rect 12048 9800 12348 9860
rect 12408 9800 12708 9860
rect 12768 9800 13068 9860
rect 13128 9800 13428 9860
rect 13488 9800 13788 9860
rect 13848 9800 14148 9860
rect 14208 9800 14508 9860
rect 14568 9800 14868 9860
rect 14928 9800 15498 9860
rect 15558 9800 15938 9860
rect 15998 9830 18078 9860
rect 18138 9830 18178 9890
rect 18238 9830 18278 9890
rect 15998 9800 18278 9830
rect 11618 9790 18278 9800
rect 8448 9700 8458 9760
rect 8518 9750 14752 9760
rect 8518 9700 11806 9750
rect 8448 9698 11806 9700
rect 11858 9698 11916 9750
rect 11968 9698 12026 9750
rect 12078 9698 12136 9750
rect 12188 9698 12246 9750
rect 12298 9698 12356 9750
rect 12408 9698 12466 9750
rect 12518 9698 12576 9750
rect 12628 9698 12686 9750
rect 12738 9698 12796 9750
rect 12848 9698 13706 9750
rect 13758 9698 13816 9750
rect 13868 9698 13926 9750
rect 13978 9698 14036 9750
rect 14088 9698 14146 9750
rect 14198 9698 14256 9750
rect 14308 9698 14366 9750
rect 14418 9698 14476 9750
rect 14528 9698 14586 9750
rect 14638 9698 14696 9750
rect 14748 9698 14752 9750
rect 8448 9690 14752 9698
rect 18338 9650 23088 9660
rect 18338 9590 18378 9650
rect 18438 9590 18478 9650
rect 18538 9590 23018 9650
rect 23078 9590 23088 9650
rect 18338 9580 23088 9590
rect 18038 9430 18278 9440
rect 11628 9420 18278 9430
rect 11628 9360 11638 9420
rect 11698 9360 11858 9420
rect 11918 9360 12078 9420
rect 12138 9360 12298 9420
rect 12358 9360 12518 9420
rect 12578 9360 12738 9420
rect 12798 9360 12958 9420
rect 13018 9360 13538 9420
rect 13598 9360 13758 9420
rect 13818 9360 13978 9420
rect 14038 9360 14198 9420
rect 14258 9360 14418 9420
rect 14478 9360 14638 9420
rect 14698 9360 14858 9420
rect 14918 9360 18078 9420
rect 18138 9360 18178 9420
rect 18238 9360 18278 9420
rect 11628 9350 18278 9360
rect 18038 9340 18278 9350
rect 9678 9310 12918 9320
rect 9678 9250 9688 9310
rect 9748 9250 11748 9310
rect 11808 9250 11968 9310
rect 12028 9250 12188 9310
rect 12248 9250 12408 9310
rect 12468 9250 12628 9310
rect 12688 9250 12848 9310
rect 12908 9250 12918 9310
rect 9678 9240 12918 9250
rect 13638 9300 18888 9310
rect 13638 9240 13648 9300
rect 13708 9240 13868 9300
rect 13928 9240 14088 9300
rect 14148 9240 14308 9300
rect 14368 9240 14528 9300
rect 14588 9240 14748 9300
rect 14808 9240 18658 9300
rect 18718 9240 18738 9300
rect 18798 9240 18818 9300
rect 18878 9240 18888 9300
rect 13638 9220 18888 9240
rect 13638 9160 13648 9220
rect 13708 9160 13868 9220
rect 13928 9160 14088 9220
rect 14148 9160 14308 9220
rect 14368 9160 14528 9220
rect 14588 9160 14748 9220
rect 14808 9160 18658 9220
rect 18718 9160 18738 9220
rect 18798 9160 18818 9220
rect 18878 9160 18888 9220
rect 13638 9140 18888 9160
rect 13638 9080 13648 9140
rect 13708 9080 13868 9140
rect 13928 9080 14088 9140
rect 14148 9080 14308 9140
rect 14368 9080 14528 9140
rect 14588 9080 14748 9140
rect 14808 9080 18658 9140
rect 18718 9080 18738 9140
rect 18798 9080 18818 9140
rect 18878 9080 18888 9140
rect 13638 9070 18888 9080
rect 23208 9130 23308 9150
rect 23208 9070 23228 9130
rect 23288 9070 23308 9130
rect 23208 9050 23308 9070
rect 19028 8770 26478 8780
rect 19028 8710 19038 8770
rect 19098 8710 26008 8770
rect 26068 8710 26088 8770
rect 26148 8710 26168 8770
rect 26228 8710 26248 8770
rect 26308 8710 26328 8770
rect 26388 8710 26408 8770
rect 26468 8710 26478 8770
rect 19028 8690 26478 8710
rect 19028 8630 19038 8690
rect 19098 8630 26008 8690
rect 26068 8630 26088 8690
rect 26148 8630 26168 8690
rect 26228 8630 26248 8690
rect 26308 8630 26328 8690
rect 26388 8630 26408 8690
rect 26468 8630 26478 8690
rect 19028 8610 26478 8630
rect 19028 8550 19038 8610
rect 19098 8550 26008 8610
rect 26068 8550 26088 8610
rect 26148 8550 26168 8610
rect 26228 8550 26248 8610
rect 26308 8550 26328 8610
rect 26388 8550 26408 8610
rect 26468 8550 26478 8610
rect 19028 8540 26478 8550
rect 19138 8500 25968 8510
rect 19138 8440 19148 8500
rect 19208 8440 25898 8500
rect 25958 8440 25968 8500
rect 19138 8430 25968 8440
rect 12908 8350 13008 8390
rect 23088 8380 23198 8400
rect 12908 8290 12928 8350
rect 12988 8310 13008 8350
rect 18098 8370 23108 8380
rect 18098 8310 18108 8370
rect 18168 8310 23108 8370
rect 23178 8310 23198 8380
rect 12988 8300 17928 8310
rect 18098 8300 23198 8310
rect 12988 8290 13258 8300
rect 12908 8250 13258 8290
rect 12908 8190 12928 8250
rect 12988 8240 13258 8250
rect 13318 8240 13478 8300
rect 13538 8240 13778 8300
rect 13838 8240 14008 8300
rect 14068 8240 14158 8300
rect 14218 8240 14378 8300
rect 14438 8240 14678 8300
rect 14738 8240 14898 8300
rect 14958 8240 15298 8300
rect 15358 8240 15628 8300
rect 15688 8240 15958 8300
rect 16018 8240 16398 8300
rect 16458 8240 16658 8300
rect 16718 8240 17178 8300
rect 17238 8240 17858 8300
rect 17918 8240 17928 8300
rect 23088 8290 23198 8300
rect 12988 8230 17928 8240
rect 18338 8230 22458 8240
rect 12988 8190 13008 8230
rect 12908 8150 13008 8190
rect 16898 8190 16978 8200
rect 16898 8130 16908 8190
rect 16968 8130 16978 8190
rect 16898 8120 16978 8130
rect 17528 8190 18178 8200
rect 17528 8130 17538 8190
rect 17598 8130 18108 8190
rect 18168 8130 18178 8190
rect 18338 8170 18378 8230
rect 18438 8170 18478 8230
rect 18538 8170 19348 8230
rect 19408 8170 19568 8230
rect 19628 8170 20008 8230
rect 20068 8170 20328 8230
rect 20388 8170 20648 8230
rect 20708 8170 21088 8230
rect 21148 8170 21408 8230
rect 21468 8170 21728 8230
rect 21788 8170 22168 8230
rect 22228 8170 22388 8230
rect 22448 8170 22458 8230
rect 18338 8160 22458 8170
rect 17528 8120 18178 8130
rect 17998 7850 18258 7860
rect 12108 7810 13208 7820
rect 12108 7750 12118 7810
rect 12178 7750 13138 7810
rect 13198 7750 13208 7810
rect 12108 7740 13208 7750
rect 15048 7800 15128 7810
rect 15048 7740 15058 7800
rect 15118 7740 15128 7800
rect 15048 7730 15128 7740
rect 16078 7800 16158 7810
rect 16078 7740 16088 7800
rect 16148 7740 16158 7800
rect 17998 7790 18008 7850
rect 18068 7790 18188 7850
rect 18248 7790 18258 7850
rect 17998 7780 18258 7790
rect 16078 7730 16158 7740
rect 22738 7590 22848 7610
rect 22738 7580 22758 7590
rect 21808 7570 21888 7580
rect 21808 7510 21818 7570
rect 21878 7510 21888 7570
rect 21808 7500 21888 7510
rect 22068 7570 22758 7580
rect 22068 7510 22078 7570
rect 22138 7520 22758 7570
rect 22828 7520 22848 7590
rect 22138 7510 22848 7520
rect 22068 7500 22848 7510
rect 18178 7490 21888 7500
rect 18178 7430 18188 7490
rect 18248 7430 21888 7490
rect 18178 7420 21888 7430
rect 18178 7380 19858 7390
rect 18178 7320 18188 7380
rect 18248 7320 18658 7380
rect 18718 7320 18738 7380
rect 18798 7320 18818 7380
rect 18878 7320 19788 7380
rect 19848 7320 19858 7380
rect 18178 7310 19858 7320
rect 21938 7320 26478 7330
rect 18288 7270 21448 7280
rect 16228 7240 16308 7250
rect 13698 7230 13778 7240
rect 12908 7170 13008 7210
rect 12908 7110 12928 7170
rect 12988 7130 13008 7170
rect 13698 7170 13708 7230
rect 13768 7220 13778 7230
rect 15228 7230 15308 7240
rect 16228 7230 16238 7240
rect 15228 7220 15238 7230
rect 13768 7180 15238 7220
rect 13768 7170 13778 7180
rect 13698 7160 13778 7170
rect 15228 7170 15238 7180
rect 15298 7190 16238 7230
rect 15298 7170 15308 7190
rect 16228 7180 16238 7190
rect 16298 7180 16308 7240
rect 16818 7230 16898 7240
rect 16228 7170 16308 7180
rect 16648 7170 16658 7230
rect 16718 7220 16728 7230
rect 16818 7220 16828 7230
rect 16718 7180 16828 7220
rect 16718 7170 16728 7180
rect 16818 7170 16828 7180
rect 16888 7170 16898 7230
rect 17458 7230 18258 7240
rect 17458 7170 17468 7230
rect 17528 7170 18188 7230
rect 18248 7170 18258 7230
rect 18288 7210 18298 7270
rect 18358 7210 21378 7270
rect 21438 7210 21448 7270
rect 21938 7260 21948 7320
rect 22008 7260 26008 7320
rect 26068 7260 26088 7320
rect 26148 7260 26168 7320
rect 26228 7260 26248 7320
rect 26308 7260 26328 7320
rect 26388 7260 26408 7320
rect 26468 7260 26478 7320
rect 21938 7250 26478 7260
rect 18288 7200 21448 7210
rect 15228 7160 15308 7170
rect 17458 7160 18258 7170
rect 18398 7160 20278 7170
rect 12988 7120 17928 7130
rect 12988 7110 13258 7120
rect 12908 7070 13258 7110
rect 12908 7010 12928 7070
rect 12988 7060 13258 7070
rect 13318 7060 13998 7120
rect 14058 7060 14158 7120
rect 14218 7060 14898 7120
rect 14958 7060 15148 7120
rect 15208 7060 15338 7120
rect 15398 7060 15418 7120
rect 15478 7060 15628 7120
rect 15688 7060 15958 7120
rect 16018 7060 16398 7120
rect 16458 7060 16788 7120
rect 16848 7060 16998 7120
rect 17058 7060 17178 7120
rect 17238 7060 17858 7120
rect 17918 7060 17928 7120
rect 18398 7100 18408 7160
rect 18468 7100 19148 7160
rect 19208 7100 20208 7160
rect 20268 7100 20278 7160
rect 18398 7090 20278 7100
rect 12988 7050 17928 7060
rect 21368 7070 21448 7080
rect 12988 7010 13008 7050
rect 18918 7040 20938 7050
rect 12908 6970 13008 7010
rect 15248 6950 15258 7010
rect 15318 6950 15328 7010
rect 18918 6980 18928 7040
rect 18988 6980 19988 7040
rect 20048 6980 20428 7040
rect 20488 6980 20868 7040
rect 20928 6980 20938 7040
rect 21368 7010 21378 7070
rect 21438 7010 21448 7070
rect 22068 7070 22848 7080
rect 21368 7000 21448 7010
rect 21498 7040 22018 7050
rect 18918 6970 20938 6980
rect 21498 6980 21508 7040
rect 21568 6980 21948 7040
rect 22008 6980 22018 7040
rect 22068 7010 22078 7070
rect 22138 7060 22848 7070
rect 22138 7010 22758 7060
rect 22068 7000 22758 7010
rect 21498 6970 22018 6980
rect 22738 6990 22758 7000
rect 22828 6990 22848 7060
rect 22738 6970 22848 6990
rect 15248 6940 15328 6950
rect 17688 6470 17768 6480
rect 16118 6440 16198 6450
rect 11938 6430 13208 6440
rect 11938 6370 11948 6430
rect 12008 6370 13138 6430
rect 13198 6370 13208 6430
rect 11938 6360 13208 6370
rect 15028 6400 15108 6410
rect 15028 6340 15038 6400
rect 15098 6340 15108 6400
rect 16118 6380 16128 6440
rect 16188 6380 16198 6440
rect 17688 6410 17698 6470
rect 17758 6410 17768 6470
rect 17688 6400 17768 6410
rect 16118 6370 16198 6380
rect 17998 6390 18368 6400
rect 15028 6330 15108 6340
rect 17998 6330 18008 6390
rect 18068 6330 18298 6390
rect 18358 6330 18368 6390
rect 17998 6320 18368 6330
rect 19238 6390 22458 6400
rect 19238 6330 19278 6390
rect 19338 6330 19378 6390
rect 19438 6330 19548 6390
rect 19608 6330 19768 6390
rect 19828 6330 20208 6390
rect 20268 6330 20648 6390
rect 20708 6330 20968 6390
rect 21028 6330 21288 6390
rect 21348 6330 21728 6390
rect 21788 6330 22168 6390
rect 22228 6330 22388 6390
rect 22448 6330 22458 6390
rect 19238 6320 22458 6330
rect 16228 6070 16308 6080
rect 16228 6060 16238 6070
rect 13658 6050 16238 6060
rect 12908 5990 13008 6030
rect 12908 5930 12928 5990
rect 12988 5950 13008 5990
rect 13658 5990 13668 6050
rect 13728 6020 15388 6050
rect 13728 5990 13738 6020
rect 13658 5980 13738 5990
rect 15378 5990 15388 6020
rect 15448 6020 16238 6050
rect 15448 5990 15458 6020
rect 16228 6010 16238 6020
rect 16298 6010 16308 6070
rect 16228 6000 16308 6010
rect 17458 6050 18478 6060
rect 15378 5980 15458 5990
rect 17458 5990 17468 6050
rect 17528 5990 18408 6050
rect 18468 5990 18478 6050
rect 17458 5980 18478 5990
rect 12988 5940 17248 5950
rect 12988 5930 13258 5940
rect 12908 5890 13258 5930
rect 12908 5830 12928 5890
rect 12988 5880 13258 5890
rect 13318 5880 13478 5940
rect 13538 5880 13778 5940
rect 13838 5880 13998 5940
rect 14058 5880 14158 5940
rect 14218 5880 14378 5940
rect 14438 5880 14678 5940
rect 14738 5880 14898 5940
rect 14958 5880 15198 5940
rect 15258 5880 15638 5940
rect 15698 5880 15968 5940
rect 16028 5880 16398 5940
rect 16458 5880 16788 5940
rect 16848 5880 17178 5940
rect 17238 5880 17248 5940
rect 22978 5890 23088 5900
rect 12988 5870 17248 5880
rect 17688 5880 23088 5890
rect 12988 5830 13008 5870
rect 12908 5790 13008 5830
rect 17688 5820 17698 5880
rect 17758 5820 22998 5880
rect 17688 5810 22998 5820
rect 23068 5810 23088 5880
rect 22978 5790 23088 5810
rect 22588 5690 22688 5730
rect 22588 5630 22608 5690
rect 22668 5650 22688 5690
rect 22668 5640 25218 5650
rect 22668 5630 23588 5640
rect 22588 5590 23588 5630
rect 22588 5530 22608 5590
rect 22668 5580 23588 5590
rect 23648 5580 24108 5640
rect 24168 5580 24628 5640
rect 24688 5580 25148 5640
rect 25208 5580 25218 5640
rect 22668 5570 25218 5580
rect 22668 5530 22688 5570
rect 22588 5490 22688 5530
rect 23388 4990 25018 5000
rect 23388 4930 23398 4990
rect 23458 4930 23918 4990
rect 23978 4930 24438 4990
rect 24498 4930 24768 4990
rect 24828 4930 24958 4990
rect 23388 4920 25018 4930
rect 23308 4810 23658 4820
rect 23308 4750 23318 4810
rect 23378 4750 23588 4810
rect 23648 4750 23658 4810
rect 23308 4740 23658 4750
rect 23828 4810 24178 4820
rect 23828 4750 23838 4810
rect 23898 4750 24108 4810
rect 24168 4750 24178 4810
rect 23828 4740 24178 4750
rect 24348 4810 24698 4820
rect 24348 4750 24358 4810
rect 24418 4750 24628 4810
rect 24688 4750 24698 4810
rect 24348 4740 24698 4750
rect 23318 4220 23488 4230
rect 23378 4160 23418 4220
rect 23478 4160 23488 4220
rect 23318 4150 23488 4160
rect 23838 4220 24008 4230
rect 23898 4160 23938 4220
rect 23998 4160 24008 4220
rect 23838 4150 24008 4160
rect 24358 4220 24528 4230
rect 24418 4160 24458 4220
rect 24518 4160 24528 4220
rect 24358 4150 24528 4160
rect 23278 4100 23598 4110
rect 23278 4048 23282 4100
rect 23334 4048 23528 4100
rect 23278 4040 23528 4048
rect 23588 4040 23598 4100
rect 23798 4100 24118 4110
rect 23798 4048 23802 4100
rect 23854 4048 24048 4100
rect 23798 4040 24048 4048
rect 24108 4040 24118 4100
rect 24318 4100 24638 4110
rect 24318 4048 24322 4100
rect 24374 4048 24568 4100
rect 24318 4040 24568 4048
rect 24628 4040 24638 4100
rect 23518 4030 23598 4040
rect 24038 4030 24118 4040
rect 24558 4030 24638 4040
rect 12218 3790 12318 3830
rect 12218 3730 12238 3790
rect 12298 3750 12318 3790
rect 12298 3740 22618 3750
rect 12298 3730 12708 3740
rect 12218 3690 12708 3730
rect 12218 3630 12238 3690
rect 12298 3680 12708 3690
rect 12768 3680 13128 3740
rect 13188 3680 13798 3740
rect 13858 3680 14368 3740
rect 14428 3680 15078 3740
rect 15138 3680 15508 3740
rect 15568 3680 15948 3740
rect 16008 3680 16198 3740
rect 16258 3680 16418 3740
rect 16478 3680 16888 3740
rect 16948 3680 17328 3740
rect 17388 3680 17948 3740
rect 18008 3680 18288 3740
rect 18348 3680 18648 3740
rect 18708 3680 19248 3740
rect 19308 3680 19588 3740
rect 19648 3680 19948 3740
rect 20008 3680 20548 3740
rect 20608 3680 20888 3740
rect 20948 3680 21248 3740
rect 21308 3680 21848 3740
rect 21908 3680 22188 3740
rect 22248 3680 22548 3740
rect 22608 3680 22618 3740
rect 12298 3670 22618 3680
rect 12298 3630 12318 3670
rect 12218 3590 12318 3630
rect 22808 3410 23308 3420
rect 22808 3350 22818 3410
rect 22878 3350 22898 3410
rect 22958 3350 22978 3410
rect 23038 3350 23248 3410
rect 12108 3340 12398 3350
rect 22808 3340 23308 3350
rect 12108 3280 12118 3340
rect 12178 3280 12328 3340
rect 12388 3280 12398 3340
rect 12108 3270 12398 3280
rect 22750 3330 23308 3340
rect 22750 3278 22754 3330
rect 22806 3278 22818 3330
rect 22750 3270 22818 3278
rect 22878 3270 22898 3330
rect 22958 3270 22978 3330
rect 23038 3270 23248 3330
rect 22750 3260 23308 3270
rect 22808 3250 23308 3260
rect 22808 3190 22818 3250
rect 22878 3190 22898 3250
rect 22958 3190 22978 3250
rect 23038 3190 23248 3250
rect 22808 3180 23308 3190
rect 23338 3410 23828 3420
rect 23398 3350 23768 3410
rect 23338 3330 23828 3350
rect 23398 3270 23768 3330
rect 23338 3250 23828 3270
rect 23398 3190 23768 3250
rect 23338 3180 23828 3190
rect 23858 3410 24348 3420
rect 23918 3350 24288 3410
rect 23858 3330 24348 3350
rect 23918 3270 24288 3330
rect 23858 3250 24348 3270
rect 23918 3190 24288 3250
rect 23858 3180 24348 3190
rect 24378 3410 26668 3420
rect 24438 3350 25178 3410
rect 25238 3350 25258 3410
rect 25318 3350 25338 3410
rect 25398 3400 26668 3410
rect 25398 3350 26548 3400
rect 24378 3330 26548 3350
rect 24438 3270 25178 3330
rect 25238 3270 25258 3330
rect 25318 3270 25338 3330
rect 25398 3320 26548 3330
rect 26628 3320 26668 3400
rect 25398 3280 26668 3320
rect 25398 3270 26548 3280
rect 24378 3250 26548 3270
rect 24438 3190 25178 3250
rect 25238 3190 25258 3250
rect 25318 3190 25338 3250
rect 25398 3200 26548 3250
rect 26628 3200 26668 3280
rect 25398 3190 26668 3200
rect 24378 3180 26668 3190
rect 12218 3010 12318 3050
rect 12218 2950 12238 3010
rect 12298 2970 12318 3010
rect 12298 2960 22618 2970
rect 12298 2950 12548 2960
rect 12218 2910 12548 2950
rect 12218 2850 12238 2910
rect 12298 2900 12548 2910
rect 12608 2900 12768 2960
rect 12828 2900 13238 2960
rect 13298 2900 13578 2960
rect 13638 2900 13798 2960
rect 13858 2900 14238 2960
rect 14298 2900 14918 2960
rect 14978 2900 15138 2960
rect 15198 2900 15608 2960
rect 15668 2900 16068 2960
rect 16128 2900 16418 2960
rect 16478 2900 16668 2960
rect 16728 2900 16888 2960
rect 16948 2900 17218 2960
rect 17278 2900 17878 2960
rect 17938 2900 18098 2960
rect 18158 2900 18668 2960
rect 18728 2900 18928 2960
rect 18988 2900 19178 2960
rect 19238 2900 19398 2960
rect 19458 2900 19948 2960
rect 20008 2900 20228 2960
rect 20288 2900 20478 2960
rect 20538 2900 20698 2960
rect 20758 2900 21248 2960
rect 21308 2900 21528 2960
rect 21588 2900 21778 2960
rect 21838 2900 21998 2960
rect 22058 2900 22548 2960
rect 22608 2900 22618 2960
rect 12298 2890 22618 2900
rect 12298 2850 12318 2890
rect 12218 2810 12318 2850
rect 23408 2760 23488 2770
rect 23928 2760 24008 2770
rect 24448 2760 24528 2770
rect 23278 2750 23418 2760
rect 23278 2698 23282 2750
rect 23334 2700 23418 2750
rect 23478 2700 23488 2760
rect 23334 2698 23488 2700
rect 23278 2690 23488 2698
rect 23798 2750 23938 2760
rect 23798 2698 23802 2750
rect 23854 2700 23938 2750
rect 23998 2700 24008 2760
rect 23854 2698 24008 2700
rect 23798 2690 24008 2698
rect 24318 2750 24458 2760
rect 24318 2698 24322 2750
rect 24374 2700 24458 2750
rect 24518 2700 24528 2760
rect 24374 2698 24528 2700
rect 24318 2690 24528 2698
rect 23318 2640 23598 2650
rect 23378 2580 23528 2640
rect 23588 2580 23598 2640
rect 23318 2570 23598 2580
rect 23838 2640 24118 2650
rect 23898 2580 24048 2640
rect 24108 2580 24118 2640
rect 23838 2570 24118 2580
rect 24358 2640 24638 2650
rect 24418 2580 24568 2640
rect 24628 2580 24638 2640
rect 24358 2570 24638 2580
rect 23263 2270 26008 2280
rect 23263 2218 23268 2270
rect 23320 2218 23788 2270
rect 23840 2218 24308 2270
rect 24360 2218 24874 2270
rect 24926 2220 26008 2270
rect 26068 2220 26088 2280
rect 26148 2220 26168 2280
rect 26228 2220 26248 2280
rect 26308 2220 26328 2280
rect 26388 2220 26408 2280
rect 26468 2220 26478 2280
rect 24926 2218 26478 2220
rect 23263 2210 26478 2218
rect 22808 1830 25408 1840
rect 22808 1770 22818 1830
rect 22878 1770 22898 1830
rect 22958 1770 22978 1830
rect 23038 1770 25178 1830
rect 25238 1770 25258 1830
rect 25318 1770 25338 1830
rect 25398 1770 25408 1830
rect 22808 1750 25408 1770
rect 22808 1690 22818 1750
rect 22878 1690 22898 1750
rect 22958 1690 22978 1750
rect 23038 1690 25178 1750
rect 25238 1690 25258 1750
rect 25318 1690 25338 1750
rect 25398 1690 25408 1750
rect 22808 1670 25408 1690
rect 22588 1610 22688 1650
rect 22588 1550 22608 1610
rect 22668 1570 22688 1610
rect 22808 1610 22818 1670
rect 22878 1610 22898 1670
rect 22958 1610 22978 1670
rect 23038 1610 25178 1670
rect 25238 1610 25258 1670
rect 25318 1610 25338 1670
rect 25398 1610 25408 1670
rect 22808 1600 25408 1610
rect 22668 1560 24918 1570
rect 22668 1550 23318 1560
rect 22588 1510 23318 1550
rect 22588 1450 22608 1510
rect 22668 1500 23318 1510
rect 23378 1500 23838 1560
rect 23898 1500 24358 1560
rect 24418 1500 24848 1560
rect 24908 1500 24918 1560
rect 22668 1490 24918 1500
rect 22668 1450 22688 1490
rect 22588 1410 22688 1450
rect 30368 1340 30528 1380
rect 11938 1330 30408 1340
rect 11938 1270 11948 1330
rect 12008 1270 30408 1330
rect 11938 1260 30408 1270
rect 30488 1260 30528 1340
rect 30368 1220 30528 1260
<< via2 >>
rect 7468 19820 7528 19880
rect 7558 19820 7618 19880
rect 7648 19820 7708 19880
rect 7468 19730 7528 19790
rect 7558 19730 7618 19790
rect 7648 19730 7708 19790
rect 22818 19720 22888 19790
rect 23318 19720 23388 19790
rect 7468 19640 7528 19700
rect 7558 19640 7618 19700
rect 7648 19640 7708 19700
rect 8938 19440 8998 19500
rect 26008 19440 26068 19500
rect 7468 18990 7528 19050
rect 7558 18990 7618 19050
rect 7648 18990 7708 19050
rect 7468 18890 7528 18950
rect 7558 18890 7618 18950
rect 7648 18890 7708 18950
rect 18198 18790 18258 18850
rect 18658 18090 18718 18150
rect 18128 17390 18188 17450
rect 18798 16690 18858 16750
rect 18998 15990 19058 16050
rect 18798 15290 18858 15350
rect 18378 14150 18438 14210
rect 18478 14150 18538 14210
rect 18378 13840 18438 13900
rect 18478 13840 18538 13900
rect 18378 13740 18438 13800
rect 18478 13740 18538 13800
rect 23228 13450 23288 13510
rect 18078 13360 18138 13420
rect 18178 13360 18238 13420
rect 18378 13120 18438 13180
rect 18478 13120 18538 13180
rect 18078 13040 18138 13100
rect 18178 13040 18238 13100
rect 18078 12940 18138 13000
rect 18178 12940 18238 13000
rect 18078 11930 18138 11990
rect 18178 11930 18238 11990
rect 23458 11510 23528 11580
rect 18078 11380 18138 11440
rect 18178 11380 18238 11440
rect 18078 11280 18138 11340
rect 18178 11280 18238 11340
rect 23458 11000 23528 11070
rect 18378 10710 18438 10770
rect 18478 10710 18538 10770
rect 18078 9930 18138 9990
rect 18178 9930 18238 9990
rect 18078 9830 18138 9890
rect 18178 9830 18238 9890
rect 18378 9590 18438 9650
rect 18478 9590 18538 9650
rect 18078 9360 18138 9420
rect 18178 9360 18238 9420
rect 23228 9070 23288 9130
rect 12928 8290 12988 8350
rect 23108 8310 23178 8380
rect 12928 8190 12988 8250
rect 18378 8170 18438 8230
rect 18478 8170 18538 8230
rect 22758 7520 22828 7590
rect 12928 7110 12988 7170
rect 12928 7010 12988 7070
rect 22758 6990 22828 7060
rect 19278 6330 19338 6390
rect 19378 6330 19438 6390
rect 12928 5930 12988 5990
rect 12928 5830 12988 5890
rect 22998 5810 23068 5880
rect 22608 5630 22668 5690
rect 22608 5530 22668 5590
rect 12238 3730 12298 3790
rect 12238 3630 12298 3690
rect 26548 3320 26628 3400
rect 26548 3200 26628 3280
rect 12238 2950 12298 3010
rect 12238 2850 12298 2910
rect 22608 1550 22668 1610
rect 22608 1450 22668 1510
rect 30408 1260 30488 1340
<< metal3 >>
rect 8918 20050 22938 32110
rect 23268 20050 26088 32110
rect 798 19880 7718 19890
rect 798 19860 7468 19880
rect 798 19780 808 19860
rect 888 19780 908 19860
rect 988 19780 1008 19860
rect 1088 19780 1108 19860
rect 1188 19820 7468 19860
rect 7528 19820 7558 19880
rect 7618 19820 7648 19880
rect 7708 19820 7718 19880
rect 1188 19790 7718 19820
rect 1188 19780 7468 19790
rect 798 19740 7468 19780
rect 798 19660 808 19740
rect 888 19660 908 19740
rect 988 19660 1008 19740
rect 1088 19660 1108 19740
rect 1188 19730 7468 19740
rect 7528 19730 7558 19790
rect 7618 19730 7648 19790
rect 7708 19730 7718 19790
rect 1188 19700 7718 19730
rect 1188 19660 7468 19700
rect 798 19640 7468 19660
rect 7528 19640 7558 19700
rect 7618 19640 7648 19700
rect 7708 19640 7718 19700
rect 798 19630 7718 19640
rect 8918 19500 9018 20050
rect 22798 19790 22908 19810
rect 22798 19720 22818 19790
rect 22888 19720 22908 19790
rect 22798 19700 22908 19720
rect 23298 19790 23408 19810
rect 23298 19720 23318 19790
rect 23388 19720 23408 19790
rect 23298 19700 23408 19720
rect 8918 19440 8938 19500
rect 8998 19440 9018 19500
rect 8918 19420 9018 19440
rect 25988 19500 26088 20050
rect 25988 19440 26008 19500
rect 26068 19440 26088 19500
rect 25988 19420 26088 19440
rect 798 19060 7718 19090
rect 798 18980 808 19060
rect 888 18980 908 19060
rect 988 18980 1008 19060
rect 1088 18980 1108 19060
rect 1188 19050 7718 19060
rect 1188 18990 7468 19050
rect 7528 18990 7558 19050
rect 7618 18990 7648 19050
rect 7708 18990 7718 19050
rect 1188 18980 7718 18990
rect 798 18960 7718 18980
rect 798 18880 808 18960
rect 888 18880 908 18960
rect 988 18880 1008 18960
rect 1088 18880 1108 18960
rect 1188 18950 7718 18960
rect 1188 18890 7468 18950
rect 7528 18890 7558 18950
rect 7618 18890 7648 18950
rect 7708 18890 7718 18950
rect 1188 18880 7718 18890
rect 798 18850 7718 18880
rect 19118 18870 19578 19040
rect 19818 18870 20278 19040
rect 20518 18870 20978 19040
rect 21218 18870 21678 19040
rect 21918 18870 22378 19040
rect 22618 18870 23078 19040
rect 23318 18870 23778 19040
rect 24018 18870 24478 19040
rect 24718 18870 25178 19040
rect 25418 18870 25878 19040
rect 19118 18860 25878 18870
rect 18188 18850 25878 18860
rect 18188 18790 18198 18850
rect 18258 18790 25878 18850
rect 18188 18780 25878 18790
rect 19118 18770 25878 18780
rect 19118 18580 19578 18770
rect 19818 18580 20278 18770
rect 20518 18580 20978 18770
rect 21218 18580 21678 18770
rect 21918 18580 22378 18770
rect 22618 18580 23078 18770
rect 23318 18580 23778 18770
rect 24018 18580 24478 18770
rect 24718 18580 25178 18770
rect 25418 18580 25878 18770
rect 25598 18340 25698 18580
rect 19118 18170 19578 18340
rect 19818 18170 20278 18340
rect 20518 18170 20978 18340
rect 21218 18170 21678 18340
rect 21918 18170 22378 18340
rect 22618 18170 23078 18340
rect 23318 18170 23778 18340
rect 24018 18170 24478 18340
rect 24718 18170 25178 18340
rect 25418 18170 25878 18340
rect 18638 18160 18738 18170
rect 18638 18080 18648 18160
rect 18728 18080 18738 18160
rect 18638 18070 18738 18080
rect 19118 18070 25878 18170
rect 19118 17880 19578 18070
rect 19818 17880 20278 18070
rect 20518 17880 20978 18070
rect 21218 17880 21678 18070
rect 21918 17880 22378 18070
rect 22618 17880 23078 18070
rect 23318 17880 23778 18070
rect 24018 17880 24478 18070
rect 24718 17880 25178 18070
rect 25418 17880 25878 18070
rect 19118 17470 19578 17640
rect 19818 17470 20278 17640
rect 20518 17470 20978 17640
rect 21218 17470 21678 17640
rect 21918 17470 22378 17640
rect 22618 17470 23078 17640
rect 23318 17470 23778 17640
rect 24018 17470 24478 17640
rect 24718 17470 25178 17640
rect 25418 17470 25878 17640
rect 19118 17460 25878 17470
rect 18118 17450 25878 17460
rect 18118 17390 18128 17450
rect 18188 17390 25878 17450
rect 18118 17380 25878 17390
rect 19118 17370 25878 17380
rect 19118 17180 19578 17370
rect 19818 17180 20278 17370
rect 20518 17180 20978 17370
rect 21218 17180 21678 17370
rect 21918 17180 22378 17370
rect 22618 17180 23078 17370
rect 23318 17180 23778 17370
rect 24018 17180 24478 17370
rect 24718 17180 25178 17370
rect 25418 17180 25878 17370
rect 25598 16940 25698 17180
rect 19118 16770 19578 16940
rect 19818 16770 20278 16940
rect 20518 16770 20978 16940
rect 21218 16770 21678 16940
rect 21918 16770 22378 16940
rect 22618 16770 23078 16940
rect 23318 16770 23778 16940
rect 24018 16770 24478 16940
rect 24718 16770 25178 16940
rect 25418 16770 25878 16940
rect 18778 16760 18878 16770
rect 18778 16680 18788 16760
rect 18868 16680 18878 16760
rect 18778 16670 18878 16680
rect 19118 16670 25878 16770
rect 19118 16480 19578 16670
rect 19818 16480 20278 16670
rect 20518 16480 20978 16670
rect 21218 16480 21678 16670
rect 21918 16480 22378 16670
rect 22618 16480 23078 16670
rect 23318 16480 23778 16670
rect 24018 16480 24478 16670
rect 24718 16480 25178 16670
rect 25418 16480 25878 16670
rect 19118 16070 19578 16240
rect 19818 16070 20278 16240
rect 20518 16070 20978 16240
rect 21218 16070 21678 16240
rect 21918 16070 22378 16240
rect 22618 16070 23078 16240
rect 23318 16070 23778 16240
rect 24018 16070 24478 16240
rect 24718 16070 25178 16240
rect 25418 16070 25878 16240
rect 19118 16060 25878 16070
rect 18988 16050 25878 16060
rect 18988 15990 18998 16050
rect 19058 15990 25878 16050
rect 18988 15980 25878 15990
rect 19118 15970 25878 15980
rect 19118 15780 19578 15970
rect 19818 15780 20278 15970
rect 20518 15780 20978 15970
rect 21218 15780 21678 15970
rect 21918 15780 22378 15970
rect 22618 15780 23078 15970
rect 23318 15780 23778 15970
rect 24018 15780 24478 15970
rect 24718 15780 25178 15970
rect 25418 15780 25878 15970
rect 25598 15540 25698 15780
rect 19118 15370 19578 15540
rect 19818 15370 20278 15540
rect 20518 15370 20978 15540
rect 21218 15370 21678 15540
rect 21918 15370 22378 15540
rect 22618 15370 23078 15540
rect 23318 15370 23778 15540
rect 24018 15370 24478 15540
rect 24718 15370 25178 15540
rect 25418 15370 25878 15540
rect 18778 15360 18878 15370
rect 18778 15280 18788 15360
rect 18868 15280 18878 15360
rect 18778 15270 18878 15280
rect 19118 15270 25878 15370
rect 19118 15080 19578 15270
rect 19818 15080 20278 15270
rect 20518 15080 20978 15270
rect 21218 15080 21678 15270
rect 21918 15080 22378 15270
rect 22618 15080 23078 15270
rect 23318 15080 23778 15270
rect 24018 15080 24478 15270
rect 24718 15080 25178 15270
rect 25418 15080 25878 15270
rect 18338 14210 18578 14260
rect 18338 14150 18378 14210
rect 18438 14150 18478 14210
rect 18538 14150 18578 14210
rect 18338 13900 18578 14150
rect 18338 13840 18378 13900
rect 18438 13840 18478 13900
rect 18538 13840 18578 13900
rect 18338 13800 18578 13840
rect 18338 13740 18378 13800
rect 18438 13740 18478 13800
rect 18538 13740 18578 13800
rect 18038 13420 18278 13440
rect 18038 13360 18078 13420
rect 18138 13360 18178 13420
rect 18238 13360 18278 13420
rect 18038 13100 18278 13360
rect 18038 13040 18078 13100
rect 18138 13040 18178 13100
rect 18238 13040 18278 13100
rect 18038 13000 18278 13040
rect 18038 12940 18078 13000
rect 18138 12940 18178 13000
rect 18238 12940 18278 13000
rect 18038 11990 18278 12940
rect 18038 11930 18078 11990
rect 18138 11930 18178 11990
rect 18238 11930 18278 11990
rect 18038 11440 18278 11930
rect 18038 11380 18078 11440
rect 18138 11380 18178 11440
rect 18238 11380 18278 11440
rect 18038 11340 18278 11380
rect 18038 11280 18078 11340
rect 18138 11280 18178 11340
rect 18238 11280 18278 11340
rect 18038 9990 18278 11280
rect 18038 9930 18078 9990
rect 18138 9930 18178 9990
rect 18238 9930 18278 9990
rect 18038 9890 18278 9930
rect 18038 9830 18078 9890
rect 18138 9830 18178 9890
rect 18238 9830 18278 9890
rect 18038 9420 18278 9830
rect 18038 9360 18078 9420
rect 18138 9360 18178 9420
rect 18238 9360 18278 9420
rect 18038 9040 18278 9360
rect 198 9010 18278 9040
rect 198 8930 208 9010
rect 288 8930 308 9010
rect 388 8930 408 9010
rect 488 8930 508 9010
rect 588 8930 18278 9010
rect 198 8910 18278 8930
rect 198 8830 208 8910
rect 288 8830 308 8910
rect 388 8830 408 8910
rect 488 8830 508 8910
rect 588 8830 18278 8910
rect 198 8800 18278 8830
rect 18338 13180 18578 13740
rect 23208 13520 23308 13530
rect 23208 13510 25848 13520
rect 23208 13450 23228 13510
rect 23288 13450 25848 13510
rect 23208 13430 25848 13450
rect 18338 13120 18378 13180
rect 18438 13120 18478 13180
rect 18538 13120 18578 13180
rect 18338 10770 18578 13120
rect 23438 11580 23548 11600
rect 23438 11510 23458 11580
rect 23528 11510 23548 11580
rect 23438 11490 23548 11510
rect 23788 11460 25848 13430
rect 23438 11070 23548 11090
rect 23438 11000 23458 11070
rect 23528 11000 23548 11070
rect 23438 10980 23548 11000
rect 18338 10710 18378 10770
rect 18438 10710 18478 10770
rect 18538 10710 18578 10770
rect 18338 9650 18578 10710
rect 18338 9590 18378 9650
rect 18438 9590 18478 9650
rect 18538 9590 18578 9650
rect 18338 8740 18578 9590
rect 23788 9150 25848 11120
rect 23208 9130 25848 9150
rect 23208 9070 23228 9130
rect 23288 9070 25848 9130
rect 23208 9060 25848 9070
rect 23208 9050 23308 9060
rect 798 8710 18578 8740
rect 798 8630 808 8710
rect 888 8630 908 8710
rect 988 8630 1008 8710
rect 1088 8630 1108 8710
rect 1188 8630 18578 8710
rect 798 8610 18578 8630
rect 798 8530 808 8610
rect 888 8530 908 8610
rect 988 8530 1008 8610
rect 1088 8530 1108 8610
rect 1188 8530 18578 8610
rect 798 8500 18578 8530
rect 798 8360 13008 8390
rect 798 8280 808 8360
rect 888 8280 908 8360
rect 988 8280 1008 8360
rect 1088 8280 1108 8360
rect 1188 8350 13008 8360
rect 1188 8290 12928 8350
rect 12988 8290 13008 8350
rect 1188 8280 13008 8290
rect 798 8260 13008 8280
rect 798 8180 808 8260
rect 888 8180 908 8260
rect 988 8180 1008 8260
rect 1088 8180 1108 8260
rect 1188 8250 13008 8260
rect 1188 8190 12928 8250
rect 12988 8190 13008 8250
rect 1188 8180 13008 8190
rect 798 8150 13008 8180
rect 18338 8230 18578 8500
rect 18338 8170 18378 8230
rect 18438 8170 18478 8230
rect 18538 8170 18578 8230
rect 18338 8160 18578 8170
rect 23088 8380 23198 8400
rect 23088 8310 23108 8380
rect 23178 8310 23198 8380
rect 23088 8290 23198 8310
rect 22738 7590 22848 7610
rect 22738 7520 22758 7590
rect 22828 7520 22848 7590
rect 22738 7500 22848 7520
rect 23088 7470 23688 8290
rect 198 7180 13008 7210
rect 198 7100 208 7180
rect 288 7100 308 7180
rect 388 7100 408 7180
rect 488 7100 508 7180
rect 588 7170 13008 7180
rect 588 7110 12928 7170
rect 12988 7110 13008 7170
rect 588 7100 13008 7110
rect 198 7080 13008 7100
rect 198 7000 208 7080
rect 288 7000 308 7080
rect 388 7000 408 7080
rect 488 7000 508 7080
rect 588 7070 13008 7080
rect 588 7010 12928 7070
rect 12988 7010 13008 7070
rect 588 7000 13008 7010
rect 198 6970 13008 7000
rect 22738 7060 22848 7080
rect 22738 6990 22758 7060
rect 22828 6990 22848 7060
rect 22738 6970 22848 6990
rect 19238 6390 19478 6400
rect 19238 6330 19278 6390
rect 19338 6330 19378 6390
rect 19438 6330 19478 6390
rect 798 6000 13008 6030
rect 798 5920 808 6000
rect 888 5920 908 6000
rect 988 5920 1008 6000
rect 1088 5920 1108 6000
rect 1188 5990 13008 6000
rect 1188 5930 12928 5990
rect 12988 5930 13008 5990
rect 1188 5920 13008 5930
rect 798 5900 13008 5920
rect 798 5820 808 5900
rect 888 5820 908 5900
rect 988 5820 1008 5900
rect 1088 5820 1108 5900
rect 1188 5890 13008 5900
rect 1188 5830 12928 5890
rect 12988 5830 13008 5890
rect 1188 5820 13008 5830
rect 798 5790 13008 5820
rect 19238 5730 19478 6330
rect 23088 5900 24188 7110
rect 22978 5880 24188 5900
rect 22978 5810 22998 5880
rect 23068 5810 24188 5880
rect 22978 5790 24188 5810
rect 198 5700 22688 5730
rect 198 5620 208 5700
rect 288 5620 308 5700
rect 388 5620 408 5700
rect 488 5620 508 5700
rect 588 5690 22688 5700
rect 588 5630 22608 5690
rect 22668 5630 22688 5690
rect 588 5620 22688 5630
rect 198 5600 22688 5620
rect 198 5520 208 5600
rect 288 5520 308 5600
rect 388 5520 408 5600
rect 488 5520 508 5600
rect 588 5590 22688 5600
rect 588 5530 22608 5590
rect 22668 5530 22688 5590
rect 588 5520 22688 5530
rect 198 5490 22688 5520
rect 198 3800 12318 3830
rect 198 3720 208 3800
rect 288 3720 308 3800
rect 388 3720 408 3800
rect 488 3720 508 3800
rect 588 3790 12318 3800
rect 588 3730 12238 3790
rect 12298 3730 12318 3790
rect 588 3720 12318 3730
rect 198 3700 12318 3720
rect 198 3620 208 3700
rect 288 3620 308 3700
rect 388 3620 408 3700
rect 488 3620 508 3700
rect 588 3690 12318 3700
rect 588 3630 12238 3690
rect 12298 3630 12318 3690
rect 588 3620 12318 3630
rect 198 3590 12318 3620
rect 26508 3400 26668 3420
rect 26508 3320 26548 3400
rect 26628 3320 26668 3400
rect 26508 3280 26668 3320
rect 26508 3200 26548 3280
rect 26628 3200 26668 3280
rect 26508 3180 26668 3200
rect 798 3020 12318 3050
rect 798 2940 808 3020
rect 888 2940 908 3020
rect 988 2940 1008 3020
rect 1088 2940 1108 3020
rect 1188 3010 12318 3020
rect 1188 2950 12238 3010
rect 12298 2950 12318 3010
rect 1188 2940 12318 2950
rect 798 2920 12318 2940
rect 798 2840 808 2920
rect 888 2840 908 2920
rect 988 2840 1008 2920
rect 1088 2840 1108 2920
rect 1188 2910 12318 2920
rect 1188 2850 12238 2910
rect 12298 2850 12318 2910
rect 1188 2840 12318 2850
rect 798 2810 12318 2840
rect 798 1620 22688 1650
rect 798 1540 808 1620
rect 888 1540 908 1620
rect 988 1540 1008 1620
rect 1088 1540 1108 1620
rect 1188 1610 22688 1620
rect 1188 1550 22608 1610
rect 22668 1550 22688 1610
rect 1188 1540 22688 1550
rect 798 1520 22688 1540
rect 798 1440 808 1520
rect 888 1440 908 1520
rect 988 1440 1008 1520
rect 1088 1440 1108 1520
rect 1188 1510 22688 1520
rect 1188 1450 22608 1510
rect 22668 1450 22688 1510
rect 1188 1440 22688 1450
rect 798 1410 22688 1440
rect 30368 1340 30528 1380
rect 30368 1260 30408 1340
rect 30488 1260 30528 1340
rect 30368 1220 30528 1260
<< via3 >>
rect 808 19780 888 19860
rect 908 19780 988 19860
rect 1008 19780 1088 19860
rect 1108 19780 1188 19860
rect 808 19660 888 19740
rect 908 19660 988 19740
rect 1008 19660 1088 19740
rect 1108 19660 1188 19740
rect 22818 19720 22888 19790
rect 23318 19720 23388 19790
rect 808 18980 888 19060
rect 908 18980 988 19060
rect 1008 18980 1088 19060
rect 1108 18980 1188 19060
rect 808 18880 888 18960
rect 908 18880 988 18960
rect 1008 18880 1088 18960
rect 1108 18880 1188 18960
rect 18648 18150 18728 18160
rect 18648 18090 18658 18150
rect 18658 18090 18718 18150
rect 18718 18090 18728 18150
rect 18648 18080 18728 18090
rect 18788 16750 18868 16760
rect 18788 16690 18798 16750
rect 18798 16690 18858 16750
rect 18858 16690 18868 16750
rect 18788 16680 18868 16690
rect 18788 15350 18868 15360
rect 18788 15290 18798 15350
rect 18798 15290 18858 15350
rect 18858 15290 18868 15350
rect 18788 15280 18868 15290
rect 208 8930 288 9010
rect 308 8930 388 9010
rect 408 8930 488 9010
rect 508 8930 588 9010
rect 208 8830 288 8910
rect 308 8830 388 8910
rect 408 8830 488 8910
rect 508 8830 588 8910
rect 23458 11510 23528 11580
rect 23458 11000 23528 11070
rect 808 8630 888 8710
rect 908 8630 988 8710
rect 1008 8630 1088 8710
rect 1108 8630 1188 8710
rect 808 8530 888 8610
rect 908 8530 988 8610
rect 1008 8530 1088 8610
rect 1108 8530 1188 8610
rect 808 8280 888 8360
rect 908 8280 988 8360
rect 1008 8280 1088 8360
rect 1108 8280 1188 8360
rect 808 8180 888 8260
rect 908 8180 988 8260
rect 1008 8180 1088 8260
rect 1108 8180 1188 8260
rect 22758 7520 22828 7590
rect 208 7100 288 7180
rect 308 7100 388 7180
rect 408 7100 488 7180
rect 508 7100 588 7180
rect 208 7000 288 7080
rect 308 7000 388 7080
rect 408 7000 488 7080
rect 508 7000 588 7080
rect 22758 6990 22828 7060
rect 808 5920 888 6000
rect 908 5920 988 6000
rect 1008 5920 1088 6000
rect 1108 5920 1188 6000
rect 808 5820 888 5900
rect 908 5820 988 5900
rect 1008 5820 1088 5900
rect 1108 5820 1188 5900
rect 208 5620 288 5700
rect 308 5620 388 5700
rect 408 5620 488 5700
rect 508 5620 588 5700
rect 208 5520 288 5600
rect 308 5520 388 5600
rect 408 5520 488 5600
rect 508 5520 588 5600
rect 208 3720 288 3800
rect 308 3720 388 3800
rect 408 3720 488 3800
rect 508 3720 588 3800
rect 208 3620 288 3700
rect 308 3620 388 3700
rect 408 3620 488 3700
rect 508 3620 588 3700
rect 26548 3320 26628 3400
rect 26548 3200 26628 3280
rect 808 2940 888 3020
rect 908 2940 988 3020
rect 1008 2940 1088 3020
rect 1108 2940 1188 3020
rect 808 2840 888 2920
rect 908 2840 988 2920
rect 1008 2840 1088 2920
rect 1108 2840 1188 2920
rect 808 1540 888 1620
rect 908 1540 988 1620
rect 1008 1540 1088 1620
rect 1108 1540 1188 1620
rect 808 1440 888 1520
rect 908 1440 988 1520
rect 1008 1440 1088 1520
rect 1108 1440 1188 1520
rect 30408 1260 30488 1340
<< mimcap >>
rect 8948 20170 22908 32080
rect 8948 20100 22818 20170
rect 22888 20100 22908 20170
rect 8948 20080 22908 20100
rect 23298 20170 26058 32080
rect 23298 20100 23318 20170
rect 23388 20100 26058 20170
rect 23298 20080 26058 20100
rect 19148 18860 19548 19010
rect 19148 18780 19318 18860
rect 19398 18780 19548 18860
rect 19148 18610 19548 18780
rect 19848 18860 20248 19010
rect 19848 18780 20008 18860
rect 20088 18780 20248 18860
rect 19848 18610 20248 18780
rect 20548 18860 20948 19010
rect 20548 18780 20708 18860
rect 20788 18780 20948 18860
rect 20548 18610 20948 18780
rect 21248 18860 21648 19010
rect 21248 18780 21408 18860
rect 21488 18780 21648 18860
rect 21248 18610 21648 18780
rect 21948 18860 22348 19010
rect 21948 18780 22108 18860
rect 22188 18780 22348 18860
rect 21948 18610 22348 18780
rect 22648 18860 23048 19010
rect 22648 18780 22808 18860
rect 22888 18780 23048 18860
rect 22648 18610 23048 18780
rect 23348 18860 23748 19010
rect 23348 18780 23508 18860
rect 23588 18780 23748 18860
rect 23348 18610 23748 18780
rect 24048 18860 24448 19010
rect 24048 18780 24208 18860
rect 24288 18780 24448 18860
rect 24048 18610 24448 18780
rect 24748 18860 25148 19010
rect 24748 18780 24908 18860
rect 24988 18780 25148 18860
rect 24748 18610 25148 18780
rect 25448 18860 25848 19010
rect 25448 18780 25608 18860
rect 25688 18780 25848 18860
rect 25448 18610 25848 18780
rect 19148 18160 19548 18310
rect 19148 18080 19318 18160
rect 19398 18080 19548 18160
rect 19148 17910 19548 18080
rect 19848 18160 20248 18310
rect 19848 18080 20008 18160
rect 20088 18080 20248 18160
rect 19848 17910 20248 18080
rect 20548 18160 20948 18310
rect 20548 18080 20708 18160
rect 20788 18080 20948 18160
rect 20548 17910 20948 18080
rect 21248 18160 21648 18310
rect 21248 18080 21408 18160
rect 21488 18080 21648 18160
rect 21248 17910 21648 18080
rect 21948 18160 22348 18310
rect 21948 18080 22108 18160
rect 22188 18080 22348 18160
rect 21948 17910 22348 18080
rect 22648 18160 23048 18310
rect 22648 18080 22808 18160
rect 22888 18080 23048 18160
rect 22648 17910 23048 18080
rect 23348 18160 23748 18310
rect 23348 18080 23508 18160
rect 23588 18080 23748 18160
rect 23348 17910 23748 18080
rect 24048 18160 24448 18310
rect 24048 18080 24208 18160
rect 24288 18080 24448 18160
rect 24048 17910 24448 18080
rect 24748 18160 25148 18310
rect 24748 18080 24908 18160
rect 24988 18080 25148 18160
rect 24748 17910 25148 18080
rect 25448 18160 25848 18310
rect 25448 18080 25608 18160
rect 25688 18080 25848 18160
rect 25448 17910 25848 18080
rect 19148 17460 19548 17610
rect 19148 17380 19318 17460
rect 19398 17380 19548 17460
rect 19148 17210 19548 17380
rect 19848 17460 20248 17610
rect 19848 17380 20008 17460
rect 20088 17380 20248 17460
rect 19848 17210 20248 17380
rect 20548 17460 20948 17610
rect 20548 17380 20708 17460
rect 20788 17380 20948 17460
rect 20548 17210 20948 17380
rect 21248 17460 21648 17610
rect 21248 17380 21408 17460
rect 21488 17380 21648 17460
rect 21248 17210 21648 17380
rect 21948 17460 22348 17610
rect 21948 17380 22108 17460
rect 22188 17380 22348 17460
rect 21948 17210 22348 17380
rect 22648 17460 23048 17610
rect 22648 17380 22808 17460
rect 22888 17380 23048 17460
rect 22648 17210 23048 17380
rect 23348 17460 23748 17610
rect 23348 17380 23508 17460
rect 23588 17380 23748 17460
rect 23348 17210 23748 17380
rect 24048 17460 24448 17610
rect 24048 17380 24208 17460
rect 24288 17380 24448 17460
rect 24048 17210 24448 17380
rect 24748 17460 25148 17610
rect 24748 17380 24908 17460
rect 24988 17380 25148 17460
rect 24748 17210 25148 17380
rect 25448 17460 25848 17610
rect 25448 17380 25608 17460
rect 25688 17380 25848 17460
rect 25448 17210 25848 17380
rect 19148 16760 19548 16910
rect 19148 16680 19318 16760
rect 19398 16680 19548 16760
rect 19148 16510 19548 16680
rect 19848 16760 20248 16910
rect 19848 16680 20008 16760
rect 20088 16680 20248 16760
rect 19848 16510 20248 16680
rect 20548 16760 20948 16910
rect 20548 16680 20708 16760
rect 20788 16680 20948 16760
rect 20548 16510 20948 16680
rect 21248 16760 21648 16910
rect 21248 16680 21408 16760
rect 21488 16680 21648 16760
rect 21248 16510 21648 16680
rect 21948 16760 22348 16910
rect 21948 16680 22108 16760
rect 22188 16680 22348 16760
rect 21948 16510 22348 16680
rect 22648 16760 23048 16910
rect 22648 16680 22808 16760
rect 22888 16680 23048 16760
rect 22648 16510 23048 16680
rect 23348 16760 23748 16910
rect 23348 16680 23508 16760
rect 23588 16680 23748 16760
rect 23348 16510 23748 16680
rect 24048 16760 24448 16910
rect 24048 16680 24208 16760
rect 24288 16680 24448 16760
rect 24048 16510 24448 16680
rect 24748 16760 25148 16910
rect 24748 16680 24908 16760
rect 24988 16680 25148 16760
rect 24748 16510 25148 16680
rect 25448 16760 25848 16910
rect 25448 16680 25608 16760
rect 25688 16680 25848 16760
rect 25448 16510 25848 16680
rect 19148 16060 19548 16210
rect 19148 15980 19318 16060
rect 19398 15980 19548 16060
rect 19148 15810 19548 15980
rect 19848 16060 20248 16210
rect 19848 15980 20008 16060
rect 20088 15980 20248 16060
rect 19848 15810 20248 15980
rect 20548 16060 20948 16210
rect 20548 15980 20708 16060
rect 20788 15980 20948 16060
rect 20548 15810 20948 15980
rect 21248 16060 21648 16210
rect 21248 15980 21408 16060
rect 21488 15980 21648 16060
rect 21248 15810 21648 15980
rect 21948 16060 22348 16210
rect 21948 15980 22108 16060
rect 22188 15980 22348 16060
rect 21948 15810 22348 15980
rect 22648 16060 23048 16210
rect 22648 15980 22808 16060
rect 22888 15980 23048 16060
rect 22648 15810 23048 15980
rect 23348 16060 23748 16210
rect 23348 15980 23508 16060
rect 23588 15980 23748 16060
rect 23348 15810 23748 15980
rect 24048 16060 24448 16210
rect 24048 15980 24208 16060
rect 24288 15980 24448 16060
rect 24048 15810 24448 15980
rect 24748 16060 25148 16210
rect 24748 15980 24908 16060
rect 24988 15980 25148 16060
rect 24748 15810 25148 15980
rect 25448 16060 25848 16210
rect 25448 15980 25608 16060
rect 25688 15980 25848 16060
rect 25448 15810 25848 15980
rect 19148 15360 19548 15510
rect 19148 15280 19318 15360
rect 19398 15280 19548 15360
rect 19148 15110 19548 15280
rect 19848 15360 20248 15510
rect 19848 15280 20008 15360
rect 20088 15280 20248 15360
rect 19848 15110 20248 15280
rect 20548 15360 20948 15510
rect 20548 15280 20708 15360
rect 20788 15280 20948 15360
rect 20548 15110 20948 15280
rect 21248 15360 21648 15510
rect 21248 15280 21408 15360
rect 21488 15280 21648 15360
rect 21248 15110 21648 15280
rect 21948 15360 22348 15510
rect 21948 15280 22108 15360
rect 22188 15280 22348 15360
rect 21948 15110 22348 15280
rect 22648 15360 23048 15510
rect 22648 15280 22808 15360
rect 22888 15280 23048 15360
rect 22648 15110 23048 15280
rect 23348 15360 23748 15510
rect 23348 15280 23508 15360
rect 23588 15280 23748 15360
rect 23348 15110 23748 15280
rect 24048 15360 24448 15510
rect 24048 15280 24208 15360
rect 24288 15280 24448 15360
rect 24048 15110 24448 15280
rect 24748 15360 25148 15510
rect 24748 15280 24908 15360
rect 24988 15280 25148 15360
rect 24748 15110 25148 15280
rect 25448 15360 25848 15510
rect 25448 15280 25608 15360
rect 25688 15280 25848 15360
rect 25448 15110 25848 15280
rect 23818 11580 25818 13490
rect 23818 11510 23838 11580
rect 23908 11510 25818 11580
rect 23818 11490 25818 11510
rect 23818 11070 25818 11090
rect 23818 11000 23838 11070
rect 23908 11000 25818 11070
rect 23818 9090 25818 11000
rect 23118 7590 23658 8260
rect 23118 7520 23138 7590
rect 23208 7520 23658 7590
rect 23118 7500 23658 7520
rect 23118 7060 24158 7080
rect 23118 6990 23138 7060
rect 23208 6990 24158 7060
rect 23118 5820 24158 6990
<< mimcapcontact >>
rect 22818 20100 22888 20170
rect 23318 20100 23388 20170
rect 19318 18780 19398 18860
rect 20008 18780 20088 18860
rect 20708 18780 20788 18860
rect 21408 18780 21488 18860
rect 22108 18780 22188 18860
rect 22808 18780 22888 18860
rect 23508 18780 23588 18860
rect 24208 18780 24288 18860
rect 24908 18780 24988 18860
rect 25608 18780 25688 18860
rect 19318 18080 19398 18160
rect 20008 18080 20088 18160
rect 20708 18080 20788 18160
rect 21408 18080 21488 18160
rect 22108 18080 22188 18160
rect 22808 18080 22888 18160
rect 23508 18080 23588 18160
rect 24208 18080 24288 18160
rect 24908 18080 24988 18160
rect 25608 18080 25688 18160
rect 19318 17380 19398 17460
rect 20008 17380 20088 17460
rect 20708 17380 20788 17460
rect 21408 17380 21488 17460
rect 22108 17380 22188 17460
rect 22808 17380 22888 17460
rect 23508 17380 23588 17460
rect 24208 17380 24288 17460
rect 24908 17380 24988 17460
rect 25608 17380 25688 17460
rect 19318 16680 19398 16760
rect 20008 16680 20088 16760
rect 20708 16680 20788 16760
rect 21408 16680 21488 16760
rect 22108 16680 22188 16760
rect 22808 16680 22888 16760
rect 23508 16680 23588 16760
rect 24208 16680 24288 16760
rect 24908 16680 24988 16760
rect 25608 16680 25688 16760
rect 19318 15980 19398 16060
rect 20008 15980 20088 16060
rect 20708 15980 20788 16060
rect 21408 15980 21488 16060
rect 22108 15980 22188 16060
rect 22808 15980 22888 16060
rect 23508 15980 23588 16060
rect 24208 15980 24288 16060
rect 24908 15980 24988 16060
rect 25608 15980 25688 16060
rect 19318 15280 19398 15360
rect 20008 15280 20088 15360
rect 20708 15280 20788 15360
rect 21408 15280 21488 15360
rect 22108 15280 22188 15360
rect 22808 15280 22888 15360
rect 23508 15280 23588 15360
rect 24208 15280 24288 15360
rect 24908 15280 24988 15360
rect 25608 15280 25688 15360
rect 23838 11510 23908 11580
rect 23838 11000 23908 11070
rect 23138 7520 23208 7590
rect 23138 6990 23208 7060
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 9040 600 44152
rect 800 19890 1200 44152
rect 798 19860 1200 19890
rect 798 19780 808 19860
rect 888 19780 908 19860
rect 988 19780 1008 19860
rect 1088 19780 1108 19860
rect 1188 19780 1200 19860
rect 798 19740 1200 19780
rect 798 19660 808 19740
rect 888 19660 908 19740
rect 988 19660 1008 19740
rect 1088 19660 1108 19740
rect 1188 19660 1200 19740
rect 22798 20170 22908 20180
rect 22798 20100 22818 20170
rect 22888 20100 22908 20170
rect 22798 19790 22908 20100
rect 22798 19720 22818 19790
rect 22888 19720 22908 19790
rect 22798 19700 22908 19720
rect 23298 20170 23408 20180
rect 23298 20100 23318 20170
rect 23388 20100 23408 20170
rect 23298 19790 23408 20100
rect 23298 19720 23318 19790
rect 23388 19720 23408 19790
rect 23298 19700 23408 19720
rect 798 19630 1200 19660
rect 800 19090 1200 19630
rect 798 19060 1200 19090
rect 798 18980 808 19060
rect 888 18980 908 19060
rect 988 18980 1008 19060
rect 1088 18980 1108 19060
rect 1188 18980 1200 19060
rect 798 18960 1200 18980
rect 798 18880 808 18960
rect 888 18880 908 18960
rect 988 18880 1008 18960
rect 1088 18880 1108 18960
rect 1188 18880 1200 18960
rect 798 18850 1200 18880
rect 800 9040 1200 18850
rect 19308 18860 25698 18870
rect 19308 18780 19318 18860
rect 19398 18780 20008 18860
rect 20088 18780 20708 18860
rect 20788 18780 21408 18860
rect 21488 18780 22108 18860
rect 22188 18780 22808 18860
rect 22888 18780 23508 18860
rect 23588 18780 24208 18860
rect 24288 18780 24908 18860
rect 24988 18780 25608 18860
rect 25688 18780 25698 18860
rect 19308 18770 25698 18780
rect 25598 18170 25698 18770
rect 18638 18160 25698 18170
rect 18638 18080 18648 18160
rect 18728 18080 19318 18160
rect 19398 18080 20008 18160
rect 20088 18080 20708 18160
rect 20788 18080 21408 18160
rect 21488 18080 22108 18160
rect 22188 18080 22808 18160
rect 22888 18080 23508 18160
rect 23588 18080 24208 18160
rect 24288 18080 24908 18160
rect 24988 18080 25608 18160
rect 25688 18080 25698 18160
rect 18638 18070 25698 18080
rect 19308 17460 25698 17470
rect 19308 17380 19318 17460
rect 19398 17380 20008 17460
rect 20088 17380 20708 17460
rect 20788 17380 21408 17460
rect 21488 17380 22108 17460
rect 22188 17380 22808 17460
rect 22888 17380 23508 17460
rect 23588 17380 24208 17460
rect 24288 17380 24908 17460
rect 24988 17380 25608 17460
rect 25688 17380 25698 17460
rect 19308 17370 25698 17380
rect 25598 16770 25698 17370
rect 18778 16760 25698 16770
rect 18778 16680 18788 16760
rect 18868 16680 19318 16760
rect 19398 16680 20008 16760
rect 20088 16680 20708 16760
rect 20788 16680 21408 16760
rect 21488 16680 22108 16760
rect 22188 16680 22808 16760
rect 22888 16680 23508 16760
rect 23588 16680 24208 16760
rect 24288 16680 24908 16760
rect 24988 16680 25608 16760
rect 25688 16680 25698 16760
rect 18778 16670 25698 16680
rect 19308 16060 25698 16070
rect 19308 15980 19318 16060
rect 19398 15980 20008 16060
rect 20088 15980 20708 16060
rect 20788 15980 21408 16060
rect 21488 15980 22108 16060
rect 22188 15980 22808 16060
rect 22888 15980 23508 16060
rect 23588 15980 24208 16060
rect 24288 15980 24908 16060
rect 24988 15980 25608 16060
rect 25688 15980 25698 16060
rect 19308 15970 25698 15980
rect 25598 15370 25698 15970
rect 18778 15360 25698 15370
rect 18778 15280 18788 15360
rect 18868 15280 19318 15360
rect 19398 15280 20008 15360
rect 20088 15280 20708 15360
rect 20788 15280 21408 15360
rect 21488 15280 22108 15360
rect 22188 15280 22808 15360
rect 22888 15280 23508 15360
rect 23588 15280 24208 15360
rect 24288 15280 24908 15360
rect 24988 15280 25608 15360
rect 25688 15280 25698 15360
rect 18778 15270 25698 15280
rect 23438 11580 23918 11600
rect 23438 11510 23458 11580
rect 23528 11510 23838 11580
rect 23908 11510 23918 11580
rect 23438 11490 23918 11510
rect 23438 11070 23918 11090
rect 23438 11000 23458 11070
rect 23528 11000 23838 11070
rect 23908 11000 23918 11070
rect 23438 10980 23918 11000
rect 198 9010 600 9040
rect 198 8930 208 9010
rect 288 8930 308 9010
rect 388 8930 408 9010
rect 488 8930 508 9010
rect 588 8930 600 9010
rect 198 8910 600 8930
rect 198 8830 208 8910
rect 288 8830 308 8910
rect 388 8830 408 8910
rect 488 8830 508 8910
rect 588 8830 600 8910
rect 198 8800 600 8830
rect 798 8800 1200 9040
rect 200 7210 600 8800
rect 800 8740 1200 8800
rect 798 8710 1200 8740
rect 798 8630 808 8710
rect 888 8630 908 8710
rect 988 8630 1008 8710
rect 1088 8630 1108 8710
rect 1188 8630 1200 8710
rect 798 8610 1200 8630
rect 798 8530 808 8610
rect 888 8530 908 8610
rect 988 8530 1008 8610
rect 1088 8530 1108 8610
rect 1188 8530 1200 8610
rect 798 8500 1200 8530
rect 800 8390 1200 8500
rect 798 8360 1200 8390
rect 798 8280 808 8360
rect 888 8280 908 8360
rect 988 8280 1008 8360
rect 1088 8280 1108 8360
rect 1188 8280 1200 8360
rect 798 8260 1200 8280
rect 798 8180 808 8260
rect 888 8180 908 8260
rect 988 8180 1008 8260
rect 1088 8180 1108 8260
rect 1188 8180 1200 8260
rect 798 8150 1200 8180
rect 800 7210 1200 8150
rect 22738 7590 23228 7610
rect 22738 7520 22758 7590
rect 22828 7520 23138 7590
rect 23208 7520 23228 7590
rect 22738 7500 23228 7520
rect 198 7180 600 7210
rect 198 7100 208 7180
rect 288 7100 308 7180
rect 388 7100 408 7180
rect 488 7100 508 7180
rect 588 7100 600 7180
rect 198 7080 600 7100
rect 198 7000 208 7080
rect 288 7000 308 7080
rect 388 7000 408 7080
rect 488 7000 508 7080
rect 588 7000 600 7080
rect 198 6970 600 7000
rect 798 6970 1200 7210
rect 22738 7060 23228 7080
rect 22738 6990 22758 7060
rect 22828 6990 23138 7060
rect 23208 6990 23228 7060
rect 22738 6970 23228 6990
rect 200 5730 600 6970
rect 800 6030 1200 6970
rect 798 6000 1200 6030
rect 798 5920 808 6000
rect 888 5920 908 6000
rect 988 5920 1008 6000
rect 1088 5920 1108 6000
rect 1188 5920 1200 6000
rect 798 5900 1200 5920
rect 798 5820 808 5900
rect 888 5820 908 5900
rect 988 5820 1008 5900
rect 1088 5820 1108 5900
rect 1188 5820 1200 5900
rect 798 5790 1200 5820
rect 800 5730 1200 5790
rect 198 5700 600 5730
rect 198 5620 208 5700
rect 288 5620 308 5700
rect 388 5620 408 5700
rect 488 5620 508 5700
rect 588 5620 600 5700
rect 198 5600 600 5620
rect 198 5520 208 5600
rect 288 5520 308 5600
rect 388 5520 408 5600
rect 488 5520 508 5600
rect 588 5520 600 5600
rect 198 5490 600 5520
rect 798 5490 1200 5730
rect 200 3830 600 5490
rect 800 3830 1200 5490
rect 198 3800 600 3830
rect 198 3720 208 3800
rect 288 3720 308 3800
rect 388 3720 408 3800
rect 488 3720 508 3800
rect 588 3720 600 3800
rect 198 3700 600 3720
rect 198 3620 208 3700
rect 288 3620 308 3700
rect 388 3620 408 3700
rect 488 3620 508 3700
rect 588 3620 600 3700
rect 198 3590 600 3620
rect 798 3590 1200 3830
rect 200 1000 600 3590
rect 800 3050 1200 3590
rect 798 3020 1200 3050
rect 798 2940 808 3020
rect 888 2940 908 3020
rect 988 2940 1008 3020
rect 1088 2940 1108 3020
rect 1188 2940 1200 3020
rect 798 2920 1200 2940
rect 798 2840 808 2920
rect 888 2840 908 2920
rect 988 2840 1008 2920
rect 1088 2840 1108 2920
rect 1188 2840 1200 2920
rect 798 2810 1200 2840
rect 800 1650 1200 2810
rect 798 1620 1200 1650
rect 798 1540 808 1620
rect 888 1540 908 1620
rect 988 1540 1008 1620
rect 1088 1540 1108 1620
rect 1188 1540 1200 1620
rect 798 1520 1200 1540
rect 798 1440 808 1520
rect 888 1440 908 1520
rect 988 1440 1008 1520
rect 1088 1440 1108 1520
rect 1188 1440 1200 1520
rect 798 1410 1200 1440
rect 800 1000 1200 1410
rect 26508 3400 26668 3420
rect 26508 3320 26548 3400
rect 26628 3320 26668 3400
rect 26508 3280 26668 3320
rect 26508 3200 26548 3280
rect 26628 3200 26668 3280
rect 26508 200 26668 3200
rect 30368 1340 30528 1380
rect 30368 1260 30408 1340
rect 30488 1260 30528 1340
rect 30368 200 30528 1260
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal1 26078 2390 26078 2390 3 FreeSans 1600 0 800 0 V_CONT
flabel metal1 18648 7760 18648 7760 7 FreeSans 1600 0 -800 0 I_IN
flabel metal2 13288 9690 13288 9690 5 FreeSans 1600 0 0 -800 PFET_GATE
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
