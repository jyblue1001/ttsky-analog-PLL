magic
tech sky130A
magscale 1 2
timestamp 1757393620
<< nwell >>
rect 38567 16457 39091 18625
rect 39347 14887 39871 18631
rect 40127 16111 40983 18633
rect 45447 16111 46303 18633
rect 46557 15777 47081 18631
rect 47347 16457 47871 18625
rect 41367 14117 45189 14641
rect 40400 11180 43130 11460
rect 43430 11180 46160 11460
rect 41500 9620 45060 10300
rect 45360 9820 46130 10100
rect 41510 9020 43150 9300
rect 43410 9020 45050 9300
<< pwell >>
rect 43240 18810 43320 19090
rect 41250 18657 42590 18810
rect 41250 17623 41403 18657
rect 42437 17623 42590 18657
rect 41250 17470 42590 17623
rect 42610 18657 43950 18810
rect 42610 17623 42763 18657
rect 43797 17623 43950 18657
rect 42610 17470 43950 17623
rect 43970 18657 45310 18810
rect 43970 17623 44123 18657
rect 45157 17623 45310 18657
rect 43970 17470 45310 17623
rect 41250 17297 42590 17450
rect 41250 16263 41403 17297
rect 42437 16263 42590 17297
rect 41250 16110 42590 16263
rect 42610 17297 43950 17450
rect 42610 16263 42763 17297
rect 43797 16263 43950 17297
rect 42610 16110 43950 16263
rect 43970 17297 45310 17450
rect 43970 16263 44123 17297
rect 45157 16263 45310 17297
rect 43970 16110 45310 16263
rect 41250 15937 42590 16090
rect 41250 14903 41403 15937
rect 42437 14903 42590 15937
rect 41250 14750 42590 14903
rect 42610 15937 43950 16090
rect 42610 14903 42763 15937
rect 43797 14903 43950 15937
rect 42610 14750 43950 14903
rect 43970 15937 45310 16090
rect 43970 14903 44123 15937
rect 45157 14903 45310 15937
rect 43970 14750 45310 14903
<< nbase >>
rect 41403 17623 42437 18657
rect 42763 17623 43797 18657
rect 44123 17623 45157 18657
rect 41403 16263 42437 17297
rect 42763 16263 43797 17297
rect 44123 16263 45157 17297
rect 41403 14903 42437 15937
rect 42763 14903 43797 15937
rect 44123 14903 45157 15937
<< nmos >>
rect 41240 13680 43240 13880
rect 43320 13680 45320 13880
rect 40820 12770 41820 13270
rect 42060 12770 43060 13270
rect 43500 12770 44500 13270
rect 44740 12770 45740 13270
rect 41440 12160 41480 12260
rect 41560 12160 41600 12260
rect 41680 12160 41720 12260
rect 41800 12160 41840 12260
rect 41920 12160 41960 12260
rect 42040 12160 42080 12260
rect 42160 12160 42200 12260
rect 42280 12160 42320 12260
rect 42400 12160 42440 12260
rect 42520 12160 42560 12260
rect 44000 12160 44040 12260
rect 44120 12160 44160 12260
rect 44240 12160 44280 12260
rect 44360 12160 44400 12260
rect 44480 12160 44520 12260
rect 44600 12160 44640 12260
rect 44720 12160 44760 12260
rect 44840 12160 44880 12260
rect 44960 12160 45000 12260
rect 45080 12160 45120 12260
<< pmos >>
rect 40600 11220 40640 11420
rect 40720 11220 40760 11420
rect 40840 11220 40880 11420
rect 40960 11220 41000 11420
rect 41080 11220 41120 11420
rect 41200 11220 41240 11420
rect 41320 11220 41360 11420
rect 41440 11220 41480 11420
rect 41560 11220 41600 11420
rect 41680 11220 41720 11420
rect 41800 11220 41840 11420
rect 41920 11220 41960 11420
rect 42040 11220 42080 11420
rect 42160 11220 42200 11420
rect 42280 11220 42320 11420
rect 42400 11220 42440 11420
rect 42520 11220 42560 11420
rect 42640 11220 42680 11420
rect 42760 11220 42800 11420
rect 42880 11220 42920 11420
rect 43640 11220 43680 11420
rect 43760 11220 43800 11420
rect 43880 11220 43920 11420
rect 44000 11220 44040 11420
rect 44120 11220 44160 11420
rect 44240 11220 44280 11420
rect 44360 11220 44400 11420
rect 44480 11220 44520 11420
rect 44600 11220 44640 11420
rect 44720 11220 44760 11420
rect 44840 11220 44880 11420
rect 44960 11220 45000 11420
rect 45080 11220 45120 11420
rect 45200 11220 45240 11420
rect 45320 11220 45360 11420
rect 45440 11220 45480 11420
rect 45560 11220 45600 11420
rect 45680 11220 45720 11420
rect 45800 11220 45840 11420
rect 45920 11220 45960 11420
rect 41700 9660 41800 10260
rect 41880 9660 41980 10260
rect 42060 9660 42160 10260
rect 42240 9660 42340 10260
rect 42420 9660 42520 10260
rect 42600 9660 42700 10260
rect 42780 9660 42880 10260
rect 42960 9660 43060 10260
rect 43140 9660 43240 10260
rect 43320 9660 43420 10260
rect 43500 9660 43600 10260
rect 43680 9660 43780 10260
rect 43860 9660 43960 10260
rect 44040 9660 44140 10260
rect 44220 9660 44320 10260
rect 44400 9660 44500 10260
rect 44580 9660 44680 10260
rect 44760 9660 44860 10260
rect 45570 9860 45600 10060
rect 45680 9860 45710 10060
rect 45790 9860 45820 10060
rect 45900 9860 45930 10060
rect 41710 9060 41740 9260
rect 41820 9060 41850 9260
rect 41930 9060 41960 9260
rect 42040 9060 42070 9260
rect 42150 9060 42180 9260
rect 42260 9060 42290 9260
rect 42370 9060 42400 9260
rect 42480 9060 42510 9260
rect 42590 9060 42620 9260
rect 42700 9060 42730 9260
rect 42810 9060 42840 9260
rect 42920 9060 42950 9260
rect 43610 9060 43640 9260
rect 43720 9060 43750 9260
rect 43830 9060 43860 9260
rect 43940 9060 43970 9260
rect 44050 9060 44080 9260
rect 44160 9060 44190 9260
rect 44270 9060 44300 9260
rect 44380 9060 44410 9260
rect 44490 9060 44520 9260
rect 44600 9060 44630 9260
rect 44710 9060 44740 9260
rect 44820 9060 44850 9260
<< ndiff >>
rect 41160 13850 41240 13880
rect 41160 13810 41180 13850
rect 41220 13810 41240 13850
rect 41160 13750 41240 13810
rect 41160 13710 41180 13750
rect 41220 13710 41240 13750
rect 41160 13680 41240 13710
rect 43240 13850 43320 13880
rect 43240 13810 43260 13850
rect 43300 13810 43320 13850
rect 43240 13750 43320 13810
rect 43240 13710 43260 13750
rect 43300 13710 43320 13750
rect 43240 13680 43320 13710
rect 45320 13850 45400 13880
rect 45320 13810 45340 13850
rect 45380 13810 45400 13850
rect 45320 13750 45400 13810
rect 45320 13710 45340 13750
rect 45380 13710 45400 13750
rect 45320 13680 45400 13710
rect 40740 13240 40820 13270
rect 40740 13200 40760 13240
rect 40800 13200 40820 13240
rect 40740 13140 40820 13200
rect 40740 13100 40760 13140
rect 40800 13100 40820 13140
rect 40740 13040 40820 13100
rect 40740 13000 40760 13040
rect 40800 13000 40820 13040
rect 40740 12940 40820 13000
rect 40740 12900 40760 12940
rect 40800 12900 40820 12940
rect 40740 12840 40820 12900
rect 40740 12800 40760 12840
rect 40800 12800 40820 12840
rect 40740 12770 40820 12800
rect 41820 13240 41900 13270
rect 41980 13240 42060 13270
rect 41820 13200 41840 13240
rect 41880 13200 41900 13240
rect 41980 13200 42000 13240
rect 42040 13200 42060 13240
rect 41820 13140 41900 13200
rect 41980 13140 42060 13200
rect 41820 13100 41840 13140
rect 41880 13100 41900 13140
rect 41980 13100 42000 13140
rect 42040 13100 42060 13140
rect 41820 13040 41900 13100
rect 41980 13040 42060 13100
rect 41820 13000 41840 13040
rect 41880 13000 41900 13040
rect 41980 13000 42000 13040
rect 42040 13000 42060 13040
rect 41820 12940 41900 13000
rect 41980 12940 42060 13000
rect 41820 12900 41840 12940
rect 41880 12900 41900 12940
rect 41980 12900 42000 12940
rect 42040 12900 42060 12940
rect 41820 12840 41900 12900
rect 41980 12840 42060 12900
rect 41820 12800 41840 12840
rect 41880 12800 41900 12840
rect 41980 12800 42000 12840
rect 42040 12800 42060 12840
rect 41820 12770 41900 12800
rect 41980 12770 42060 12800
rect 43060 13240 43140 13270
rect 43060 13200 43080 13240
rect 43120 13200 43140 13240
rect 43060 13140 43140 13200
rect 43060 13100 43080 13140
rect 43120 13100 43140 13140
rect 43060 13040 43140 13100
rect 43060 13000 43080 13040
rect 43120 13000 43140 13040
rect 43060 12940 43140 13000
rect 43060 12900 43080 12940
rect 43120 12900 43140 12940
rect 43060 12840 43140 12900
rect 43060 12800 43080 12840
rect 43120 12800 43140 12840
rect 43060 12770 43140 12800
rect 43420 13240 43500 13270
rect 43420 13200 43440 13240
rect 43480 13200 43500 13240
rect 43420 13140 43500 13200
rect 43420 13100 43440 13140
rect 43480 13100 43500 13140
rect 43420 13040 43500 13100
rect 43420 13000 43440 13040
rect 43480 13000 43500 13040
rect 43420 12940 43500 13000
rect 43420 12900 43440 12940
rect 43480 12900 43500 12940
rect 43420 12840 43500 12900
rect 43420 12800 43440 12840
rect 43480 12800 43500 12840
rect 43420 12770 43500 12800
rect 44500 13240 44580 13270
rect 44660 13240 44740 13270
rect 44500 13200 44520 13240
rect 44560 13200 44580 13240
rect 44660 13200 44680 13240
rect 44720 13200 44740 13240
rect 44500 13140 44580 13200
rect 44660 13140 44740 13200
rect 44500 13100 44520 13140
rect 44560 13100 44580 13140
rect 44660 13100 44680 13140
rect 44720 13100 44740 13140
rect 44500 13040 44580 13100
rect 44660 13040 44740 13100
rect 44500 13000 44520 13040
rect 44560 13000 44580 13040
rect 44660 13000 44680 13040
rect 44720 13000 44740 13040
rect 44500 12940 44580 13000
rect 44660 12940 44740 13000
rect 44500 12900 44520 12940
rect 44560 12900 44580 12940
rect 44660 12900 44680 12940
rect 44720 12900 44740 12940
rect 44500 12840 44580 12900
rect 44660 12840 44740 12900
rect 44500 12800 44520 12840
rect 44560 12800 44580 12840
rect 44660 12800 44680 12840
rect 44720 12800 44740 12840
rect 44500 12770 44580 12800
rect 44660 12770 44740 12800
rect 45740 13240 45820 13270
rect 45740 13200 45760 13240
rect 45800 13200 45820 13240
rect 45740 13140 45820 13200
rect 45740 13100 45760 13140
rect 45800 13100 45820 13140
rect 45740 13040 45820 13100
rect 45740 13000 45760 13040
rect 45800 13000 45820 13040
rect 45740 12940 45820 13000
rect 45740 12900 45760 12940
rect 45800 12900 45820 12940
rect 45740 12840 45820 12900
rect 45740 12800 45760 12840
rect 45800 12800 45820 12840
rect 45740 12770 45820 12800
rect 41360 12230 41440 12260
rect 41360 12190 41380 12230
rect 41420 12190 41440 12230
rect 41360 12160 41440 12190
rect 41480 12230 41560 12260
rect 41480 12190 41500 12230
rect 41540 12190 41560 12230
rect 41480 12160 41560 12190
rect 41600 12230 41680 12260
rect 41600 12190 41620 12230
rect 41660 12190 41680 12230
rect 41600 12160 41680 12190
rect 41720 12230 41800 12260
rect 41720 12190 41740 12230
rect 41780 12190 41800 12230
rect 41720 12160 41800 12190
rect 41840 12230 41920 12260
rect 41840 12190 41860 12230
rect 41900 12190 41920 12230
rect 41840 12160 41920 12190
rect 41960 12230 42040 12260
rect 41960 12190 41980 12230
rect 42020 12190 42040 12230
rect 41960 12160 42040 12190
rect 42080 12230 42160 12260
rect 42080 12190 42100 12230
rect 42140 12190 42160 12230
rect 42080 12160 42160 12190
rect 42200 12230 42280 12260
rect 42200 12190 42220 12230
rect 42260 12190 42280 12230
rect 42200 12160 42280 12190
rect 42320 12230 42400 12260
rect 42320 12190 42340 12230
rect 42380 12190 42400 12230
rect 42320 12160 42400 12190
rect 42440 12230 42520 12260
rect 42440 12190 42460 12230
rect 42500 12190 42520 12230
rect 42440 12160 42520 12190
rect 42560 12230 42640 12260
rect 42560 12190 42580 12230
rect 42620 12190 42640 12230
rect 42560 12160 42640 12190
rect 43920 12230 44000 12260
rect 43920 12190 43940 12230
rect 43980 12190 44000 12230
rect 43920 12160 44000 12190
rect 44040 12230 44120 12260
rect 44040 12190 44060 12230
rect 44100 12190 44120 12230
rect 44040 12160 44120 12190
rect 44160 12230 44240 12260
rect 44160 12190 44180 12230
rect 44220 12190 44240 12230
rect 44160 12160 44240 12190
rect 44280 12230 44360 12260
rect 44280 12190 44300 12230
rect 44340 12190 44360 12230
rect 44280 12160 44360 12190
rect 44400 12230 44480 12260
rect 44400 12190 44420 12230
rect 44460 12190 44480 12230
rect 44400 12160 44480 12190
rect 44520 12230 44600 12260
rect 44520 12190 44540 12230
rect 44580 12190 44600 12230
rect 44520 12160 44600 12190
rect 44640 12230 44720 12260
rect 44640 12190 44660 12230
rect 44700 12190 44720 12230
rect 44640 12160 44720 12190
rect 44760 12230 44840 12260
rect 44760 12190 44780 12230
rect 44820 12190 44840 12230
rect 44760 12160 44840 12190
rect 44880 12230 44960 12260
rect 44880 12190 44900 12230
rect 44940 12190 44960 12230
rect 44880 12160 44960 12190
rect 45000 12230 45080 12260
rect 45000 12190 45020 12230
rect 45060 12190 45080 12230
rect 45000 12160 45080 12190
rect 45120 12230 45200 12260
rect 45120 12190 45140 12230
rect 45180 12190 45200 12230
rect 45120 12160 45200 12190
<< pdiff >>
rect 41580 18426 42260 18480
rect 41580 18392 41632 18426
rect 41666 18392 41722 18426
rect 41756 18392 41812 18426
rect 41846 18392 41902 18426
rect 41936 18392 41992 18426
rect 42026 18392 42082 18426
rect 42116 18392 42172 18426
rect 42206 18392 42260 18426
rect 41580 18336 42260 18392
rect 41580 18302 41632 18336
rect 41666 18302 41722 18336
rect 41756 18302 41812 18336
rect 41846 18302 41902 18336
rect 41936 18302 41992 18336
rect 42026 18302 42082 18336
rect 42116 18302 42172 18336
rect 42206 18302 42260 18336
rect 41580 18246 42260 18302
rect 41580 18212 41632 18246
rect 41666 18212 41722 18246
rect 41756 18212 41812 18246
rect 41846 18212 41902 18246
rect 41936 18212 41992 18246
rect 42026 18212 42082 18246
rect 42116 18212 42172 18246
rect 42206 18212 42260 18246
rect 41580 18156 42260 18212
rect 41580 18122 41632 18156
rect 41666 18122 41722 18156
rect 41756 18122 41812 18156
rect 41846 18122 41902 18156
rect 41936 18122 41992 18156
rect 42026 18122 42082 18156
rect 42116 18122 42172 18156
rect 42206 18122 42260 18156
rect 41580 18066 42260 18122
rect 41580 18032 41632 18066
rect 41666 18032 41722 18066
rect 41756 18032 41812 18066
rect 41846 18032 41902 18066
rect 41936 18032 41992 18066
rect 42026 18032 42082 18066
rect 42116 18032 42172 18066
rect 42206 18032 42260 18066
rect 41580 17976 42260 18032
rect 41580 17942 41632 17976
rect 41666 17942 41722 17976
rect 41756 17942 41812 17976
rect 41846 17942 41902 17976
rect 41936 17942 41992 17976
rect 42026 17942 42082 17976
rect 42116 17942 42172 17976
rect 42206 17942 42260 17976
rect 41580 17886 42260 17942
rect 41580 17852 41632 17886
rect 41666 17852 41722 17886
rect 41756 17852 41812 17886
rect 41846 17852 41902 17886
rect 41936 17852 41992 17886
rect 42026 17852 42082 17886
rect 42116 17852 42172 17886
rect 42206 17852 42260 17886
rect 41580 17800 42260 17852
rect 42940 18426 43620 18480
rect 42940 18392 42992 18426
rect 43026 18392 43082 18426
rect 43116 18392 43172 18426
rect 43206 18392 43262 18426
rect 43296 18392 43352 18426
rect 43386 18392 43442 18426
rect 43476 18392 43532 18426
rect 43566 18392 43620 18426
rect 42940 18336 43620 18392
rect 42940 18302 42992 18336
rect 43026 18302 43082 18336
rect 43116 18302 43172 18336
rect 43206 18302 43262 18336
rect 43296 18302 43352 18336
rect 43386 18302 43442 18336
rect 43476 18302 43532 18336
rect 43566 18302 43620 18336
rect 42940 18246 43620 18302
rect 42940 18212 42992 18246
rect 43026 18212 43082 18246
rect 43116 18212 43172 18246
rect 43206 18212 43262 18246
rect 43296 18212 43352 18246
rect 43386 18212 43442 18246
rect 43476 18212 43532 18246
rect 43566 18212 43620 18246
rect 42940 18156 43620 18212
rect 42940 18122 42992 18156
rect 43026 18122 43082 18156
rect 43116 18122 43172 18156
rect 43206 18122 43262 18156
rect 43296 18122 43352 18156
rect 43386 18122 43442 18156
rect 43476 18122 43532 18156
rect 43566 18122 43620 18156
rect 42940 18066 43620 18122
rect 42940 18032 42992 18066
rect 43026 18032 43082 18066
rect 43116 18032 43172 18066
rect 43206 18032 43262 18066
rect 43296 18032 43352 18066
rect 43386 18032 43442 18066
rect 43476 18032 43532 18066
rect 43566 18032 43620 18066
rect 42940 17976 43620 18032
rect 42940 17942 42992 17976
rect 43026 17942 43082 17976
rect 43116 17942 43172 17976
rect 43206 17942 43262 17976
rect 43296 17942 43352 17976
rect 43386 17942 43442 17976
rect 43476 17942 43532 17976
rect 43566 17942 43620 17976
rect 42940 17886 43620 17942
rect 42940 17852 42992 17886
rect 43026 17852 43082 17886
rect 43116 17852 43172 17886
rect 43206 17852 43262 17886
rect 43296 17852 43352 17886
rect 43386 17852 43442 17886
rect 43476 17852 43532 17886
rect 43566 17852 43620 17886
rect 42940 17800 43620 17852
rect 44300 18426 44980 18480
rect 44300 18392 44352 18426
rect 44386 18392 44442 18426
rect 44476 18392 44532 18426
rect 44566 18392 44622 18426
rect 44656 18392 44712 18426
rect 44746 18392 44802 18426
rect 44836 18392 44892 18426
rect 44926 18392 44980 18426
rect 44300 18336 44980 18392
rect 44300 18302 44352 18336
rect 44386 18302 44442 18336
rect 44476 18302 44532 18336
rect 44566 18302 44622 18336
rect 44656 18302 44712 18336
rect 44746 18302 44802 18336
rect 44836 18302 44892 18336
rect 44926 18302 44980 18336
rect 44300 18246 44980 18302
rect 44300 18212 44352 18246
rect 44386 18212 44442 18246
rect 44476 18212 44532 18246
rect 44566 18212 44622 18246
rect 44656 18212 44712 18246
rect 44746 18212 44802 18246
rect 44836 18212 44892 18246
rect 44926 18212 44980 18246
rect 44300 18156 44980 18212
rect 44300 18122 44352 18156
rect 44386 18122 44442 18156
rect 44476 18122 44532 18156
rect 44566 18122 44622 18156
rect 44656 18122 44712 18156
rect 44746 18122 44802 18156
rect 44836 18122 44892 18156
rect 44926 18122 44980 18156
rect 44300 18066 44980 18122
rect 44300 18032 44352 18066
rect 44386 18032 44442 18066
rect 44476 18032 44532 18066
rect 44566 18032 44622 18066
rect 44656 18032 44712 18066
rect 44746 18032 44802 18066
rect 44836 18032 44892 18066
rect 44926 18032 44980 18066
rect 44300 17976 44980 18032
rect 44300 17942 44352 17976
rect 44386 17942 44442 17976
rect 44476 17942 44532 17976
rect 44566 17942 44622 17976
rect 44656 17942 44712 17976
rect 44746 17942 44802 17976
rect 44836 17942 44892 17976
rect 44926 17942 44980 17976
rect 44300 17886 44980 17942
rect 44300 17852 44352 17886
rect 44386 17852 44442 17886
rect 44476 17852 44532 17886
rect 44566 17852 44622 17886
rect 44656 17852 44712 17886
rect 44746 17852 44802 17886
rect 44836 17852 44892 17886
rect 44926 17852 44980 17886
rect 44300 17800 44980 17852
rect 41580 17066 42260 17120
rect 41580 17032 41632 17066
rect 41666 17032 41722 17066
rect 41756 17032 41812 17066
rect 41846 17032 41902 17066
rect 41936 17032 41992 17066
rect 42026 17032 42082 17066
rect 42116 17032 42172 17066
rect 42206 17032 42260 17066
rect 41580 16976 42260 17032
rect 41580 16942 41632 16976
rect 41666 16942 41722 16976
rect 41756 16942 41812 16976
rect 41846 16942 41902 16976
rect 41936 16942 41992 16976
rect 42026 16942 42082 16976
rect 42116 16942 42172 16976
rect 42206 16942 42260 16976
rect 41580 16886 42260 16942
rect 41580 16852 41632 16886
rect 41666 16852 41722 16886
rect 41756 16852 41812 16886
rect 41846 16852 41902 16886
rect 41936 16852 41992 16886
rect 42026 16852 42082 16886
rect 42116 16852 42172 16886
rect 42206 16852 42260 16886
rect 41580 16796 42260 16852
rect 41580 16762 41632 16796
rect 41666 16762 41722 16796
rect 41756 16762 41812 16796
rect 41846 16762 41902 16796
rect 41936 16762 41992 16796
rect 42026 16762 42082 16796
rect 42116 16762 42172 16796
rect 42206 16762 42260 16796
rect 41580 16706 42260 16762
rect 41580 16672 41632 16706
rect 41666 16672 41722 16706
rect 41756 16672 41812 16706
rect 41846 16672 41902 16706
rect 41936 16672 41992 16706
rect 42026 16672 42082 16706
rect 42116 16672 42172 16706
rect 42206 16672 42260 16706
rect 41580 16616 42260 16672
rect 41580 16582 41632 16616
rect 41666 16582 41722 16616
rect 41756 16582 41812 16616
rect 41846 16582 41902 16616
rect 41936 16582 41992 16616
rect 42026 16582 42082 16616
rect 42116 16582 42172 16616
rect 42206 16582 42260 16616
rect 41580 16526 42260 16582
rect 41580 16492 41632 16526
rect 41666 16492 41722 16526
rect 41756 16492 41812 16526
rect 41846 16492 41902 16526
rect 41936 16492 41992 16526
rect 42026 16492 42082 16526
rect 42116 16492 42172 16526
rect 42206 16492 42260 16526
rect 41580 16440 42260 16492
rect 42940 17066 43620 17120
rect 42940 17032 42992 17066
rect 43026 17032 43082 17066
rect 43116 17032 43172 17066
rect 43206 17032 43262 17066
rect 43296 17032 43352 17066
rect 43386 17032 43442 17066
rect 43476 17032 43532 17066
rect 43566 17032 43620 17066
rect 42940 16976 43620 17032
rect 42940 16942 42992 16976
rect 43026 16942 43082 16976
rect 43116 16942 43172 16976
rect 43206 16942 43262 16976
rect 43296 16942 43352 16976
rect 43386 16942 43442 16976
rect 43476 16942 43532 16976
rect 43566 16942 43620 16976
rect 42940 16886 43620 16942
rect 42940 16852 42992 16886
rect 43026 16852 43082 16886
rect 43116 16852 43172 16886
rect 43206 16852 43262 16886
rect 43296 16852 43352 16886
rect 43386 16852 43442 16886
rect 43476 16852 43532 16886
rect 43566 16852 43620 16886
rect 42940 16796 43620 16852
rect 42940 16762 42992 16796
rect 43026 16762 43082 16796
rect 43116 16762 43172 16796
rect 43206 16762 43262 16796
rect 43296 16762 43352 16796
rect 43386 16762 43442 16796
rect 43476 16762 43532 16796
rect 43566 16762 43620 16796
rect 42940 16706 43620 16762
rect 42940 16672 42992 16706
rect 43026 16672 43082 16706
rect 43116 16672 43172 16706
rect 43206 16672 43262 16706
rect 43296 16672 43352 16706
rect 43386 16672 43442 16706
rect 43476 16672 43532 16706
rect 43566 16672 43620 16706
rect 42940 16616 43620 16672
rect 42940 16582 42992 16616
rect 43026 16582 43082 16616
rect 43116 16582 43172 16616
rect 43206 16582 43262 16616
rect 43296 16582 43352 16616
rect 43386 16582 43442 16616
rect 43476 16582 43532 16616
rect 43566 16582 43620 16616
rect 42940 16526 43620 16582
rect 42940 16492 42992 16526
rect 43026 16492 43082 16526
rect 43116 16492 43172 16526
rect 43206 16492 43262 16526
rect 43296 16492 43352 16526
rect 43386 16492 43442 16526
rect 43476 16492 43532 16526
rect 43566 16492 43620 16526
rect 42940 16440 43620 16492
rect 44300 17066 44980 17120
rect 44300 17032 44352 17066
rect 44386 17032 44442 17066
rect 44476 17032 44532 17066
rect 44566 17032 44622 17066
rect 44656 17032 44712 17066
rect 44746 17032 44802 17066
rect 44836 17032 44892 17066
rect 44926 17032 44980 17066
rect 44300 16976 44980 17032
rect 44300 16942 44352 16976
rect 44386 16942 44442 16976
rect 44476 16942 44532 16976
rect 44566 16942 44622 16976
rect 44656 16942 44712 16976
rect 44746 16942 44802 16976
rect 44836 16942 44892 16976
rect 44926 16942 44980 16976
rect 44300 16886 44980 16942
rect 44300 16852 44352 16886
rect 44386 16852 44442 16886
rect 44476 16852 44532 16886
rect 44566 16852 44622 16886
rect 44656 16852 44712 16886
rect 44746 16852 44802 16886
rect 44836 16852 44892 16886
rect 44926 16852 44980 16886
rect 44300 16796 44980 16852
rect 44300 16762 44352 16796
rect 44386 16762 44442 16796
rect 44476 16762 44532 16796
rect 44566 16762 44622 16796
rect 44656 16762 44712 16796
rect 44746 16762 44802 16796
rect 44836 16762 44892 16796
rect 44926 16762 44980 16796
rect 44300 16706 44980 16762
rect 44300 16672 44352 16706
rect 44386 16672 44442 16706
rect 44476 16672 44532 16706
rect 44566 16672 44622 16706
rect 44656 16672 44712 16706
rect 44746 16672 44802 16706
rect 44836 16672 44892 16706
rect 44926 16672 44980 16706
rect 44300 16616 44980 16672
rect 44300 16582 44352 16616
rect 44386 16582 44442 16616
rect 44476 16582 44532 16616
rect 44566 16582 44622 16616
rect 44656 16582 44712 16616
rect 44746 16582 44802 16616
rect 44836 16582 44892 16616
rect 44926 16582 44980 16616
rect 44300 16526 44980 16582
rect 44300 16492 44352 16526
rect 44386 16492 44442 16526
rect 44476 16492 44532 16526
rect 44566 16492 44622 16526
rect 44656 16492 44712 16526
rect 44746 16492 44802 16526
rect 44836 16492 44892 16526
rect 44926 16492 44980 16526
rect 44300 16440 44980 16492
rect 41580 15706 42260 15760
rect 41580 15672 41632 15706
rect 41666 15672 41722 15706
rect 41756 15672 41812 15706
rect 41846 15672 41902 15706
rect 41936 15672 41992 15706
rect 42026 15672 42082 15706
rect 42116 15672 42172 15706
rect 42206 15672 42260 15706
rect 41580 15616 42260 15672
rect 41580 15582 41632 15616
rect 41666 15582 41722 15616
rect 41756 15582 41812 15616
rect 41846 15582 41902 15616
rect 41936 15582 41992 15616
rect 42026 15582 42082 15616
rect 42116 15582 42172 15616
rect 42206 15582 42260 15616
rect 41580 15526 42260 15582
rect 41580 15492 41632 15526
rect 41666 15492 41722 15526
rect 41756 15492 41812 15526
rect 41846 15492 41902 15526
rect 41936 15492 41992 15526
rect 42026 15492 42082 15526
rect 42116 15492 42172 15526
rect 42206 15492 42260 15526
rect 41580 15436 42260 15492
rect 41580 15402 41632 15436
rect 41666 15402 41722 15436
rect 41756 15402 41812 15436
rect 41846 15402 41902 15436
rect 41936 15402 41992 15436
rect 42026 15402 42082 15436
rect 42116 15402 42172 15436
rect 42206 15402 42260 15436
rect 41580 15346 42260 15402
rect 41580 15312 41632 15346
rect 41666 15312 41722 15346
rect 41756 15312 41812 15346
rect 41846 15312 41902 15346
rect 41936 15312 41992 15346
rect 42026 15312 42082 15346
rect 42116 15312 42172 15346
rect 42206 15312 42260 15346
rect 41580 15256 42260 15312
rect 41580 15222 41632 15256
rect 41666 15222 41722 15256
rect 41756 15222 41812 15256
rect 41846 15222 41902 15256
rect 41936 15222 41992 15256
rect 42026 15222 42082 15256
rect 42116 15222 42172 15256
rect 42206 15222 42260 15256
rect 41580 15166 42260 15222
rect 41580 15132 41632 15166
rect 41666 15132 41722 15166
rect 41756 15132 41812 15166
rect 41846 15132 41902 15166
rect 41936 15132 41992 15166
rect 42026 15132 42082 15166
rect 42116 15132 42172 15166
rect 42206 15132 42260 15166
rect 41580 15080 42260 15132
rect 42940 15706 43620 15760
rect 42940 15672 42992 15706
rect 43026 15672 43082 15706
rect 43116 15672 43172 15706
rect 43206 15672 43262 15706
rect 43296 15672 43352 15706
rect 43386 15672 43442 15706
rect 43476 15672 43532 15706
rect 43566 15672 43620 15706
rect 42940 15616 43620 15672
rect 42940 15582 42992 15616
rect 43026 15582 43082 15616
rect 43116 15582 43172 15616
rect 43206 15582 43262 15616
rect 43296 15582 43352 15616
rect 43386 15582 43442 15616
rect 43476 15582 43532 15616
rect 43566 15582 43620 15616
rect 42940 15526 43620 15582
rect 42940 15492 42992 15526
rect 43026 15492 43082 15526
rect 43116 15492 43172 15526
rect 43206 15492 43262 15526
rect 43296 15492 43352 15526
rect 43386 15492 43442 15526
rect 43476 15492 43532 15526
rect 43566 15492 43620 15526
rect 42940 15436 43620 15492
rect 42940 15402 42992 15436
rect 43026 15402 43082 15436
rect 43116 15402 43172 15436
rect 43206 15402 43262 15436
rect 43296 15402 43352 15436
rect 43386 15402 43442 15436
rect 43476 15402 43532 15436
rect 43566 15402 43620 15436
rect 42940 15346 43620 15402
rect 42940 15312 42992 15346
rect 43026 15312 43082 15346
rect 43116 15312 43172 15346
rect 43206 15312 43262 15346
rect 43296 15312 43352 15346
rect 43386 15312 43442 15346
rect 43476 15312 43532 15346
rect 43566 15312 43620 15346
rect 42940 15256 43620 15312
rect 42940 15222 42992 15256
rect 43026 15222 43082 15256
rect 43116 15222 43172 15256
rect 43206 15222 43262 15256
rect 43296 15222 43352 15256
rect 43386 15222 43442 15256
rect 43476 15222 43532 15256
rect 43566 15222 43620 15256
rect 42940 15166 43620 15222
rect 42940 15132 42992 15166
rect 43026 15132 43082 15166
rect 43116 15132 43172 15166
rect 43206 15132 43262 15166
rect 43296 15132 43352 15166
rect 43386 15132 43442 15166
rect 43476 15132 43532 15166
rect 43566 15132 43620 15166
rect 42940 15080 43620 15132
rect 44300 15706 44980 15760
rect 44300 15672 44352 15706
rect 44386 15672 44442 15706
rect 44476 15672 44532 15706
rect 44566 15672 44622 15706
rect 44656 15672 44712 15706
rect 44746 15672 44802 15706
rect 44836 15672 44892 15706
rect 44926 15672 44980 15706
rect 44300 15616 44980 15672
rect 44300 15582 44352 15616
rect 44386 15582 44442 15616
rect 44476 15582 44532 15616
rect 44566 15582 44622 15616
rect 44656 15582 44712 15616
rect 44746 15582 44802 15616
rect 44836 15582 44892 15616
rect 44926 15582 44980 15616
rect 44300 15526 44980 15582
rect 44300 15492 44352 15526
rect 44386 15492 44442 15526
rect 44476 15492 44532 15526
rect 44566 15492 44622 15526
rect 44656 15492 44712 15526
rect 44746 15492 44802 15526
rect 44836 15492 44892 15526
rect 44926 15492 44980 15526
rect 44300 15436 44980 15492
rect 44300 15402 44352 15436
rect 44386 15402 44442 15436
rect 44476 15402 44532 15436
rect 44566 15402 44622 15436
rect 44656 15402 44712 15436
rect 44746 15402 44802 15436
rect 44836 15402 44892 15436
rect 44926 15402 44980 15436
rect 44300 15346 44980 15402
rect 44300 15312 44352 15346
rect 44386 15312 44442 15346
rect 44476 15312 44532 15346
rect 44566 15312 44622 15346
rect 44656 15312 44712 15346
rect 44746 15312 44802 15346
rect 44836 15312 44892 15346
rect 44926 15312 44980 15346
rect 44300 15256 44980 15312
rect 44300 15222 44352 15256
rect 44386 15222 44442 15256
rect 44476 15222 44532 15256
rect 44566 15222 44622 15256
rect 44656 15222 44712 15256
rect 44746 15222 44802 15256
rect 44836 15222 44892 15256
rect 44926 15222 44980 15256
rect 44300 15166 44980 15222
rect 44300 15132 44352 15166
rect 44386 15132 44442 15166
rect 44476 15132 44532 15166
rect 44566 15132 44622 15166
rect 44656 15132 44712 15166
rect 44746 15132 44802 15166
rect 44836 15132 44892 15166
rect 44926 15132 44980 15166
rect 44300 15080 44980 15132
rect 40520 11390 40600 11420
rect 40520 11350 40540 11390
rect 40580 11350 40600 11390
rect 40520 11290 40600 11350
rect 40520 11250 40540 11290
rect 40580 11250 40600 11290
rect 40520 11220 40600 11250
rect 40640 11390 40720 11420
rect 40640 11350 40660 11390
rect 40700 11350 40720 11390
rect 40640 11290 40720 11350
rect 40640 11250 40660 11290
rect 40700 11250 40720 11290
rect 40640 11220 40720 11250
rect 40760 11390 40840 11420
rect 40760 11350 40780 11390
rect 40820 11350 40840 11390
rect 40760 11290 40840 11350
rect 40760 11250 40780 11290
rect 40820 11250 40840 11290
rect 40760 11220 40840 11250
rect 40880 11390 40960 11420
rect 40880 11350 40900 11390
rect 40940 11350 40960 11390
rect 40880 11290 40960 11350
rect 40880 11250 40900 11290
rect 40940 11250 40960 11290
rect 40880 11220 40960 11250
rect 41000 11390 41080 11420
rect 41000 11350 41020 11390
rect 41060 11350 41080 11390
rect 41000 11290 41080 11350
rect 41000 11250 41020 11290
rect 41060 11250 41080 11290
rect 41000 11220 41080 11250
rect 41120 11390 41200 11420
rect 41120 11350 41140 11390
rect 41180 11350 41200 11390
rect 41120 11290 41200 11350
rect 41120 11250 41140 11290
rect 41180 11250 41200 11290
rect 41120 11220 41200 11250
rect 41240 11390 41320 11420
rect 41240 11350 41260 11390
rect 41300 11350 41320 11390
rect 41240 11290 41320 11350
rect 41240 11250 41260 11290
rect 41300 11250 41320 11290
rect 41240 11220 41320 11250
rect 41360 11390 41440 11420
rect 41360 11350 41380 11390
rect 41420 11350 41440 11390
rect 41360 11290 41440 11350
rect 41360 11250 41380 11290
rect 41420 11250 41440 11290
rect 41360 11220 41440 11250
rect 41480 11390 41560 11420
rect 41480 11350 41500 11390
rect 41540 11350 41560 11390
rect 41480 11290 41560 11350
rect 41480 11250 41500 11290
rect 41540 11250 41560 11290
rect 41480 11220 41560 11250
rect 41600 11390 41680 11420
rect 41600 11350 41620 11390
rect 41660 11350 41680 11390
rect 41600 11290 41680 11350
rect 41600 11250 41620 11290
rect 41660 11250 41680 11290
rect 41600 11220 41680 11250
rect 41720 11390 41800 11420
rect 41720 11350 41740 11390
rect 41780 11350 41800 11390
rect 41720 11290 41800 11350
rect 41720 11250 41740 11290
rect 41780 11250 41800 11290
rect 41720 11220 41800 11250
rect 41840 11390 41920 11420
rect 41840 11350 41860 11390
rect 41900 11350 41920 11390
rect 41840 11290 41920 11350
rect 41840 11250 41860 11290
rect 41900 11250 41920 11290
rect 41840 11220 41920 11250
rect 41960 11390 42040 11420
rect 41960 11350 41980 11390
rect 42020 11350 42040 11390
rect 41960 11290 42040 11350
rect 41960 11250 41980 11290
rect 42020 11250 42040 11290
rect 41960 11220 42040 11250
rect 42080 11390 42160 11420
rect 42080 11350 42100 11390
rect 42140 11350 42160 11390
rect 42080 11290 42160 11350
rect 42080 11250 42100 11290
rect 42140 11250 42160 11290
rect 42080 11220 42160 11250
rect 42200 11390 42280 11420
rect 42200 11350 42220 11390
rect 42260 11350 42280 11390
rect 42200 11290 42280 11350
rect 42200 11250 42220 11290
rect 42260 11250 42280 11290
rect 42200 11220 42280 11250
rect 42320 11390 42400 11420
rect 42320 11350 42340 11390
rect 42380 11350 42400 11390
rect 42320 11290 42400 11350
rect 42320 11250 42340 11290
rect 42380 11250 42400 11290
rect 42320 11220 42400 11250
rect 42440 11390 42520 11420
rect 42440 11350 42460 11390
rect 42500 11350 42520 11390
rect 42440 11290 42520 11350
rect 42440 11250 42460 11290
rect 42500 11250 42520 11290
rect 42440 11220 42520 11250
rect 42560 11390 42640 11420
rect 42560 11350 42580 11390
rect 42620 11350 42640 11390
rect 42560 11290 42640 11350
rect 42560 11250 42580 11290
rect 42620 11250 42640 11290
rect 42560 11220 42640 11250
rect 42680 11390 42760 11420
rect 42680 11350 42700 11390
rect 42740 11350 42760 11390
rect 42680 11290 42760 11350
rect 42680 11250 42700 11290
rect 42740 11250 42760 11290
rect 42680 11220 42760 11250
rect 42800 11390 42880 11420
rect 42800 11350 42820 11390
rect 42860 11350 42880 11390
rect 42800 11290 42880 11350
rect 42800 11250 42820 11290
rect 42860 11250 42880 11290
rect 42800 11220 42880 11250
rect 42920 11390 43000 11420
rect 42920 11350 42940 11390
rect 42980 11350 43000 11390
rect 42920 11290 43000 11350
rect 42920 11250 42940 11290
rect 42980 11250 43000 11290
rect 42920 11220 43000 11250
rect 43560 11390 43640 11420
rect 43560 11350 43580 11390
rect 43620 11350 43640 11390
rect 43560 11290 43640 11350
rect 43560 11250 43580 11290
rect 43620 11250 43640 11290
rect 43560 11220 43640 11250
rect 43680 11390 43760 11420
rect 43680 11350 43700 11390
rect 43740 11350 43760 11390
rect 43680 11290 43760 11350
rect 43680 11250 43700 11290
rect 43740 11250 43760 11290
rect 43680 11220 43760 11250
rect 43800 11390 43880 11420
rect 43800 11350 43820 11390
rect 43860 11350 43880 11390
rect 43800 11290 43880 11350
rect 43800 11250 43820 11290
rect 43860 11250 43880 11290
rect 43800 11220 43880 11250
rect 43920 11390 44000 11420
rect 43920 11350 43940 11390
rect 43980 11350 44000 11390
rect 43920 11290 44000 11350
rect 43920 11250 43940 11290
rect 43980 11250 44000 11290
rect 43920 11220 44000 11250
rect 44040 11390 44120 11420
rect 44040 11350 44060 11390
rect 44100 11350 44120 11390
rect 44040 11290 44120 11350
rect 44040 11250 44060 11290
rect 44100 11250 44120 11290
rect 44040 11220 44120 11250
rect 44160 11390 44240 11420
rect 44160 11350 44180 11390
rect 44220 11350 44240 11390
rect 44160 11290 44240 11350
rect 44160 11250 44180 11290
rect 44220 11250 44240 11290
rect 44160 11220 44240 11250
rect 44280 11390 44360 11420
rect 44280 11350 44300 11390
rect 44340 11350 44360 11390
rect 44280 11290 44360 11350
rect 44280 11250 44300 11290
rect 44340 11250 44360 11290
rect 44280 11220 44360 11250
rect 44400 11390 44480 11420
rect 44400 11350 44420 11390
rect 44460 11350 44480 11390
rect 44400 11290 44480 11350
rect 44400 11250 44420 11290
rect 44460 11250 44480 11290
rect 44400 11220 44480 11250
rect 44520 11390 44600 11420
rect 44520 11350 44540 11390
rect 44580 11350 44600 11390
rect 44520 11290 44600 11350
rect 44520 11250 44540 11290
rect 44580 11250 44600 11290
rect 44520 11220 44600 11250
rect 44640 11390 44720 11420
rect 44640 11350 44660 11390
rect 44700 11350 44720 11390
rect 44640 11290 44720 11350
rect 44640 11250 44660 11290
rect 44700 11250 44720 11290
rect 44640 11220 44720 11250
rect 44760 11390 44840 11420
rect 44760 11350 44780 11390
rect 44820 11350 44840 11390
rect 44760 11290 44840 11350
rect 44760 11250 44780 11290
rect 44820 11250 44840 11290
rect 44760 11220 44840 11250
rect 44880 11390 44960 11420
rect 44880 11350 44900 11390
rect 44940 11350 44960 11390
rect 44880 11290 44960 11350
rect 44880 11250 44900 11290
rect 44940 11250 44960 11290
rect 44880 11220 44960 11250
rect 45000 11390 45080 11420
rect 45000 11350 45020 11390
rect 45060 11350 45080 11390
rect 45000 11290 45080 11350
rect 45000 11250 45020 11290
rect 45060 11250 45080 11290
rect 45000 11220 45080 11250
rect 45120 11390 45200 11420
rect 45120 11350 45140 11390
rect 45180 11350 45200 11390
rect 45120 11290 45200 11350
rect 45120 11250 45140 11290
rect 45180 11250 45200 11290
rect 45120 11220 45200 11250
rect 45240 11390 45320 11420
rect 45240 11350 45260 11390
rect 45300 11350 45320 11390
rect 45240 11290 45320 11350
rect 45240 11250 45260 11290
rect 45300 11250 45320 11290
rect 45240 11220 45320 11250
rect 45360 11390 45440 11420
rect 45360 11350 45380 11390
rect 45420 11350 45440 11390
rect 45360 11290 45440 11350
rect 45360 11250 45380 11290
rect 45420 11250 45440 11290
rect 45360 11220 45440 11250
rect 45480 11390 45560 11420
rect 45480 11350 45500 11390
rect 45540 11350 45560 11390
rect 45480 11290 45560 11350
rect 45480 11250 45500 11290
rect 45540 11250 45560 11290
rect 45480 11220 45560 11250
rect 45600 11390 45680 11420
rect 45600 11350 45620 11390
rect 45660 11350 45680 11390
rect 45600 11290 45680 11350
rect 45600 11250 45620 11290
rect 45660 11250 45680 11290
rect 45600 11220 45680 11250
rect 45720 11390 45800 11420
rect 45720 11350 45740 11390
rect 45780 11350 45800 11390
rect 45720 11290 45800 11350
rect 45720 11250 45740 11290
rect 45780 11250 45800 11290
rect 45720 11220 45800 11250
rect 45840 11390 45920 11420
rect 45840 11350 45860 11390
rect 45900 11350 45920 11390
rect 45840 11290 45920 11350
rect 45840 11250 45860 11290
rect 45900 11250 45920 11290
rect 45840 11220 45920 11250
rect 45960 11390 46040 11420
rect 45960 11350 45980 11390
rect 46020 11350 46040 11390
rect 45960 11290 46040 11350
rect 45960 11250 45980 11290
rect 46020 11250 46040 11290
rect 45960 11220 46040 11250
rect 41620 10230 41700 10260
rect 41620 10190 41640 10230
rect 41680 10190 41700 10230
rect 41620 10130 41700 10190
rect 41620 10090 41640 10130
rect 41680 10090 41700 10130
rect 41620 10030 41700 10090
rect 41620 9990 41640 10030
rect 41680 9990 41700 10030
rect 41620 9930 41700 9990
rect 41620 9890 41640 9930
rect 41680 9890 41700 9930
rect 41620 9830 41700 9890
rect 41620 9790 41640 9830
rect 41680 9790 41700 9830
rect 41620 9730 41700 9790
rect 41620 9690 41640 9730
rect 41680 9690 41700 9730
rect 41620 9660 41700 9690
rect 41800 10230 41880 10260
rect 41800 10190 41820 10230
rect 41860 10190 41880 10230
rect 41800 10130 41880 10190
rect 41800 10090 41820 10130
rect 41860 10090 41880 10130
rect 41800 10030 41880 10090
rect 41800 9990 41820 10030
rect 41860 9990 41880 10030
rect 41800 9930 41880 9990
rect 41800 9890 41820 9930
rect 41860 9890 41880 9930
rect 41800 9830 41880 9890
rect 41800 9790 41820 9830
rect 41860 9790 41880 9830
rect 41800 9730 41880 9790
rect 41800 9690 41820 9730
rect 41860 9690 41880 9730
rect 41800 9660 41880 9690
rect 41980 10230 42060 10260
rect 41980 10190 42000 10230
rect 42040 10190 42060 10230
rect 41980 10130 42060 10190
rect 41980 10090 42000 10130
rect 42040 10090 42060 10130
rect 41980 10030 42060 10090
rect 41980 9990 42000 10030
rect 42040 9990 42060 10030
rect 41980 9930 42060 9990
rect 41980 9890 42000 9930
rect 42040 9890 42060 9930
rect 41980 9830 42060 9890
rect 41980 9790 42000 9830
rect 42040 9790 42060 9830
rect 41980 9730 42060 9790
rect 41980 9690 42000 9730
rect 42040 9690 42060 9730
rect 41980 9660 42060 9690
rect 42160 10230 42240 10260
rect 42160 10190 42180 10230
rect 42220 10190 42240 10230
rect 42160 10130 42240 10190
rect 42160 10090 42180 10130
rect 42220 10090 42240 10130
rect 42160 10030 42240 10090
rect 42160 9990 42180 10030
rect 42220 9990 42240 10030
rect 42160 9930 42240 9990
rect 42160 9890 42180 9930
rect 42220 9890 42240 9930
rect 42160 9830 42240 9890
rect 42160 9790 42180 9830
rect 42220 9790 42240 9830
rect 42160 9730 42240 9790
rect 42160 9690 42180 9730
rect 42220 9690 42240 9730
rect 42160 9660 42240 9690
rect 42340 10230 42420 10260
rect 42340 10190 42360 10230
rect 42400 10190 42420 10230
rect 42340 10130 42420 10190
rect 42340 10090 42360 10130
rect 42400 10090 42420 10130
rect 42340 10030 42420 10090
rect 42340 9990 42360 10030
rect 42400 9990 42420 10030
rect 42340 9930 42420 9990
rect 42340 9890 42360 9930
rect 42400 9890 42420 9930
rect 42340 9830 42420 9890
rect 42340 9790 42360 9830
rect 42400 9790 42420 9830
rect 42340 9730 42420 9790
rect 42340 9690 42360 9730
rect 42400 9690 42420 9730
rect 42340 9660 42420 9690
rect 42520 10230 42600 10260
rect 42520 10190 42540 10230
rect 42580 10190 42600 10230
rect 42520 10130 42600 10190
rect 42520 10090 42540 10130
rect 42580 10090 42600 10130
rect 42520 10030 42600 10090
rect 42520 9990 42540 10030
rect 42580 9990 42600 10030
rect 42520 9930 42600 9990
rect 42520 9890 42540 9930
rect 42580 9890 42600 9930
rect 42520 9830 42600 9890
rect 42520 9790 42540 9830
rect 42580 9790 42600 9830
rect 42520 9730 42600 9790
rect 42520 9690 42540 9730
rect 42580 9690 42600 9730
rect 42520 9660 42600 9690
rect 42700 10230 42780 10260
rect 42700 10190 42720 10230
rect 42760 10190 42780 10230
rect 42700 10130 42780 10190
rect 42700 10090 42720 10130
rect 42760 10090 42780 10130
rect 42700 10030 42780 10090
rect 42700 9990 42720 10030
rect 42760 9990 42780 10030
rect 42700 9930 42780 9990
rect 42700 9890 42720 9930
rect 42760 9890 42780 9930
rect 42700 9830 42780 9890
rect 42700 9790 42720 9830
rect 42760 9790 42780 9830
rect 42700 9730 42780 9790
rect 42700 9690 42720 9730
rect 42760 9690 42780 9730
rect 42700 9660 42780 9690
rect 42880 10230 42960 10260
rect 42880 10190 42900 10230
rect 42940 10190 42960 10230
rect 42880 10130 42960 10190
rect 42880 10090 42900 10130
rect 42940 10090 42960 10130
rect 42880 10030 42960 10090
rect 42880 9990 42900 10030
rect 42940 9990 42960 10030
rect 42880 9930 42960 9990
rect 42880 9890 42900 9930
rect 42940 9890 42960 9930
rect 42880 9830 42960 9890
rect 42880 9790 42900 9830
rect 42940 9790 42960 9830
rect 42880 9730 42960 9790
rect 42880 9690 42900 9730
rect 42940 9690 42960 9730
rect 42880 9660 42960 9690
rect 43060 10230 43140 10260
rect 43060 10190 43080 10230
rect 43120 10190 43140 10230
rect 43060 10130 43140 10190
rect 43060 10090 43080 10130
rect 43120 10090 43140 10130
rect 43060 10030 43140 10090
rect 43060 9990 43080 10030
rect 43120 9990 43140 10030
rect 43060 9930 43140 9990
rect 43060 9890 43080 9930
rect 43120 9890 43140 9930
rect 43060 9830 43140 9890
rect 43060 9790 43080 9830
rect 43120 9790 43140 9830
rect 43060 9730 43140 9790
rect 43060 9690 43080 9730
rect 43120 9690 43140 9730
rect 43060 9660 43140 9690
rect 43240 10230 43320 10260
rect 43240 10190 43260 10230
rect 43300 10190 43320 10230
rect 43240 10130 43320 10190
rect 43240 10090 43260 10130
rect 43300 10090 43320 10130
rect 43240 10030 43320 10090
rect 43240 9990 43260 10030
rect 43300 9990 43320 10030
rect 43240 9930 43320 9990
rect 43240 9890 43260 9930
rect 43300 9890 43320 9930
rect 43240 9830 43320 9890
rect 43240 9790 43260 9830
rect 43300 9790 43320 9830
rect 43240 9730 43320 9790
rect 43240 9690 43260 9730
rect 43300 9690 43320 9730
rect 43240 9660 43320 9690
rect 43420 10230 43500 10260
rect 43420 10190 43440 10230
rect 43480 10190 43500 10230
rect 43420 10130 43500 10190
rect 43420 10090 43440 10130
rect 43480 10090 43500 10130
rect 43420 10030 43500 10090
rect 43420 9990 43440 10030
rect 43480 9990 43500 10030
rect 43420 9930 43500 9990
rect 43420 9890 43440 9930
rect 43480 9890 43500 9930
rect 43420 9830 43500 9890
rect 43420 9790 43440 9830
rect 43480 9790 43500 9830
rect 43420 9730 43500 9790
rect 43420 9690 43440 9730
rect 43480 9690 43500 9730
rect 43420 9660 43500 9690
rect 43600 10230 43680 10260
rect 43600 10190 43620 10230
rect 43660 10190 43680 10230
rect 43600 10130 43680 10190
rect 43600 10090 43620 10130
rect 43660 10090 43680 10130
rect 43600 10030 43680 10090
rect 43600 9990 43620 10030
rect 43660 9990 43680 10030
rect 43600 9930 43680 9990
rect 43600 9890 43620 9930
rect 43660 9890 43680 9930
rect 43600 9830 43680 9890
rect 43600 9790 43620 9830
rect 43660 9790 43680 9830
rect 43600 9730 43680 9790
rect 43600 9690 43620 9730
rect 43660 9690 43680 9730
rect 43600 9660 43680 9690
rect 43780 10230 43860 10260
rect 43780 10190 43800 10230
rect 43840 10190 43860 10230
rect 43780 10130 43860 10190
rect 43780 10090 43800 10130
rect 43840 10090 43860 10130
rect 43780 10030 43860 10090
rect 43780 9990 43800 10030
rect 43840 9990 43860 10030
rect 43780 9930 43860 9990
rect 43780 9890 43800 9930
rect 43840 9890 43860 9930
rect 43780 9830 43860 9890
rect 43780 9790 43800 9830
rect 43840 9790 43860 9830
rect 43780 9730 43860 9790
rect 43780 9690 43800 9730
rect 43840 9690 43860 9730
rect 43780 9660 43860 9690
rect 43960 10230 44040 10260
rect 43960 10190 43980 10230
rect 44020 10190 44040 10230
rect 43960 10130 44040 10190
rect 43960 10090 43980 10130
rect 44020 10090 44040 10130
rect 43960 10030 44040 10090
rect 43960 9990 43980 10030
rect 44020 9990 44040 10030
rect 43960 9930 44040 9990
rect 43960 9890 43980 9930
rect 44020 9890 44040 9930
rect 43960 9830 44040 9890
rect 43960 9790 43980 9830
rect 44020 9790 44040 9830
rect 43960 9730 44040 9790
rect 43960 9690 43980 9730
rect 44020 9690 44040 9730
rect 43960 9660 44040 9690
rect 44140 10230 44220 10260
rect 44140 10190 44160 10230
rect 44200 10190 44220 10230
rect 44140 10130 44220 10190
rect 44140 10090 44160 10130
rect 44200 10090 44220 10130
rect 44140 10030 44220 10090
rect 44140 9990 44160 10030
rect 44200 9990 44220 10030
rect 44140 9930 44220 9990
rect 44140 9890 44160 9930
rect 44200 9890 44220 9930
rect 44140 9830 44220 9890
rect 44140 9790 44160 9830
rect 44200 9790 44220 9830
rect 44140 9730 44220 9790
rect 44140 9690 44160 9730
rect 44200 9690 44220 9730
rect 44140 9660 44220 9690
rect 44320 10230 44400 10260
rect 44320 10190 44340 10230
rect 44380 10190 44400 10230
rect 44320 10130 44400 10190
rect 44320 10090 44340 10130
rect 44380 10090 44400 10130
rect 44320 10030 44400 10090
rect 44320 9990 44340 10030
rect 44380 9990 44400 10030
rect 44320 9930 44400 9990
rect 44320 9890 44340 9930
rect 44380 9890 44400 9930
rect 44320 9830 44400 9890
rect 44320 9790 44340 9830
rect 44380 9790 44400 9830
rect 44320 9730 44400 9790
rect 44320 9690 44340 9730
rect 44380 9690 44400 9730
rect 44320 9660 44400 9690
rect 44500 10230 44580 10260
rect 44500 10190 44520 10230
rect 44560 10190 44580 10230
rect 44500 10130 44580 10190
rect 44500 10090 44520 10130
rect 44560 10090 44580 10130
rect 44500 10030 44580 10090
rect 44500 9990 44520 10030
rect 44560 9990 44580 10030
rect 44500 9930 44580 9990
rect 44500 9890 44520 9930
rect 44560 9890 44580 9930
rect 44500 9830 44580 9890
rect 44500 9790 44520 9830
rect 44560 9790 44580 9830
rect 44500 9730 44580 9790
rect 44500 9690 44520 9730
rect 44560 9690 44580 9730
rect 44500 9660 44580 9690
rect 44680 10230 44760 10260
rect 44680 10190 44700 10230
rect 44740 10190 44760 10230
rect 44680 10130 44760 10190
rect 44680 10090 44700 10130
rect 44740 10090 44760 10130
rect 44680 10030 44760 10090
rect 44680 9990 44700 10030
rect 44740 9990 44760 10030
rect 44680 9930 44760 9990
rect 44680 9890 44700 9930
rect 44740 9890 44760 9930
rect 44680 9830 44760 9890
rect 44680 9790 44700 9830
rect 44740 9790 44760 9830
rect 44680 9730 44760 9790
rect 44680 9690 44700 9730
rect 44740 9690 44760 9730
rect 44680 9660 44760 9690
rect 44860 10230 44940 10260
rect 44860 10190 44880 10230
rect 44920 10190 44940 10230
rect 44860 10130 44940 10190
rect 44860 10090 44880 10130
rect 44920 10090 44940 10130
rect 44860 10030 44940 10090
rect 44860 9990 44880 10030
rect 44920 9990 44940 10030
rect 44860 9930 44940 9990
rect 44860 9890 44880 9930
rect 44920 9890 44940 9930
rect 44860 9830 44940 9890
rect 45480 10030 45570 10060
rect 45480 9990 45510 10030
rect 45550 9990 45570 10030
rect 45480 9930 45570 9990
rect 45480 9890 45510 9930
rect 45550 9890 45570 9930
rect 45480 9860 45570 9890
rect 45600 10030 45680 10060
rect 45600 9990 45620 10030
rect 45660 9990 45680 10030
rect 45600 9930 45680 9990
rect 45600 9890 45620 9930
rect 45660 9890 45680 9930
rect 45600 9860 45680 9890
rect 45710 10030 45790 10060
rect 45710 9990 45730 10030
rect 45770 9990 45790 10030
rect 45710 9930 45790 9990
rect 45710 9890 45730 9930
rect 45770 9890 45790 9930
rect 45710 9860 45790 9890
rect 45820 10030 45900 10060
rect 45820 9990 45840 10030
rect 45880 9990 45900 10030
rect 45820 9930 45900 9990
rect 45820 9890 45840 9930
rect 45880 9890 45900 9930
rect 45820 9860 45900 9890
rect 45930 10030 46010 10060
rect 45930 9990 45950 10030
rect 45990 9990 46010 10030
rect 45930 9930 46010 9990
rect 45930 9890 45950 9930
rect 45990 9890 46010 9930
rect 45930 9860 46010 9890
rect 44860 9790 44880 9830
rect 44920 9790 44940 9830
rect 44860 9730 44940 9790
rect 44860 9690 44880 9730
rect 44920 9690 44940 9730
rect 44860 9660 44940 9690
rect 41630 9230 41710 9260
rect 41630 9190 41650 9230
rect 41690 9190 41710 9230
rect 41630 9130 41710 9190
rect 41630 9090 41650 9130
rect 41690 9090 41710 9130
rect 41630 9060 41710 9090
rect 41740 9230 41820 9260
rect 41740 9190 41760 9230
rect 41800 9190 41820 9230
rect 41740 9130 41820 9190
rect 41740 9090 41760 9130
rect 41800 9090 41820 9130
rect 41740 9060 41820 9090
rect 41850 9230 41930 9260
rect 41850 9190 41870 9230
rect 41910 9190 41930 9230
rect 41850 9130 41930 9190
rect 41850 9090 41870 9130
rect 41910 9090 41930 9130
rect 41850 9060 41930 9090
rect 41960 9230 42040 9260
rect 41960 9190 41980 9230
rect 42020 9190 42040 9230
rect 41960 9130 42040 9190
rect 41960 9090 41980 9130
rect 42020 9090 42040 9130
rect 41960 9060 42040 9090
rect 42070 9230 42150 9260
rect 42070 9190 42090 9230
rect 42130 9190 42150 9230
rect 42070 9130 42150 9190
rect 42070 9090 42090 9130
rect 42130 9090 42150 9130
rect 42070 9060 42150 9090
rect 42180 9230 42260 9260
rect 42180 9190 42200 9230
rect 42240 9190 42260 9230
rect 42180 9130 42260 9190
rect 42180 9090 42200 9130
rect 42240 9090 42260 9130
rect 42180 9060 42260 9090
rect 42290 9230 42370 9260
rect 42290 9190 42310 9230
rect 42350 9190 42370 9230
rect 42290 9130 42370 9190
rect 42290 9090 42310 9130
rect 42350 9090 42370 9130
rect 42290 9060 42370 9090
rect 42400 9230 42480 9260
rect 42400 9190 42420 9230
rect 42460 9190 42480 9230
rect 42400 9130 42480 9190
rect 42400 9090 42420 9130
rect 42460 9090 42480 9130
rect 42400 9060 42480 9090
rect 42510 9230 42590 9260
rect 42510 9190 42530 9230
rect 42570 9190 42590 9230
rect 42510 9130 42590 9190
rect 42510 9090 42530 9130
rect 42570 9090 42590 9130
rect 42510 9060 42590 9090
rect 42620 9230 42700 9260
rect 42620 9190 42640 9230
rect 42680 9190 42700 9230
rect 42620 9130 42700 9190
rect 42620 9090 42640 9130
rect 42680 9090 42700 9130
rect 42620 9060 42700 9090
rect 42730 9230 42810 9260
rect 42730 9190 42750 9230
rect 42790 9190 42810 9230
rect 42730 9130 42810 9190
rect 42730 9090 42750 9130
rect 42790 9090 42810 9130
rect 42730 9060 42810 9090
rect 42840 9230 42920 9260
rect 42840 9190 42860 9230
rect 42900 9190 42920 9230
rect 42840 9130 42920 9190
rect 42840 9090 42860 9130
rect 42900 9090 42920 9130
rect 42840 9060 42920 9090
rect 42950 9230 43030 9260
rect 42950 9190 42970 9230
rect 43010 9190 43030 9230
rect 42950 9130 43030 9190
rect 42950 9090 42970 9130
rect 43010 9090 43030 9130
rect 42950 9060 43030 9090
rect 43530 9230 43610 9260
rect 43530 9190 43550 9230
rect 43590 9190 43610 9230
rect 43530 9130 43610 9190
rect 43530 9090 43550 9130
rect 43590 9090 43610 9130
rect 43530 9060 43610 9090
rect 43640 9230 43720 9260
rect 43640 9190 43660 9230
rect 43700 9190 43720 9230
rect 43640 9130 43720 9190
rect 43640 9090 43660 9130
rect 43700 9090 43720 9130
rect 43640 9060 43720 9090
rect 43750 9230 43830 9260
rect 43750 9190 43770 9230
rect 43810 9190 43830 9230
rect 43750 9130 43830 9190
rect 43750 9090 43770 9130
rect 43810 9090 43830 9130
rect 43750 9060 43830 9090
rect 43860 9230 43940 9260
rect 43860 9190 43880 9230
rect 43920 9190 43940 9230
rect 43860 9130 43940 9190
rect 43860 9090 43880 9130
rect 43920 9090 43940 9130
rect 43860 9060 43940 9090
rect 43970 9230 44050 9260
rect 43970 9190 43990 9230
rect 44030 9190 44050 9230
rect 43970 9130 44050 9190
rect 43970 9090 43990 9130
rect 44030 9090 44050 9130
rect 43970 9060 44050 9090
rect 44080 9230 44160 9260
rect 44080 9190 44100 9230
rect 44140 9190 44160 9230
rect 44080 9130 44160 9190
rect 44080 9090 44100 9130
rect 44140 9090 44160 9130
rect 44080 9060 44160 9090
rect 44190 9230 44270 9260
rect 44190 9190 44210 9230
rect 44250 9190 44270 9230
rect 44190 9130 44270 9190
rect 44190 9090 44210 9130
rect 44250 9090 44270 9130
rect 44190 9060 44270 9090
rect 44300 9230 44380 9260
rect 44300 9190 44320 9230
rect 44360 9190 44380 9230
rect 44300 9130 44380 9190
rect 44300 9090 44320 9130
rect 44360 9090 44380 9130
rect 44300 9060 44380 9090
rect 44410 9230 44490 9260
rect 44410 9190 44430 9230
rect 44470 9190 44490 9230
rect 44410 9130 44490 9190
rect 44410 9090 44430 9130
rect 44470 9090 44490 9130
rect 44410 9060 44490 9090
rect 44520 9230 44600 9260
rect 44520 9190 44540 9230
rect 44580 9190 44600 9230
rect 44520 9130 44600 9190
rect 44520 9090 44540 9130
rect 44580 9090 44600 9130
rect 44520 9060 44600 9090
rect 44630 9230 44710 9260
rect 44630 9190 44650 9230
rect 44690 9190 44710 9230
rect 44630 9130 44710 9190
rect 44630 9090 44650 9130
rect 44690 9090 44710 9130
rect 44630 9060 44710 9090
rect 44740 9230 44820 9260
rect 44740 9190 44760 9230
rect 44800 9190 44820 9230
rect 44740 9130 44820 9190
rect 44740 9090 44760 9130
rect 44800 9090 44820 9130
rect 44740 9060 44820 9090
rect 44850 9230 44930 9260
rect 44850 9190 44870 9230
rect 44910 9190 44930 9230
rect 44850 9130 44930 9190
rect 44850 9090 44870 9130
rect 44910 9090 44930 9130
rect 44850 9060 44930 9090
<< ndiffc >>
rect 41180 13810 41220 13850
rect 41180 13710 41220 13750
rect 43260 13810 43300 13850
rect 43260 13710 43300 13750
rect 45340 13810 45380 13850
rect 45340 13710 45380 13750
rect 40760 13200 40800 13240
rect 40760 13100 40800 13140
rect 40760 13000 40800 13040
rect 40760 12900 40800 12940
rect 40760 12800 40800 12840
rect 41840 13200 41880 13240
rect 42000 13200 42040 13240
rect 41840 13100 41880 13140
rect 42000 13100 42040 13140
rect 41840 13000 41880 13040
rect 42000 13000 42040 13040
rect 41840 12900 41880 12940
rect 42000 12900 42040 12940
rect 41840 12800 41880 12840
rect 42000 12800 42040 12840
rect 43080 13200 43120 13240
rect 43080 13100 43120 13140
rect 43080 13000 43120 13040
rect 43080 12900 43120 12940
rect 43080 12800 43120 12840
rect 43440 13200 43480 13240
rect 43440 13100 43480 13140
rect 43440 13000 43480 13040
rect 43440 12900 43480 12940
rect 43440 12800 43480 12840
rect 44520 13200 44560 13240
rect 44680 13200 44720 13240
rect 44520 13100 44560 13140
rect 44680 13100 44720 13140
rect 44520 13000 44560 13040
rect 44680 13000 44720 13040
rect 44520 12900 44560 12940
rect 44680 12900 44720 12940
rect 44520 12800 44560 12840
rect 44680 12800 44720 12840
rect 45760 13200 45800 13240
rect 45760 13100 45800 13140
rect 45760 13000 45800 13040
rect 45760 12900 45800 12940
rect 45760 12800 45800 12840
rect 41380 12190 41420 12230
rect 41500 12190 41540 12230
rect 41620 12190 41660 12230
rect 41740 12190 41780 12230
rect 41860 12190 41900 12230
rect 41980 12190 42020 12230
rect 42100 12190 42140 12230
rect 42220 12190 42260 12230
rect 42340 12190 42380 12230
rect 42460 12190 42500 12230
rect 42580 12190 42620 12230
rect 43940 12190 43980 12230
rect 44060 12190 44100 12230
rect 44180 12190 44220 12230
rect 44300 12190 44340 12230
rect 44420 12190 44460 12230
rect 44540 12190 44580 12230
rect 44660 12190 44700 12230
rect 44780 12190 44820 12230
rect 44900 12190 44940 12230
rect 45020 12190 45060 12230
rect 45140 12190 45180 12230
<< pdiffc >>
rect 41632 18392 41666 18426
rect 41722 18392 41756 18426
rect 41812 18392 41846 18426
rect 41902 18392 41936 18426
rect 41992 18392 42026 18426
rect 42082 18392 42116 18426
rect 42172 18392 42206 18426
rect 41632 18302 41666 18336
rect 41722 18302 41756 18336
rect 41812 18302 41846 18336
rect 41902 18302 41936 18336
rect 41992 18302 42026 18336
rect 42082 18302 42116 18336
rect 42172 18302 42206 18336
rect 41632 18212 41666 18246
rect 41722 18212 41756 18246
rect 41812 18212 41846 18246
rect 41902 18212 41936 18246
rect 41992 18212 42026 18246
rect 42082 18212 42116 18246
rect 42172 18212 42206 18246
rect 41632 18122 41666 18156
rect 41722 18122 41756 18156
rect 41812 18122 41846 18156
rect 41902 18122 41936 18156
rect 41992 18122 42026 18156
rect 42082 18122 42116 18156
rect 42172 18122 42206 18156
rect 41632 18032 41666 18066
rect 41722 18032 41756 18066
rect 41812 18032 41846 18066
rect 41902 18032 41936 18066
rect 41992 18032 42026 18066
rect 42082 18032 42116 18066
rect 42172 18032 42206 18066
rect 41632 17942 41666 17976
rect 41722 17942 41756 17976
rect 41812 17942 41846 17976
rect 41902 17942 41936 17976
rect 41992 17942 42026 17976
rect 42082 17942 42116 17976
rect 42172 17942 42206 17976
rect 41632 17852 41666 17886
rect 41722 17852 41756 17886
rect 41812 17852 41846 17886
rect 41902 17852 41936 17886
rect 41992 17852 42026 17886
rect 42082 17852 42116 17886
rect 42172 17852 42206 17886
rect 42992 18392 43026 18426
rect 43082 18392 43116 18426
rect 43172 18392 43206 18426
rect 43262 18392 43296 18426
rect 43352 18392 43386 18426
rect 43442 18392 43476 18426
rect 43532 18392 43566 18426
rect 42992 18302 43026 18336
rect 43082 18302 43116 18336
rect 43172 18302 43206 18336
rect 43262 18302 43296 18336
rect 43352 18302 43386 18336
rect 43442 18302 43476 18336
rect 43532 18302 43566 18336
rect 42992 18212 43026 18246
rect 43082 18212 43116 18246
rect 43172 18212 43206 18246
rect 43262 18212 43296 18246
rect 43352 18212 43386 18246
rect 43442 18212 43476 18246
rect 43532 18212 43566 18246
rect 42992 18122 43026 18156
rect 43082 18122 43116 18156
rect 43172 18122 43206 18156
rect 43262 18122 43296 18156
rect 43352 18122 43386 18156
rect 43442 18122 43476 18156
rect 43532 18122 43566 18156
rect 42992 18032 43026 18066
rect 43082 18032 43116 18066
rect 43172 18032 43206 18066
rect 43262 18032 43296 18066
rect 43352 18032 43386 18066
rect 43442 18032 43476 18066
rect 43532 18032 43566 18066
rect 42992 17942 43026 17976
rect 43082 17942 43116 17976
rect 43172 17942 43206 17976
rect 43262 17942 43296 17976
rect 43352 17942 43386 17976
rect 43442 17942 43476 17976
rect 43532 17942 43566 17976
rect 42992 17852 43026 17886
rect 43082 17852 43116 17886
rect 43172 17852 43206 17886
rect 43262 17852 43296 17886
rect 43352 17852 43386 17886
rect 43442 17852 43476 17886
rect 43532 17852 43566 17886
rect 44352 18392 44386 18426
rect 44442 18392 44476 18426
rect 44532 18392 44566 18426
rect 44622 18392 44656 18426
rect 44712 18392 44746 18426
rect 44802 18392 44836 18426
rect 44892 18392 44926 18426
rect 44352 18302 44386 18336
rect 44442 18302 44476 18336
rect 44532 18302 44566 18336
rect 44622 18302 44656 18336
rect 44712 18302 44746 18336
rect 44802 18302 44836 18336
rect 44892 18302 44926 18336
rect 44352 18212 44386 18246
rect 44442 18212 44476 18246
rect 44532 18212 44566 18246
rect 44622 18212 44656 18246
rect 44712 18212 44746 18246
rect 44802 18212 44836 18246
rect 44892 18212 44926 18246
rect 44352 18122 44386 18156
rect 44442 18122 44476 18156
rect 44532 18122 44566 18156
rect 44622 18122 44656 18156
rect 44712 18122 44746 18156
rect 44802 18122 44836 18156
rect 44892 18122 44926 18156
rect 44352 18032 44386 18066
rect 44442 18032 44476 18066
rect 44532 18032 44566 18066
rect 44622 18032 44656 18066
rect 44712 18032 44746 18066
rect 44802 18032 44836 18066
rect 44892 18032 44926 18066
rect 44352 17942 44386 17976
rect 44442 17942 44476 17976
rect 44532 17942 44566 17976
rect 44622 17942 44656 17976
rect 44712 17942 44746 17976
rect 44802 17942 44836 17976
rect 44892 17942 44926 17976
rect 44352 17852 44386 17886
rect 44442 17852 44476 17886
rect 44532 17852 44566 17886
rect 44622 17852 44656 17886
rect 44712 17852 44746 17886
rect 44802 17852 44836 17886
rect 44892 17852 44926 17886
rect 41632 17032 41666 17066
rect 41722 17032 41756 17066
rect 41812 17032 41846 17066
rect 41902 17032 41936 17066
rect 41992 17032 42026 17066
rect 42082 17032 42116 17066
rect 42172 17032 42206 17066
rect 41632 16942 41666 16976
rect 41722 16942 41756 16976
rect 41812 16942 41846 16976
rect 41902 16942 41936 16976
rect 41992 16942 42026 16976
rect 42082 16942 42116 16976
rect 42172 16942 42206 16976
rect 41632 16852 41666 16886
rect 41722 16852 41756 16886
rect 41812 16852 41846 16886
rect 41902 16852 41936 16886
rect 41992 16852 42026 16886
rect 42082 16852 42116 16886
rect 42172 16852 42206 16886
rect 41632 16762 41666 16796
rect 41722 16762 41756 16796
rect 41812 16762 41846 16796
rect 41902 16762 41936 16796
rect 41992 16762 42026 16796
rect 42082 16762 42116 16796
rect 42172 16762 42206 16796
rect 41632 16672 41666 16706
rect 41722 16672 41756 16706
rect 41812 16672 41846 16706
rect 41902 16672 41936 16706
rect 41992 16672 42026 16706
rect 42082 16672 42116 16706
rect 42172 16672 42206 16706
rect 41632 16582 41666 16616
rect 41722 16582 41756 16616
rect 41812 16582 41846 16616
rect 41902 16582 41936 16616
rect 41992 16582 42026 16616
rect 42082 16582 42116 16616
rect 42172 16582 42206 16616
rect 41632 16492 41666 16526
rect 41722 16492 41756 16526
rect 41812 16492 41846 16526
rect 41902 16492 41936 16526
rect 41992 16492 42026 16526
rect 42082 16492 42116 16526
rect 42172 16492 42206 16526
rect 42992 17032 43026 17066
rect 43082 17032 43116 17066
rect 43172 17032 43206 17066
rect 43262 17032 43296 17066
rect 43352 17032 43386 17066
rect 43442 17032 43476 17066
rect 43532 17032 43566 17066
rect 42992 16942 43026 16976
rect 43082 16942 43116 16976
rect 43172 16942 43206 16976
rect 43262 16942 43296 16976
rect 43352 16942 43386 16976
rect 43442 16942 43476 16976
rect 43532 16942 43566 16976
rect 42992 16852 43026 16886
rect 43082 16852 43116 16886
rect 43172 16852 43206 16886
rect 43262 16852 43296 16886
rect 43352 16852 43386 16886
rect 43442 16852 43476 16886
rect 43532 16852 43566 16886
rect 42992 16762 43026 16796
rect 43082 16762 43116 16796
rect 43172 16762 43206 16796
rect 43262 16762 43296 16796
rect 43352 16762 43386 16796
rect 43442 16762 43476 16796
rect 43532 16762 43566 16796
rect 42992 16672 43026 16706
rect 43082 16672 43116 16706
rect 43172 16672 43206 16706
rect 43262 16672 43296 16706
rect 43352 16672 43386 16706
rect 43442 16672 43476 16706
rect 43532 16672 43566 16706
rect 42992 16582 43026 16616
rect 43082 16582 43116 16616
rect 43172 16582 43206 16616
rect 43262 16582 43296 16616
rect 43352 16582 43386 16616
rect 43442 16582 43476 16616
rect 43532 16582 43566 16616
rect 42992 16492 43026 16526
rect 43082 16492 43116 16526
rect 43172 16492 43206 16526
rect 43262 16492 43296 16526
rect 43352 16492 43386 16526
rect 43442 16492 43476 16526
rect 43532 16492 43566 16526
rect 44352 17032 44386 17066
rect 44442 17032 44476 17066
rect 44532 17032 44566 17066
rect 44622 17032 44656 17066
rect 44712 17032 44746 17066
rect 44802 17032 44836 17066
rect 44892 17032 44926 17066
rect 44352 16942 44386 16976
rect 44442 16942 44476 16976
rect 44532 16942 44566 16976
rect 44622 16942 44656 16976
rect 44712 16942 44746 16976
rect 44802 16942 44836 16976
rect 44892 16942 44926 16976
rect 44352 16852 44386 16886
rect 44442 16852 44476 16886
rect 44532 16852 44566 16886
rect 44622 16852 44656 16886
rect 44712 16852 44746 16886
rect 44802 16852 44836 16886
rect 44892 16852 44926 16886
rect 44352 16762 44386 16796
rect 44442 16762 44476 16796
rect 44532 16762 44566 16796
rect 44622 16762 44656 16796
rect 44712 16762 44746 16796
rect 44802 16762 44836 16796
rect 44892 16762 44926 16796
rect 44352 16672 44386 16706
rect 44442 16672 44476 16706
rect 44532 16672 44566 16706
rect 44622 16672 44656 16706
rect 44712 16672 44746 16706
rect 44802 16672 44836 16706
rect 44892 16672 44926 16706
rect 44352 16582 44386 16616
rect 44442 16582 44476 16616
rect 44532 16582 44566 16616
rect 44622 16582 44656 16616
rect 44712 16582 44746 16616
rect 44802 16582 44836 16616
rect 44892 16582 44926 16616
rect 44352 16492 44386 16526
rect 44442 16492 44476 16526
rect 44532 16492 44566 16526
rect 44622 16492 44656 16526
rect 44712 16492 44746 16526
rect 44802 16492 44836 16526
rect 44892 16492 44926 16526
rect 41632 15672 41666 15706
rect 41722 15672 41756 15706
rect 41812 15672 41846 15706
rect 41902 15672 41936 15706
rect 41992 15672 42026 15706
rect 42082 15672 42116 15706
rect 42172 15672 42206 15706
rect 41632 15582 41666 15616
rect 41722 15582 41756 15616
rect 41812 15582 41846 15616
rect 41902 15582 41936 15616
rect 41992 15582 42026 15616
rect 42082 15582 42116 15616
rect 42172 15582 42206 15616
rect 41632 15492 41666 15526
rect 41722 15492 41756 15526
rect 41812 15492 41846 15526
rect 41902 15492 41936 15526
rect 41992 15492 42026 15526
rect 42082 15492 42116 15526
rect 42172 15492 42206 15526
rect 41632 15402 41666 15436
rect 41722 15402 41756 15436
rect 41812 15402 41846 15436
rect 41902 15402 41936 15436
rect 41992 15402 42026 15436
rect 42082 15402 42116 15436
rect 42172 15402 42206 15436
rect 41632 15312 41666 15346
rect 41722 15312 41756 15346
rect 41812 15312 41846 15346
rect 41902 15312 41936 15346
rect 41992 15312 42026 15346
rect 42082 15312 42116 15346
rect 42172 15312 42206 15346
rect 41632 15222 41666 15256
rect 41722 15222 41756 15256
rect 41812 15222 41846 15256
rect 41902 15222 41936 15256
rect 41992 15222 42026 15256
rect 42082 15222 42116 15256
rect 42172 15222 42206 15256
rect 41632 15132 41666 15166
rect 41722 15132 41756 15166
rect 41812 15132 41846 15166
rect 41902 15132 41936 15166
rect 41992 15132 42026 15166
rect 42082 15132 42116 15166
rect 42172 15132 42206 15166
rect 42992 15672 43026 15706
rect 43082 15672 43116 15706
rect 43172 15672 43206 15706
rect 43262 15672 43296 15706
rect 43352 15672 43386 15706
rect 43442 15672 43476 15706
rect 43532 15672 43566 15706
rect 42992 15582 43026 15616
rect 43082 15582 43116 15616
rect 43172 15582 43206 15616
rect 43262 15582 43296 15616
rect 43352 15582 43386 15616
rect 43442 15582 43476 15616
rect 43532 15582 43566 15616
rect 42992 15492 43026 15526
rect 43082 15492 43116 15526
rect 43172 15492 43206 15526
rect 43262 15492 43296 15526
rect 43352 15492 43386 15526
rect 43442 15492 43476 15526
rect 43532 15492 43566 15526
rect 42992 15402 43026 15436
rect 43082 15402 43116 15436
rect 43172 15402 43206 15436
rect 43262 15402 43296 15436
rect 43352 15402 43386 15436
rect 43442 15402 43476 15436
rect 43532 15402 43566 15436
rect 42992 15312 43026 15346
rect 43082 15312 43116 15346
rect 43172 15312 43206 15346
rect 43262 15312 43296 15346
rect 43352 15312 43386 15346
rect 43442 15312 43476 15346
rect 43532 15312 43566 15346
rect 42992 15222 43026 15256
rect 43082 15222 43116 15256
rect 43172 15222 43206 15256
rect 43262 15222 43296 15256
rect 43352 15222 43386 15256
rect 43442 15222 43476 15256
rect 43532 15222 43566 15256
rect 42992 15132 43026 15166
rect 43082 15132 43116 15166
rect 43172 15132 43206 15166
rect 43262 15132 43296 15166
rect 43352 15132 43386 15166
rect 43442 15132 43476 15166
rect 43532 15132 43566 15166
rect 44352 15672 44386 15706
rect 44442 15672 44476 15706
rect 44532 15672 44566 15706
rect 44622 15672 44656 15706
rect 44712 15672 44746 15706
rect 44802 15672 44836 15706
rect 44892 15672 44926 15706
rect 44352 15582 44386 15616
rect 44442 15582 44476 15616
rect 44532 15582 44566 15616
rect 44622 15582 44656 15616
rect 44712 15582 44746 15616
rect 44802 15582 44836 15616
rect 44892 15582 44926 15616
rect 44352 15492 44386 15526
rect 44442 15492 44476 15526
rect 44532 15492 44566 15526
rect 44622 15492 44656 15526
rect 44712 15492 44746 15526
rect 44802 15492 44836 15526
rect 44892 15492 44926 15526
rect 44352 15402 44386 15436
rect 44442 15402 44476 15436
rect 44532 15402 44566 15436
rect 44622 15402 44656 15436
rect 44712 15402 44746 15436
rect 44802 15402 44836 15436
rect 44892 15402 44926 15436
rect 44352 15312 44386 15346
rect 44442 15312 44476 15346
rect 44532 15312 44566 15346
rect 44622 15312 44656 15346
rect 44712 15312 44746 15346
rect 44802 15312 44836 15346
rect 44892 15312 44926 15346
rect 44352 15222 44386 15256
rect 44442 15222 44476 15256
rect 44532 15222 44566 15256
rect 44622 15222 44656 15256
rect 44712 15222 44746 15256
rect 44802 15222 44836 15256
rect 44892 15222 44926 15256
rect 44352 15132 44386 15166
rect 44442 15132 44476 15166
rect 44532 15132 44566 15166
rect 44622 15132 44656 15166
rect 44712 15132 44746 15166
rect 44802 15132 44836 15166
rect 44892 15132 44926 15166
rect 40540 11350 40580 11390
rect 40540 11250 40580 11290
rect 40660 11350 40700 11390
rect 40660 11250 40700 11290
rect 40780 11350 40820 11390
rect 40780 11250 40820 11290
rect 40900 11350 40940 11390
rect 40900 11250 40940 11290
rect 41020 11350 41060 11390
rect 41020 11250 41060 11290
rect 41140 11350 41180 11390
rect 41140 11250 41180 11290
rect 41260 11350 41300 11390
rect 41260 11250 41300 11290
rect 41380 11350 41420 11390
rect 41380 11250 41420 11290
rect 41500 11350 41540 11390
rect 41500 11250 41540 11290
rect 41620 11350 41660 11390
rect 41620 11250 41660 11290
rect 41740 11350 41780 11390
rect 41740 11250 41780 11290
rect 41860 11350 41900 11390
rect 41860 11250 41900 11290
rect 41980 11350 42020 11390
rect 41980 11250 42020 11290
rect 42100 11350 42140 11390
rect 42100 11250 42140 11290
rect 42220 11350 42260 11390
rect 42220 11250 42260 11290
rect 42340 11350 42380 11390
rect 42340 11250 42380 11290
rect 42460 11350 42500 11390
rect 42460 11250 42500 11290
rect 42580 11350 42620 11390
rect 42580 11250 42620 11290
rect 42700 11350 42740 11390
rect 42700 11250 42740 11290
rect 42820 11350 42860 11390
rect 42820 11250 42860 11290
rect 42940 11350 42980 11390
rect 42940 11250 42980 11290
rect 43580 11350 43620 11390
rect 43580 11250 43620 11290
rect 43700 11350 43740 11390
rect 43700 11250 43740 11290
rect 43820 11350 43860 11390
rect 43820 11250 43860 11290
rect 43940 11350 43980 11390
rect 43940 11250 43980 11290
rect 44060 11350 44100 11390
rect 44060 11250 44100 11290
rect 44180 11350 44220 11390
rect 44180 11250 44220 11290
rect 44300 11350 44340 11390
rect 44300 11250 44340 11290
rect 44420 11350 44460 11390
rect 44420 11250 44460 11290
rect 44540 11350 44580 11390
rect 44540 11250 44580 11290
rect 44660 11350 44700 11390
rect 44660 11250 44700 11290
rect 44780 11350 44820 11390
rect 44780 11250 44820 11290
rect 44900 11350 44940 11390
rect 44900 11250 44940 11290
rect 45020 11350 45060 11390
rect 45020 11250 45060 11290
rect 45140 11350 45180 11390
rect 45140 11250 45180 11290
rect 45260 11350 45300 11390
rect 45260 11250 45300 11290
rect 45380 11350 45420 11390
rect 45380 11250 45420 11290
rect 45500 11350 45540 11390
rect 45500 11250 45540 11290
rect 45620 11350 45660 11390
rect 45620 11250 45660 11290
rect 45740 11350 45780 11390
rect 45740 11250 45780 11290
rect 45860 11350 45900 11390
rect 45860 11250 45900 11290
rect 45980 11350 46020 11390
rect 45980 11250 46020 11290
rect 41640 10190 41680 10230
rect 41640 10090 41680 10130
rect 41640 9990 41680 10030
rect 41640 9890 41680 9930
rect 41640 9790 41680 9830
rect 41640 9690 41680 9730
rect 41820 10190 41860 10230
rect 41820 10090 41860 10130
rect 41820 9990 41860 10030
rect 41820 9890 41860 9930
rect 41820 9790 41860 9830
rect 41820 9690 41860 9730
rect 42000 10190 42040 10230
rect 42000 10090 42040 10130
rect 42000 9990 42040 10030
rect 42000 9890 42040 9930
rect 42000 9790 42040 9830
rect 42000 9690 42040 9730
rect 42180 10190 42220 10230
rect 42180 10090 42220 10130
rect 42180 9990 42220 10030
rect 42180 9890 42220 9930
rect 42180 9790 42220 9830
rect 42180 9690 42220 9730
rect 42360 10190 42400 10230
rect 42360 10090 42400 10130
rect 42360 9990 42400 10030
rect 42360 9890 42400 9930
rect 42360 9790 42400 9830
rect 42360 9690 42400 9730
rect 42540 10190 42580 10230
rect 42540 10090 42580 10130
rect 42540 9990 42580 10030
rect 42540 9890 42580 9930
rect 42540 9790 42580 9830
rect 42540 9690 42580 9730
rect 42720 10190 42760 10230
rect 42720 10090 42760 10130
rect 42720 9990 42760 10030
rect 42720 9890 42760 9930
rect 42720 9790 42760 9830
rect 42720 9690 42760 9730
rect 42900 10190 42940 10230
rect 42900 10090 42940 10130
rect 42900 9990 42940 10030
rect 42900 9890 42940 9930
rect 42900 9790 42940 9830
rect 42900 9690 42940 9730
rect 43080 10190 43120 10230
rect 43080 10090 43120 10130
rect 43080 9990 43120 10030
rect 43080 9890 43120 9930
rect 43080 9790 43120 9830
rect 43080 9690 43120 9730
rect 43260 10190 43300 10230
rect 43260 10090 43300 10130
rect 43260 9990 43300 10030
rect 43260 9890 43300 9930
rect 43260 9790 43300 9830
rect 43260 9690 43300 9730
rect 43440 10190 43480 10230
rect 43440 10090 43480 10130
rect 43440 9990 43480 10030
rect 43440 9890 43480 9930
rect 43440 9790 43480 9830
rect 43440 9690 43480 9730
rect 43620 10190 43660 10230
rect 43620 10090 43660 10130
rect 43620 9990 43660 10030
rect 43620 9890 43660 9930
rect 43620 9790 43660 9830
rect 43620 9690 43660 9730
rect 43800 10190 43840 10230
rect 43800 10090 43840 10130
rect 43800 9990 43840 10030
rect 43800 9890 43840 9930
rect 43800 9790 43840 9830
rect 43800 9690 43840 9730
rect 43980 10190 44020 10230
rect 43980 10090 44020 10130
rect 43980 9990 44020 10030
rect 43980 9890 44020 9930
rect 43980 9790 44020 9830
rect 43980 9690 44020 9730
rect 44160 10190 44200 10230
rect 44160 10090 44200 10130
rect 44160 9990 44200 10030
rect 44160 9890 44200 9930
rect 44160 9790 44200 9830
rect 44160 9690 44200 9730
rect 44340 10190 44380 10230
rect 44340 10090 44380 10130
rect 44340 9990 44380 10030
rect 44340 9890 44380 9930
rect 44340 9790 44380 9830
rect 44340 9690 44380 9730
rect 44520 10190 44560 10230
rect 44520 10090 44560 10130
rect 44520 9990 44560 10030
rect 44520 9890 44560 9930
rect 44520 9790 44560 9830
rect 44520 9690 44560 9730
rect 44700 10190 44740 10230
rect 44700 10090 44740 10130
rect 44700 9990 44740 10030
rect 44700 9890 44740 9930
rect 44700 9790 44740 9830
rect 44700 9690 44740 9730
rect 44880 10190 44920 10230
rect 44880 10090 44920 10130
rect 44880 9990 44920 10030
rect 44880 9890 44920 9930
rect 45510 9990 45550 10030
rect 45510 9890 45550 9930
rect 45620 9990 45660 10030
rect 45620 9890 45660 9930
rect 45730 9990 45770 10030
rect 45730 9890 45770 9930
rect 45840 9990 45880 10030
rect 45840 9890 45880 9930
rect 45950 9990 45990 10030
rect 45950 9890 45990 9930
rect 44880 9790 44920 9830
rect 44880 9690 44920 9730
rect 41650 9190 41690 9230
rect 41650 9090 41690 9130
rect 41760 9190 41800 9230
rect 41760 9090 41800 9130
rect 41870 9190 41910 9230
rect 41870 9090 41910 9130
rect 41980 9190 42020 9230
rect 41980 9090 42020 9130
rect 42090 9190 42130 9230
rect 42090 9090 42130 9130
rect 42200 9190 42240 9230
rect 42200 9090 42240 9130
rect 42310 9190 42350 9230
rect 42310 9090 42350 9130
rect 42420 9190 42460 9230
rect 42420 9090 42460 9130
rect 42530 9190 42570 9230
rect 42530 9090 42570 9130
rect 42640 9190 42680 9230
rect 42640 9090 42680 9130
rect 42750 9190 42790 9230
rect 42750 9090 42790 9130
rect 42860 9190 42900 9230
rect 42860 9090 42900 9130
rect 42970 9190 43010 9230
rect 42970 9090 43010 9130
rect 43550 9190 43590 9230
rect 43550 9090 43590 9130
rect 43660 9190 43700 9230
rect 43660 9090 43700 9130
rect 43770 9190 43810 9230
rect 43770 9090 43810 9130
rect 43880 9190 43920 9230
rect 43880 9090 43920 9130
rect 43990 9190 44030 9230
rect 43990 9090 44030 9130
rect 44100 9190 44140 9230
rect 44100 9090 44140 9130
rect 44210 9190 44250 9230
rect 44210 9090 44250 9130
rect 44320 9190 44360 9230
rect 44320 9090 44360 9130
rect 44430 9190 44470 9230
rect 44430 9090 44470 9130
rect 44540 9190 44580 9230
rect 44540 9090 44580 9130
rect 44650 9190 44690 9230
rect 44650 9090 44690 9130
rect 44760 9190 44800 9230
rect 44760 9090 44800 9130
rect 44870 9190 44910 9230
rect 44870 9090 44910 9130
<< psubdiff >>
rect 43230 19070 43330 19100
rect 43230 19030 43260 19070
rect 43300 19030 43330 19070
rect 43230 18990 43330 19030
rect 43230 18950 43260 18990
rect 43300 18950 43330 18990
rect 43230 18910 43330 18950
rect 43230 18870 43260 18910
rect 43300 18870 43330 18910
rect 43230 18840 43330 18870
rect 41276 18752 42564 18784
rect 41276 18718 41410 18752
rect 41444 18718 41500 18752
rect 41534 18718 41590 18752
rect 41624 18718 41680 18752
rect 41714 18718 41770 18752
rect 41804 18718 41860 18752
rect 41894 18718 41950 18752
rect 41984 18718 42040 18752
rect 42074 18718 42130 18752
rect 42164 18718 42220 18752
rect 42254 18718 42310 18752
rect 42344 18718 42400 18752
rect 42434 18718 42564 18752
rect 41276 18683 42564 18718
rect 41276 18668 41377 18683
rect 41276 18634 41309 18668
rect 41343 18634 41377 18668
rect 41276 18578 41377 18634
rect 42463 18668 42564 18683
rect 42463 18634 42496 18668
rect 42530 18634 42564 18668
rect 41276 18544 41309 18578
rect 41343 18544 41377 18578
rect 41276 18488 41377 18544
rect 41276 18454 41309 18488
rect 41343 18454 41377 18488
rect 41276 18398 41377 18454
rect 41276 18364 41309 18398
rect 41343 18364 41377 18398
rect 41276 18308 41377 18364
rect 41276 18274 41309 18308
rect 41343 18274 41377 18308
rect 41276 18218 41377 18274
rect 41276 18184 41309 18218
rect 41343 18184 41377 18218
rect 41276 18128 41377 18184
rect 41276 18094 41309 18128
rect 41343 18094 41377 18128
rect 41276 18038 41377 18094
rect 41276 18004 41309 18038
rect 41343 18004 41377 18038
rect 41276 17948 41377 18004
rect 41276 17914 41309 17948
rect 41343 17914 41377 17948
rect 41276 17858 41377 17914
rect 41276 17824 41309 17858
rect 41343 17824 41377 17858
rect 41276 17768 41377 17824
rect 41276 17734 41309 17768
rect 41343 17734 41377 17768
rect 41276 17678 41377 17734
rect 41276 17644 41309 17678
rect 41343 17644 41377 17678
rect 42463 18578 42564 18634
rect 42463 18544 42496 18578
rect 42530 18544 42564 18578
rect 42463 18488 42564 18544
rect 42463 18454 42496 18488
rect 42530 18454 42564 18488
rect 42463 18398 42564 18454
rect 42463 18364 42496 18398
rect 42530 18364 42564 18398
rect 42463 18308 42564 18364
rect 42463 18274 42496 18308
rect 42530 18274 42564 18308
rect 42463 18218 42564 18274
rect 42463 18184 42496 18218
rect 42530 18184 42564 18218
rect 42463 18128 42564 18184
rect 42463 18094 42496 18128
rect 42530 18094 42564 18128
rect 42463 18038 42564 18094
rect 42463 18004 42496 18038
rect 42530 18004 42564 18038
rect 42463 17948 42564 18004
rect 42463 17914 42496 17948
rect 42530 17914 42564 17948
rect 42463 17858 42564 17914
rect 42463 17824 42496 17858
rect 42530 17824 42564 17858
rect 42463 17768 42564 17824
rect 42463 17734 42496 17768
rect 42530 17734 42564 17768
rect 42463 17678 42564 17734
rect 41276 17597 41377 17644
rect 42463 17644 42496 17678
rect 42530 17644 42564 17678
rect 42463 17597 42564 17644
rect 41276 17588 42564 17597
rect 41276 17554 41309 17588
rect 41343 17565 42496 17588
rect 41343 17554 41410 17565
rect 41276 17531 41410 17554
rect 41444 17531 41500 17565
rect 41534 17531 41590 17565
rect 41624 17531 41680 17565
rect 41714 17531 41770 17565
rect 41804 17531 41860 17565
rect 41894 17531 41950 17565
rect 41984 17531 42040 17565
rect 42074 17531 42130 17565
rect 42164 17531 42220 17565
rect 42254 17531 42310 17565
rect 42344 17531 42400 17565
rect 42434 17554 42496 17565
rect 42530 17554 42564 17588
rect 42434 17531 42564 17554
rect 41276 17496 42564 17531
rect 42636 18752 43924 18784
rect 42636 18718 42770 18752
rect 42804 18718 42860 18752
rect 42894 18718 42950 18752
rect 42984 18718 43040 18752
rect 43074 18718 43130 18752
rect 43164 18718 43220 18752
rect 43254 18718 43310 18752
rect 43344 18718 43400 18752
rect 43434 18718 43490 18752
rect 43524 18718 43580 18752
rect 43614 18718 43670 18752
rect 43704 18718 43760 18752
rect 43794 18718 43924 18752
rect 42636 18683 43924 18718
rect 42636 18668 42737 18683
rect 42636 18634 42669 18668
rect 42703 18634 42737 18668
rect 42636 18578 42737 18634
rect 43823 18668 43924 18683
rect 43823 18634 43856 18668
rect 43890 18634 43924 18668
rect 42636 18544 42669 18578
rect 42703 18544 42737 18578
rect 42636 18488 42737 18544
rect 42636 18454 42669 18488
rect 42703 18454 42737 18488
rect 42636 18398 42737 18454
rect 42636 18364 42669 18398
rect 42703 18364 42737 18398
rect 42636 18308 42737 18364
rect 42636 18274 42669 18308
rect 42703 18274 42737 18308
rect 42636 18218 42737 18274
rect 42636 18184 42669 18218
rect 42703 18184 42737 18218
rect 42636 18128 42737 18184
rect 42636 18094 42669 18128
rect 42703 18094 42737 18128
rect 42636 18038 42737 18094
rect 42636 18004 42669 18038
rect 42703 18004 42737 18038
rect 42636 17948 42737 18004
rect 42636 17914 42669 17948
rect 42703 17914 42737 17948
rect 42636 17858 42737 17914
rect 42636 17824 42669 17858
rect 42703 17824 42737 17858
rect 42636 17768 42737 17824
rect 42636 17734 42669 17768
rect 42703 17734 42737 17768
rect 42636 17678 42737 17734
rect 42636 17644 42669 17678
rect 42703 17644 42737 17678
rect 43823 18578 43924 18634
rect 43823 18544 43856 18578
rect 43890 18544 43924 18578
rect 43823 18488 43924 18544
rect 43823 18454 43856 18488
rect 43890 18454 43924 18488
rect 43823 18398 43924 18454
rect 43823 18364 43856 18398
rect 43890 18364 43924 18398
rect 43823 18308 43924 18364
rect 43823 18274 43856 18308
rect 43890 18274 43924 18308
rect 43823 18218 43924 18274
rect 43823 18184 43856 18218
rect 43890 18184 43924 18218
rect 43823 18128 43924 18184
rect 43823 18094 43856 18128
rect 43890 18094 43924 18128
rect 43823 18038 43924 18094
rect 43823 18004 43856 18038
rect 43890 18004 43924 18038
rect 43823 17948 43924 18004
rect 43823 17914 43856 17948
rect 43890 17914 43924 17948
rect 43823 17858 43924 17914
rect 43823 17824 43856 17858
rect 43890 17824 43924 17858
rect 43823 17768 43924 17824
rect 43823 17734 43856 17768
rect 43890 17734 43924 17768
rect 43823 17678 43924 17734
rect 42636 17597 42737 17644
rect 43823 17644 43856 17678
rect 43890 17644 43924 17678
rect 43823 17597 43924 17644
rect 42636 17588 43924 17597
rect 42636 17554 42669 17588
rect 42703 17565 43856 17588
rect 42703 17554 42770 17565
rect 42636 17531 42770 17554
rect 42804 17531 42860 17565
rect 42894 17531 42950 17565
rect 42984 17531 43040 17565
rect 43074 17531 43130 17565
rect 43164 17531 43220 17565
rect 43254 17531 43310 17565
rect 43344 17531 43400 17565
rect 43434 17531 43490 17565
rect 43524 17531 43580 17565
rect 43614 17531 43670 17565
rect 43704 17531 43760 17565
rect 43794 17554 43856 17565
rect 43890 17554 43924 17588
rect 43794 17531 43924 17554
rect 42636 17496 43924 17531
rect 43996 18752 45284 18784
rect 43996 18718 44130 18752
rect 44164 18718 44220 18752
rect 44254 18718 44310 18752
rect 44344 18718 44400 18752
rect 44434 18718 44490 18752
rect 44524 18718 44580 18752
rect 44614 18718 44670 18752
rect 44704 18718 44760 18752
rect 44794 18718 44850 18752
rect 44884 18718 44940 18752
rect 44974 18718 45030 18752
rect 45064 18718 45120 18752
rect 45154 18718 45284 18752
rect 43996 18683 45284 18718
rect 43996 18668 44097 18683
rect 43996 18634 44029 18668
rect 44063 18634 44097 18668
rect 43996 18578 44097 18634
rect 45183 18668 45284 18683
rect 45183 18634 45216 18668
rect 45250 18634 45284 18668
rect 43996 18544 44029 18578
rect 44063 18544 44097 18578
rect 43996 18488 44097 18544
rect 43996 18454 44029 18488
rect 44063 18454 44097 18488
rect 43996 18398 44097 18454
rect 43996 18364 44029 18398
rect 44063 18364 44097 18398
rect 43996 18308 44097 18364
rect 43996 18274 44029 18308
rect 44063 18274 44097 18308
rect 43996 18218 44097 18274
rect 43996 18184 44029 18218
rect 44063 18184 44097 18218
rect 43996 18128 44097 18184
rect 43996 18094 44029 18128
rect 44063 18094 44097 18128
rect 43996 18038 44097 18094
rect 43996 18004 44029 18038
rect 44063 18004 44097 18038
rect 43996 17948 44097 18004
rect 43996 17914 44029 17948
rect 44063 17914 44097 17948
rect 43996 17858 44097 17914
rect 43996 17824 44029 17858
rect 44063 17824 44097 17858
rect 43996 17768 44097 17824
rect 43996 17734 44029 17768
rect 44063 17734 44097 17768
rect 43996 17678 44097 17734
rect 43996 17644 44029 17678
rect 44063 17644 44097 17678
rect 45183 18578 45284 18634
rect 45183 18544 45216 18578
rect 45250 18544 45284 18578
rect 45183 18488 45284 18544
rect 45183 18454 45216 18488
rect 45250 18454 45284 18488
rect 45183 18398 45284 18454
rect 45183 18364 45216 18398
rect 45250 18364 45284 18398
rect 45183 18308 45284 18364
rect 45183 18274 45216 18308
rect 45250 18274 45284 18308
rect 45183 18218 45284 18274
rect 45183 18184 45216 18218
rect 45250 18184 45284 18218
rect 45183 18128 45284 18184
rect 45183 18094 45216 18128
rect 45250 18094 45284 18128
rect 45183 18038 45284 18094
rect 45183 18004 45216 18038
rect 45250 18004 45284 18038
rect 45183 17948 45284 18004
rect 45183 17914 45216 17948
rect 45250 17914 45284 17948
rect 45183 17858 45284 17914
rect 45183 17824 45216 17858
rect 45250 17824 45284 17858
rect 45183 17768 45284 17824
rect 45183 17734 45216 17768
rect 45250 17734 45284 17768
rect 45183 17678 45284 17734
rect 43996 17597 44097 17644
rect 45183 17644 45216 17678
rect 45250 17644 45284 17678
rect 45183 17597 45284 17644
rect 43996 17588 45284 17597
rect 43996 17554 44029 17588
rect 44063 17565 45216 17588
rect 44063 17554 44130 17565
rect 43996 17531 44130 17554
rect 44164 17531 44220 17565
rect 44254 17531 44310 17565
rect 44344 17531 44400 17565
rect 44434 17531 44490 17565
rect 44524 17531 44580 17565
rect 44614 17531 44670 17565
rect 44704 17531 44760 17565
rect 44794 17531 44850 17565
rect 44884 17531 44940 17565
rect 44974 17531 45030 17565
rect 45064 17531 45120 17565
rect 45154 17554 45216 17565
rect 45250 17554 45284 17588
rect 45154 17531 45284 17554
rect 43996 17496 45284 17531
rect 41276 17392 42564 17424
rect 41276 17358 41410 17392
rect 41444 17358 41500 17392
rect 41534 17358 41590 17392
rect 41624 17358 41680 17392
rect 41714 17358 41770 17392
rect 41804 17358 41860 17392
rect 41894 17358 41950 17392
rect 41984 17358 42040 17392
rect 42074 17358 42130 17392
rect 42164 17358 42220 17392
rect 42254 17358 42310 17392
rect 42344 17358 42400 17392
rect 42434 17358 42564 17392
rect 41276 17323 42564 17358
rect 41276 17308 41377 17323
rect 41276 17274 41309 17308
rect 41343 17274 41377 17308
rect 41276 17218 41377 17274
rect 42463 17308 42564 17323
rect 42463 17274 42496 17308
rect 42530 17274 42564 17308
rect 41276 17184 41309 17218
rect 41343 17184 41377 17218
rect 41276 17128 41377 17184
rect 41276 17094 41309 17128
rect 41343 17094 41377 17128
rect 41276 17038 41377 17094
rect 41276 17004 41309 17038
rect 41343 17004 41377 17038
rect 41276 16948 41377 17004
rect 41276 16914 41309 16948
rect 41343 16914 41377 16948
rect 41276 16858 41377 16914
rect 41276 16824 41309 16858
rect 41343 16824 41377 16858
rect 41276 16768 41377 16824
rect 41276 16734 41309 16768
rect 41343 16734 41377 16768
rect 41276 16678 41377 16734
rect 41276 16644 41309 16678
rect 41343 16644 41377 16678
rect 41276 16588 41377 16644
rect 41276 16554 41309 16588
rect 41343 16554 41377 16588
rect 41276 16498 41377 16554
rect 41276 16464 41309 16498
rect 41343 16464 41377 16498
rect 41276 16408 41377 16464
rect 41276 16374 41309 16408
rect 41343 16374 41377 16408
rect 41276 16318 41377 16374
rect 41276 16284 41309 16318
rect 41343 16284 41377 16318
rect 42463 17218 42564 17274
rect 42463 17184 42496 17218
rect 42530 17184 42564 17218
rect 42463 17128 42564 17184
rect 42463 17094 42496 17128
rect 42530 17094 42564 17128
rect 42463 17038 42564 17094
rect 42463 17004 42496 17038
rect 42530 17004 42564 17038
rect 42463 16948 42564 17004
rect 42463 16914 42496 16948
rect 42530 16914 42564 16948
rect 42463 16858 42564 16914
rect 42463 16824 42496 16858
rect 42530 16824 42564 16858
rect 42463 16768 42564 16824
rect 42463 16734 42496 16768
rect 42530 16734 42564 16768
rect 42463 16678 42564 16734
rect 42463 16644 42496 16678
rect 42530 16644 42564 16678
rect 42463 16588 42564 16644
rect 42463 16554 42496 16588
rect 42530 16554 42564 16588
rect 42463 16498 42564 16554
rect 42463 16464 42496 16498
rect 42530 16464 42564 16498
rect 42463 16408 42564 16464
rect 42463 16374 42496 16408
rect 42530 16374 42564 16408
rect 42463 16318 42564 16374
rect 41276 16237 41377 16284
rect 42463 16284 42496 16318
rect 42530 16284 42564 16318
rect 42463 16237 42564 16284
rect 41276 16228 42564 16237
rect 41276 16194 41309 16228
rect 41343 16205 42496 16228
rect 41343 16194 41410 16205
rect 41276 16171 41410 16194
rect 41444 16171 41500 16205
rect 41534 16171 41590 16205
rect 41624 16171 41680 16205
rect 41714 16171 41770 16205
rect 41804 16171 41860 16205
rect 41894 16171 41950 16205
rect 41984 16171 42040 16205
rect 42074 16171 42130 16205
rect 42164 16171 42220 16205
rect 42254 16171 42310 16205
rect 42344 16171 42400 16205
rect 42434 16194 42496 16205
rect 42530 16194 42564 16228
rect 42434 16171 42564 16194
rect 41276 16136 42564 16171
rect 42636 17392 43924 17424
rect 42636 17358 42770 17392
rect 42804 17358 42860 17392
rect 42894 17358 42950 17392
rect 42984 17358 43040 17392
rect 43074 17358 43130 17392
rect 43164 17358 43220 17392
rect 43254 17358 43310 17392
rect 43344 17358 43400 17392
rect 43434 17358 43490 17392
rect 43524 17358 43580 17392
rect 43614 17358 43670 17392
rect 43704 17358 43760 17392
rect 43794 17358 43924 17392
rect 42636 17323 43924 17358
rect 42636 17308 42737 17323
rect 42636 17274 42669 17308
rect 42703 17274 42737 17308
rect 42636 17218 42737 17274
rect 43823 17308 43924 17323
rect 43823 17274 43856 17308
rect 43890 17274 43924 17308
rect 42636 17184 42669 17218
rect 42703 17184 42737 17218
rect 42636 17128 42737 17184
rect 42636 17094 42669 17128
rect 42703 17094 42737 17128
rect 42636 17038 42737 17094
rect 42636 17004 42669 17038
rect 42703 17004 42737 17038
rect 42636 16948 42737 17004
rect 42636 16914 42669 16948
rect 42703 16914 42737 16948
rect 42636 16858 42737 16914
rect 42636 16824 42669 16858
rect 42703 16824 42737 16858
rect 42636 16768 42737 16824
rect 42636 16734 42669 16768
rect 42703 16734 42737 16768
rect 42636 16678 42737 16734
rect 42636 16644 42669 16678
rect 42703 16644 42737 16678
rect 42636 16588 42737 16644
rect 42636 16554 42669 16588
rect 42703 16554 42737 16588
rect 42636 16498 42737 16554
rect 42636 16464 42669 16498
rect 42703 16464 42737 16498
rect 42636 16408 42737 16464
rect 42636 16374 42669 16408
rect 42703 16374 42737 16408
rect 42636 16318 42737 16374
rect 42636 16284 42669 16318
rect 42703 16284 42737 16318
rect 43823 17218 43924 17274
rect 43823 17184 43856 17218
rect 43890 17184 43924 17218
rect 43823 17128 43924 17184
rect 43823 17094 43856 17128
rect 43890 17094 43924 17128
rect 43823 17038 43924 17094
rect 43823 17004 43856 17038
rect 43890 17004 43924 17038
rect 43823 16948 43924 17004
rect 43823 16914 43856 16948
rect 43890 16914 43924 16948
rect 43823 16858 43924 16914
rect 43823 16824 43856 16858
rect 43890 16824 43924 16858
rect 43823 16768 43924 16824
rect 43823 16734 43856 16768
rect 43890 16734 43924 16768
rect 43823 16678 43924 16734
rect 43823 16644 43856 16678
rect 43890 16644 43924 16678
rect 43823 16588 43924 16644
rect 43823 16554 43856 16588
rect 43890 16554 43924 16588
rect 43823 16498 43924 16554
rect 43823 16464 43856 16498
rect 43890 16464 43924 16498
rect 43823 16408 43924 16464
rect 43823 16374 43856 16408
rect 43890 16374 43924 16408
rect 43823 16318 43924 16374
rect 42636 16237 42737 16284
rect 43823 16284 43856 16318
rect 43890 16284 43924 16318
rect 43823 16237 43924 16284
rect 42636 16228 43924 16237
rect 42636 16194 42669 16228
rect 42703 16205 43856 16228
rect 42703 16194 42770 16205
rect 42636 16171 42770 16194
rect 42804 16171 42860 16205
rect 42894 16171 42950 16205
rect 42984 16171 43040 16205
rect 43074 16171 43130 16205
rect 43164 16171 43220 16205
rect 43254 16171 43310 16205
rect 43344 16171 43400 16205
rect 43434 16171 43490 16205
rect 43524 16171 43580 16205
rect 43614 16171 43670 16205
rect 43704 16171 43760 16205
rect 43794 16194 43856 16205
rect 43890 16194 43924 16228
rect 43794 16171 43924 16194
rect 42636 16136 43924 16171
rect 43996 17392 45284 17424
rect 43996 17358 44130 17392
rect 44164 17358 44220 17392
rect 44254 17358 44310 17392
rect 44344 17358 44400 17392
rect 44434 17358 44490 17392
rect 44524 17358 44580 17392
rect 44614 17358 44670 17392
rect 44704 17358 44760 17392
rect 44794 17358 44850 17392
rect 44884 17358 44940 17392
rect 44974 17358 45030 17392
rect 45064 17358 45120 17392
rect 45154 17358 45284 17392
rect 43996 17323 45284 17358
rect 43996 17308 44097 17323
rect 43996 17274 44029 17308
rect 44063 17274 44097 17308
rect 43996 17218 44097 17274
rect 45183 17308 45284 17323
rect 45183 17274 45216 17308
rect 45250 17274 45284 17308
rect 43996 17184 44029 17218
rect 44063 17184 44097 17218
rect 43996 17128 44097 17184
rect 43996 17094 44029 17128
rect 44063 17094 44097 17128
rect 43996 17038 44097 17094
rect 43996 17004 44029 17038
rect 44063 17004 44097 17038
rect 43996 16948 44097 17004
rect 43996 16914 44029 16948
rect 44063 16914 44097 16948
rect 43996 16858 44097 16914
rect 43996 16824 44029 16858
rect 44063 16824 44097 16858
rect 43996 16768 44097 16824
rect 43996 16734 44029 16768
rect 44063 16734 44097 16768
rect 43996 16678 44097 16734
rect 43996 16644 44029 16678
rect 44063 16644 44097 16678
rect 43996 16588 44097 16644
rect 43996 16554 44029 16588
rect 44063 16554 44097 16588
rect 43996 16498 44097 16554
rect 43996 16464 44029 16498
rect 44063 16464 44097 16498
rect 43996 16408 44097 16464
rect 43996 16374 44029 16408
rect 44063 16374 44097 16408
rect 43996 16318 44097 16374
rect 43996 16284 44029 16318
rect 44063 16284 44097 16318
rect 45183 17218 45284 17274
rect 45183 17184 45216 17218
rect 45250 17184 45284 17218
rect 45183 17128 45284 17184
rect 45183 17094 45216 17128
rect 45250 17094 45284 17128
rect 45183 17038 45284 17094
rect 45183 17004 45216 17038
rect 45250 17004 45284 17038
rect 45183 16948 45284 17004
rect 45183 16914 45216 16948
rect 45250 16914 45284 16948
rect 45183 16858 45284 16914
rect 45183 16824 45216 16858
rect 45250 16824 45284 16858
rect 45183 16768 45284 16824
rect 45183 16734 45216 16768
rect 45250 16734 45284 16768
rect 45183 16678 45284 16734
rect 45183 16644 45216 16678
rect 45250 16644 45284 16678
rect 45183 16588 45284 16644
rect 45183 16554 45216 16588
rect 45250 16554 45284 16588
rect 45183 16498 45284 16554
rect 45183 16464 45216 16498
rect 45250 16464 45284 16498
rect 45183 16408 45284 16464
rect 45183 16374 45216 16408
rect 45250 16374 45284 16408
rect 45183 16318 45284 16374
rect 43996 16237 44097 16284
rect 45183 16284 45216 16318
rect 45250 16284 45284 16318
rect 45183 16237 45284 16284
rect 43996 16228 45284 16237
rect 43996 16194 44029 16228
rect 44063 16205 45216 16228
rect 44063 16194 44130 16205
rect 43996 16171 44130 16194
rect 44164 16171 44220 16205
rect 44254 16171 44310 16205
rect 44344 16171 44400 16205
rect 44434 16171 44490 16205
rect 44524 16171 44580 16205
rect 44614 16171 44670 16205
rect 44704 16171 44760 16205
rect 44794 16171 44850 16205
rect 44884 16171 44940 16205
rect 44974 16171 45030 16205
rect 45064 16171 45120 16205
rect 45154 16194 45216 16205
rect 45250 16194 45284 16228
rect 45154 16171 45284 16194
rect 43996 16136 45284 16171
rect 41276 16032 42564 16064
rect 41276 15998 41410 16032
rect 41444 15998 41500 16032
rect 41534 15998 41590 16032
rect 41624 15998 41680 16032
rect 41714 15998 41770 16032
rect 41804 15998 41860 16032
rect 41894 15998 41950 16032
rect 41984 15998 42040 16032
rect 42074 15998 42130 16032
rect 42164 15998 42220 16032
rect 42254 15998 42310 16032
rect 42344 15998 42400 16032
rect 42434 15998 42564 16032
rect 41276 15963 42564 15998
rect 41276 15948 41377 15963
rect 41276 15914 41309 15948
rect 41343 15914 41377 15948
rect 41276 15858 41377 15914
rect 42463 15948 42564 15963
rect 42463 15914 42496 15948
rect 42530 15914 42564 15948
rect 41276 15824 41309 15858
rect 41343 15824 41377 15858
rect 41276 15768 41377 15824
rect 41276 15734 41309 15768
rect 41343 15734 41377 15768
rect 41276 15678 41377 15734
rect 41276 15644 41309 15678
rect 41343 15644 41377 15678
rect 41276 15588 41377 15644
rect 41276 15554 41309 15588
rect 41343 15554 41377 15588
rect 41276 15498 41377 15554
rect 41276 15464 41309 15498
rect 41343 15464 41377 15498
rect 41276 15408 41377 15464
rect 41276 15374 41309 15408
rect 41343 15374 41377 15408
rect 41276 15318 41377 15374
rect 41276 15284 41309 15318
rect 41343 15284 41377 15318
rect 41276 15228 41377 15284
rect 41276 15194 41309 15228
rect 41343 15194 41377 15228
rect 41276 15138 41377 15194
rect 41276 15104 41309 15138
rect 41343 15104 41377 15138
rect 41276 15048 41377 15104
rect 41276 15014 41309 15048
rect 41343 15014 41377 15048
rect 41276 14958 41377 15014
rect 41276 14924 41309 14958
rect 41343 14924 41377 14958
rect 42463 15858 42564 15914
rect 42463 15824 42496 15858
rect 42530 15824 42564 15858
rect 42463 15768 42564 15824
rect 42463 15734 42496 15768
rect 42530 15734 42564 15768
rect 42463 15678 42564 15734
rect 42463 15644 42496 15678
rect 42530 15644 42564 15678
rect 42463 15588 42564 15644
rect 42463 15554 42496 15588
rect 42530 15554 42564 15588
rect 42463 15498 42564 15554
rect 42463 15464 42496 15498
rect 42530 15464 42564 15498
rect 42463 15408 42564 15464
rect 42463 15374 42496 15408
rect 42530 15374 42564 15408
rect 42463 15318 42564 15374
rect 42463 15284 42496 15318
rect 42530 15284 42564 15318
rect 42463 15228 42564 15284
rect 42463 15194 42496 15228
rect 42530 15194 42564 15228
rect 42463 15138 42564 15194
rect 42463 15104 42496 15138
rect 42530 15104 42564 15138
rect 42463 15048 42564 15104
rect 42463 15014 42496 15048
rect 42530 15014 42564 15048
rect 42463 14958 42564 15014
rect 41276 14877 41377 14924
rect 42463 14924 42496 14958
rect 42530 14924 42564 14958
rect 42463 14877 42564 14924
rect 41276 14868 42564 14877
rect 41276 14834 41309 14868
rect 41343 14845 42496 14868
rect 41343 14834 41410 14845
rect 41276 14811 41410 14834
rect 41444 14811 41500 14845
rect 41534 14811 41590 14845
rect 41624 14811 41680 14845
rect 41714 14811 41770 14845
rect 41804 14811 41860 14845
rect 41894 14811 41950 14845
rect 41984 14811 42040 14845
rect 42074 14811 42130 14845
rect 42164 14811 42220 14845
rect 42254 14811 42310 14845
rect 42344 14811 42400 14845
rect 42434 14834 42496 14845
rect 42530 14834 42564 14868
rect 42434 14811 42564 14834
rect 41276 14776 42564 14811
rect 42636 16032 43924 16064
rect 42636 15998 42770 16032
rect 42804 15998 42860 16032
rect 42894 15998 42950 16032
rect 42984 15998 43040 16032
rect 43074 15998 43130 16032
rect 43164 15998 43220 16032
rect 43254 15998 43310 16032
rect 43344 15998 43400 16032
rect 43434 15998 43490 16032
rect 43524 15998 43580 16032
rect 43614 15998 43670 16032
rect 43704 15998 43760 16032
rect 43794 15998 43924 16032
rect 42636 15963 43924 15998
rect 42636 15948 42737 15963
rect 42636 15914 42669 15948
rect 42703 15914 42737 15948
rect 42636 15858 42737 15914
rect 43823 15948 43924 15963
rect 43823 15914 43856 15948
rect 43890 15914 43924 15948
rect 42636 15824 42669 15858
rect 42703 15824 42737 15858
rect 42636 15768 42737 15824
rect 42636 15734 42669 15768
rect 42703 15734 42737 15768
rect 42636 15678 42737 15734
rect 42636 15644 42669 15678
rect 42703 15644 42737 15678
rect 42636 15588 42737 15644
rect 42636 15554 42669 15588
rect 42703 15554 42737 15588
rect 42636 15498 42737 15554
rect 42636 15464 42669 15498
rect 42703 15464 42737 15498
rect 42636 15408 42737 15464
rect 42636 15374 42669 15408
rect 42703 15374 42737 15408
rect 42636 15318 42737 15374
rect 42636 15284 42669 15318
rect 42703 15284 42737 15318
rect 42636 15228 42737 15284
rect 42636 15194 42669 15228
rect 42703 15194 42737 15228
rect 42636 15138 42737 15194
rect 42636 15104 42669 15138
rect 42703 15104 42737 15138
rect 42636 15048 42737 15104
rect 42636 15014 42669 15048
rect 42703 15014 42737 15048
rect 42636 14958 42737 15014
rect 42636 14924 42669 14958
rect 42703 14924 42737 14958
rect 43823 15858 43924 15914
rect 43823 15824 43856 15858
rect 43890 15824 43924 15858
rect 43823 15768 43924 15824
rect 43823 15734 43856 15768
rect 43890 15734 43924 15768
rect 43823 15678 43924 15734
rect 43823 15644 43856 15678
rect 43890 15644 43924 15678
rect 43823 15588 43924 15644
rect 43823 15554 43856 15588
rect 43890 15554 43924 15588
rect 43823 15498 43924 15554
rect 43823 15464 43856 15498
rect 43890 15464 43924 15498
rect 43823 15408 43924 15464
rect 43823 15374 43856 15408
rect 43890 15374 43924 15408
rect 43823 15318 43924 15374
rect 43823 15284 43856 15318
rect 43890 15284 43924 15318
rect 43823 15228 43924 15284
rect 43823 15194 43856 15228
rect 43890 15194 43924 15228
rect 43823 15138 43924 15194
rect 43823 15104 43856 15138
rect 43890 15104 43924 15138
rect 43823 15048 43924 15104
rect 43823 15014 43856 15048
rect 43890 15014 43924 15048
rect 43823 14958 43924 15014
rect 42636 14877 42737 14924
rect 43823 14924 43856 14958
rect 43890 14924 43924 14958
rect 43823 14877 43924 14924
rect 42636 14868 43924 14877
rect 42636 14834 42669 14868
rect 42703 14845 43856 14868
rect 42703 14834 42770 14845
rect 42636 14811 42770 14834
rect 42804 14811 42860 14845
rect 42894 14811 42950 14845
rect 42984 14811 43040 14845
rect 43074 14811 43130 14845
rect 43164 14811 43220 14845
rect 43254 14811 43310 14845
rect 43344 14811 43400 14845
rect 43434 14811 43490 14845
rect 43524 14811 43580 14845
rect 43614 14811 43670 14845
rect 43704 14811 43760 14845
rect 43794 14834 43856 14845
rect 43890 14834 43924 14868
rect 43794 14811 43924 14834
rect 42636 14776 43924 14811
rect 43996 16032 45284 16064
rect 43996 15998 44130 16032
rect 44164 15998 44220 16032
rect 44254 15998 44310 16032
rect 44344 15998 44400 16032
rect 44434 15998 44490 16032
rect 44524 15998 44580 16032
rect 44614 15998 44670 16032
rect 44704 15998 44760 16032
rect 44794 15998 44850 16032
rect 44884 15998 44940 16032
rect 44974 15998 45030 16032
rect 45064 15998 45120 16032
rect 45154 15998 45284 16032
rect 43996 15963 45284 15998
rect 43996 15948 44097 15963
rect 43996 15914 44029 15948
rect 44063 15914 44097 15948
rect 43996 15858 44097 15914
rect 45183 15948 45284 15963
rect 45183 15914 45216 15948
rect 45250 15914 45284 15948
rect 43996 15824 44029 15858
rect 44063 15824 44097 15858
rect 43996 15768 44097 15824
rect 43996 15734 44029 15768
rect 44063 15734 44097 15768
rect 43996 15678 44097 15734
rect 43996 15644 44029 15678
rect 44063 15644 44097 15678
rect 43996 15588 44097 15644
rect 43996 15554 44029 15588
rect 44063 15554 44097 15588
rect 43996 15498 44097 15554
rect 43996 15464 44029 15498
rect 44063 15464 44097 15498
rect 43996 15408 44097 15464
rect 43996 15374 44029 15408
rect 44063 15374 44097 15408
rect 43996 15318 44097 15374
rect 43996 15284 44029 15318
rect 44063 15284 44097 15318
rect 43996 15228 44097 15284
rect 43996 15194 44029 15228
rect 44063 15194 44097 15228
rect 43996 15138 44097 15194
rect 43996 15104 44029 15138
rect 44063 15104 44097 15138
rect 43996 15048 44097 15104
rect 43996 15014 44029 15048
rect 44063 15014 44097 15048
rect 43996 14958 44097 15014
rect 43996 14924 44029 14958
rect 44063 14924 44097 14958
rect 45183 15858 45284 15914
rect 45183 15824 45216 15858
rect 45250 15824 45284 15858
rect 45183 15768 45284 15824
rect 45183 15734 45216 15768
rect 45250 15734 45284 15768
rect 45183 15678 45284 15734
rect 45183 15644 45216 15678
rect 45250 15644 45284 15678
rect 45183 15588 45284 15644
rect 45183 15554 45216 15588
rect 45250 15554 45284 15588
rect 45183 15498 45284 15554
rect 45183 15464 45216 15498
rect 45250 15464 45284 15498
rect 45183 15408 45284 15464
rect 45183 15374 45216 15408
rect 45250 15374 45284 15408
rect 45183 15318 45284 15374
rect 45183 15284 45216 15318
rect 45250 15284 45284 15318
rect 45183 15228 45284 15284
rect 45183 15194 45216 15228
rect 45250 15194 45284 15228
rect 45183 15138 45284 15194
rect 45183 15104 45216 15138
rect 45250 15104 45284 15138
rect 45183 15048 45284 15104
rect 45183 15014 45216 15048
rect 45250 15014 45284 15048
rect 45183 14958 45284 15014
rect 43996 14877 44097 14924
rect 45183 14924 45216 14958
rect 45250 14924 45284 14958
rect 45183 14877 45284 14924
rect 43996 14868 45284 14877
rect 43996 14834 44029 14868
rect 44063 14845 45216 14868
rect 44063 14834 44130 14845
rect 43996 14811 44130 14834
rect 44164 14811 44220 14845
rect 44254 14811 44310 14845
rect 44344 14811 44400 14845
rect 44434 14811 44490 14845
rect 44524 14811 44580 14845
rect 44614 14811 44670 14845
rect 44704 14811 44760 14845
rect 44794 14811 44850 14845
rect 44884 14811 44940 14845
rect 44974 14811 45030 14845
rect 45064 14811 45120 14845
rect 45154 14834 45216 14845
rect 45250 14834 45284 14868
rect 45154 14811 45284 14834
rect 43996 14776 45284 14811
rect 45400 13850 45480 13880
rect 45400 13810 45420 13850
rect 45460 13810 45480 13850
rect 45400 13750 45480 13810
rect 45400 13710 45420 13750
rect 45460 13710 45480 13750
rect 45400 13680 45480 13710
rect 41900 13240 41980 13270
rect 41900 13200 41920 13240
rect 41960 13200 41980 13240
rect 41900 13140 41980 13200
rect 41900 13100 41920 13140
rect 41960 13100 41980 13140
rect 41900 13040 41980 13100
rect 41900 13000 41920 13040
rect 41960 13000 41980 13040
rect 41900 12940 41980 13000
rect 41900 12900 41920 12940
rect 41960 12900 41980 12940
rect 41900 12840 41980 12900
rect 41900 12800 41920 12840
rect 41960 12800 41980 12840
rect 41900 12770 41980 12800
rect 44580 13240 44660 13270
rect 44580 13200 44600 13240
rect 44640 13200 44660 13240
rect 44580 13140 44660 13200
rect 44580 13100 44600 13140
rect 44640 13100 44660 13140
rect 44580 13040 44660 13100
rect 44580 13000 44600 13040
rect 44640 13000 44660 13040
rect 44580 12940 44660 13000
rect 44580 12900 44600 12940
rect 44640 12900 44660 12940
rect 44580 12840 44660 12900
rect 44580 12800 44600 12840
rect 44640 12800 44660 12840
rect 44580 12770 44660 12800
rect 42800 12320 42880 12350
rect 42800 12280 42820 12320
rect 42860 12280 42880 12320
rect 42800 12240 42880 12280
rect 42800 12200 42820 12240
rect 42860 12200 42880 12240
rect 42800 12160 42880 12200
rect 42800 12120 42820 12160
rect 42860 12120 42880 12160
rect 42800 12090 42880 12120
rect 43680 12320 43760 12350
rect 43680 12280 43700 12320
rect 43740 12280 43760 12320
rect 43680 12240 43760 12280
rect 43680 12200 43700 12240
rect 43740 12200 43760 12240
rect 43680 12160 43760 12200
rect 43680 12120 43700 12160
rect 43740 12120 43760 12160
rect 43680 12090 43760 12120
<< nsubdiff >>
rect 38603 18555 38699 18589
rect 38959 18555 39055 18589
rect 38603 18493 38637 18555
rect 39021 18493 39055 18555
rect 38603 16527 38637 16589
rect 39021 16527 39055 16589
rect 38603 16493 38699 16527
rect 38959 16493 39055 16527
rect 39383 18561 39479 18595
rect 39739 18561 39835 18595
rect 39383 18499 39417 18561
rect 39801 18499 39835 18561
rect 39383 14957 39417 15019
rect 40163 18563 40259 18597
rect 40851 18563 40947 18597
rect 40163 18501 40197 18563
rect 40913 18501 40947 18563
rect 40163 16181 40197 16243
rect 41439 18602 42401 18621
rect 41439 18568 41550 18602
rect 41584 18568 41640 18602
rect 41674 18568 41730 18602
rect 41764 18568 41820 18602
rect 41854 18568 41910 18602
rect 41944 18568 42000 18602
rect 42034 18568 42090 18602
rect 42124 18568 42180 18602
rect 42214 18568 42270 18602
rect 42304 18568 42401 18602
rect 41439 18549 42401 18568
rect 41439 18508 41511 18549
rect 41439 18474 41458 18508
rect 41492 18474 41511 18508
rect 42329 18489 42401 18549
rect 41439 18418 41511 18474
rect 41439 18384 41458 18418
rect 41492 18384 41511 18418
rect 41439 18328 41511 18384
rect 41439 18294 41458 18328
rect 41492 18294 41511 18328
rect 41439 18238 41511 18294
rect 41439 18204 41458 18238
rect 41492 18204 41511 18238
rect 41439 18148 41511 18204
rect 41439 18114 41458 18148
rect 41492 18114 41511 18148
rect 41439 18058 41511 18114
rect 41439 18024 41458 18058
rect 41492 18024 41511 18058
rect 41439 17968 41511 18024
rect 41439 17934 41458 17968
rect 41492 17934 41511 17968
rect 41439 17878 41511 17934
rect 41439 17844 41458 17878
rect 41492 17844 41511 17878
rect 41439 17788 41511 17844
rect 42329 18455 42348 18489
rect 42382 18455 42401 18489
rect 42329 18399 42401 18455
rect 42329 18365 42348 18399
rect 42382 18365 42401 18399
rect 42329 18309 42401 18365
rect 42329 18275 42348 18309
rect 42382 18275 42401 18309
rect 42329 18219 42401 18275
rect 42329 18185 42348 18219
rect 42382 18185 42401 18219
rect 42329 18129 42401 18185
rect 42329 18095 42348 18129
rect 42382 18095 42401 18129
rect 42329 18039 42401 18095
rect 42329 18005 42348 18039
rect 42382 18005 42401 18039
rect 42329 17949 42401 18005
rect 42329 17915 42348 17949
rect 42382 17915 42401 17949
rect 42329 17859 42401 17915
rect 42329 17825 42348 17859
rect 42382 17825 42401 17859
rect 41439 17754 41458 17788
rect 41492 17754 41511 17788
rect 41439 17731 41511 17754
rect 42329 17769 42401 17825
rect 42329 17735 42348 17769
rect 42382 17735 42401 17769
rect 42329 17731 42401 17735
rect 41439 17712 42401 17731
rect 41439 17678 41516 17712
rect 41550 17678 41606 17712
rect 41640 17678 41696 17712
rect 41730 17678 41786 17712
rect 41820 17678 41876 17712
rect 41910 17678 41966 17712
rect 42000 17678 42056 17712
rect 42090 17678 42146 17712
rect 42180 17678 42236 17712
rect 42270 17678 42401 17712
rect 41439 17659 42401 17678
rect 42799 18602 43761 18621
rect 42799 18568 42910 18602
rect 42944 18568 43000 18602
rect 43034 18568 43090 18602
rect 43124 18568 43180 18602
rect 43214 18568 43270 18602
rect 43304 18568 43360 18602
rect 43394 18568 43450 18602
rect 43484 18568 43540 18602
rect 43574 18568 43630 18602
rect 43664 18568 43761 18602
rect 42799 18549 43761 18568
rect 42799 18508 42871 18549
rect 42799 18474 42818 18508
rect 42852 18474 42871 18508
rect 43689 18489 43761 18549
rect 42799 18418 42871 18474
rect 42799 18384 42818 18418
rect 42852 18384 42871 18418
rect 42799 18328 42871 18384
rect 42799 18294 42818 18328
rect 42852 18294 42871 18328
rect 42799 18238 42871 18294
rect 42799 18204 42818 18238
rect 42852 18204 42871 18238
rect 42799 18148 42871 18204
rect 42799 18114 42818 18148
rect 42852 18114 42871 18148
rect 42799 18058 42871 18114
rect 42799 18024 42818 18058
rect 42852 18024 42871 18058
rect 42799 17968 42871 18024
rect 42799 17934 42818 17968
rect 42852 17934 42871 17968
rect 42799 17878 42871 17934
rect 42799 17844 42818 17878
rect 42852 17844 42871 17878
rect 42799 17788 42871 17844
rect 43689 18455 43708 18489
rect 43742 18455 43761 18489
rect 43689 18399 43761 18455
rect 43689 18365 43708 18399
rect 43742 18365 43761 18399
rect 43689 18309 43761 18365
rect 43689 18275 43708 18309
rect 43742 18275 43761 18309
rect 43689 18219 43761 18275
rect 43689 18185 43708 18219
rect 43742 18185 43761 18219
rect 43689 18129 43761 18185
rect 43689 18095 43708 18129
rect 43742 18095 43761 18129
rect 43689 18039 43761 18095
rect 43689 18005 43708 18039
rect 43742 18005 43761 18039
rect 43689 17949 43761 18005
rect 43689 17915 43708 17949
rect 43742 17915 43761 17949
rect 43689 17859 43761 17915
rect 43689 17825 43708 17859
rect 43742 17825 43761 17859
rect 42799 17754 42818 17788
rect 42852 17754 42871 17788
rect 42799 17731 42871 17754
rect 43689 17769 43761 17825
rect 43689 17735 43708 17769
rect 43742 17735 43761 17769
rect 43689 17731 43761 17735
rect 42799 17712 43761 17731
rect 42799 17678 42876 17712
rect 42910 17678 42966 17712
rect 43000 17678 43056 17712
rect 43090 17678 43146 17712
rect 43180 17678 43236 17712
rect 43270 17678 43326 17712
rect 43360 17678 43416 17712
rect 43450 17678 43506 17712
rect 43540 17678 43596 17712
rect 43630 17678 43761 17712
rect 42799 17659 43761 17678
rect 44159 18602 45121 18621
rect 44159 18568 44270 18602
rect 44304 18568 44360 18602
rect 44394 18568 44450 18602
rect 44484 18568 44540 18602
rect 44574 18568 44630 18602
rect 44664 18568 44720 18602
rect 44754 18568 44810 18602
rect 44844 18568 44900 18602
rect 44934 18568 44990 18602
rect 45024 18568 45121 18602
rect 44159 18549 45121 18568
rect 44159 18508 44231 18549
rect 44159 18474 44178 18508
rect 44212 18474 44231 18508
rect 45049 18489 45121 18549
rect 44159 18418 44231 18474
rect 44159 18384 44178 18418
rect 44212 18384 44231 18418
rect 44159 18328 44231 18384
rect 44159 18294 44178 18328
rect 44212 18294 44231 18328
rect 44159 18238 44231 18294
rect 44159 18204 44178 18238
rect 44212 18204 44231 18238
rect 44159 18148 44231 18204
rect 44159 18114 44178 18148
rect 44212 18114 44231 18148
rect 44159 18058 44231 18114
rect 44159 18024 44178 18058
rect 44212 18024 44231 18058
rect 44159 17968 44231 18024
rect 44159 17934 44178 17968
rect 44212 17934 44231 17968
rect 44159 17878 44231 17934
rect 44159 17844 44178 17878
rect 44212 17844 44231 17878
rect 44159 17788 44231 17844
rect 45049 18455 45068 18489
rect 45102 18455 45121 18489
rect 45049 18399 45121 18455
rect 45049 18365 45068 18399
rect 45102 18365 45121 18399
rect 45049 18309 45121 18365
rect 45049 18275 45068 18309
rect 45102 18275 45121 18309
rect 45049 18219 45121 18275
rect 45049 18185 45068 18219
rect 45102 18185 45121 18219
rect 45049 18129 45121 18185
rect 45049 18095 45068 18129
rect 45102 18095 45121 18129
rect 45049 18039 45121 18095
rect 45049 18005 45068 18039
rect 45102 18005 45121 18039
rect 45049 17949 45121 18005
rect 45049 17915 45068 17949
rect 45102 17915 45121 17949
rect 45049 17859 45121 17915
rect 45049 17825 45068 17859
rect 45102 17825 45121 17859
rect 44159 17754 44178 17788
rect 44212 17754 44231 17788
rect 44159 17731 44231 17754
rect 45049 17769 45121 17825
rect 45049 17735 45068 17769
rect 45102 17735 45121 17769
rect 45049 17731 45121 17735
rect 44159 17712 45121 17731
rect 44159 17678 44236 17712
rect 44270 17678 44326 17712
rect 44360 17678 44416 17712
rect 44450 17678 44506 17712
rect 44540 17678 44596 17712
rect 44630 17678 44686 17712
rect 44720 17678 44776 17712
rect 44810 17678 44866 17712
rect 44900 17678 44956 17712
rect 44990 17678 45121 17712
rect 44159 17659 45121 17678
rect 45483 18563 45579 18597
rect 46171 18563 46267 18597
rect 45483 18501 45517 18563
rect 40913 16181 40947 16243
rect 40163 16147 40259 16181
rect 40851 16147 40947 16181
rect 41439 17242 42401 17261
rect 41439 17208 41550 17242
rect 41584 17208 41640 17242
rect 41674 17208 41730 17242
rect 41764 17208 41820 17242
rect 41854 17208 41910 17242
rect 41944 17208 42000 17242
rect 42034 17208 42090 17242
rect 42124 17208 42180 17242
rect 42214 17208 42270 17242
rect 42304 17208 42401 17242
rect 41439 17189 42401 17208
rect 41439 17148 41511 17189
rect 41439 17114 41458 17148
rect 41492 17114 41511 17148
rect 42329 17129 42401 17189
rect 41439 17058 41511 17114
rect 41439 17024 41458 17058
rect 41492 17024 41511 17058
rect 41439 16968 41511 17024
rect 41439 16934 41458 16968
rect 41492 16934 41511 16968
rect 41439 16878 41511 16934
rect 41439 16844 41458 16878
rect 41492 16844 41511 16878
rect 41439 16788 41511 16844
rect 41439 16754 41458 16788
rect 41492 16754 41511 16788
rect 41439 16698 41511 16754
rect 41439 16664 41458 16698
rect 41492 16664 41511 16698
rect 41439 16608 41511 16664
rect 41439 16574 41458 16608
rect 41492 16574 41511 16608
rect 41439 16518 41511 16574
rect 41439 16484 41458 16518
rect 41492 16484 41511 16518
rect 41439 16428 41511 16484
rect 42329 17095 42348 17129
rect 42382 17095 42401 17129
rect 42329 17039 42401 17095
rect 42329 17005 42348 17039
rect 42382 17005 42401 17039
rect 42329 16949 42401 17005
rect 42329 16915 42348 16949
rect 42382 16915 42401 16949
rect 42329 16859 42401 16915
rect 42329 16825 42348 16859
rect 42382 16825 42401 16859
rect 42329 16769 42401 16825
rect 42329 16735 42348 16769
rect 42382 16735 42401 16769
rect 42329 16679 42401 16735
rect 42329 16645 42348 16679
rect 42382 16645 42401 16679
rect 42329 16589 42401 16645
rect 42329 16555 42348 16589
rect 42382 16555 42401 16589
rect 42329 16499 42401 16555
rect 42329 16465 42348 16499
rect 42382 16465 42401 16499
rect 41439 16394 41458 16428
rect 41492 16394 41511 16428
rect 41439 16371 41511 16394
rect 42329 16409 42401 16465
rect 42329 16375 42348 16409
rect 42382 16375 42401 16409
rect 42329 16371 42401 16375
rect 41439 16352 42401 16371
rect 41439 16318 41516 16352
rect 41550 16318 41606 16352
rect 41640 16318 41696 16352
rect 41730 16318 41786 16352
rect 41820 16318 41876 16352
rect 41910 16318 41966 16352
rect 42000 16318 42056 16352
rect 42090 16318 42146 16352
rect 42180 16318 42236 16352
rect 42270 16318 42401 16352
rect 41439 16299 42401 16318
rect 42799 17242 43761 17261
rect 42799 17208 42910 17242
rect 42944 17208 43000 17242
rect 43034 17208 43090 17242
rect 43124 17208 43180 17242
rect 43214 17208 43270 17242
rect 43304 17208 43360 17242
rect 43394 17208 43450 17242
rect 43484 17208 43540 17242
rect 43574 17208 43630 17242
rect 43664 17208 43761 17242
rect 42799 17189 43761 17208
rect 42799 17148 42871 17189
rect 42799 17114 42818 17148
rect 42852 17114 42871 17148
rect 43689 17129 43761 17189
rect 42799 17058 42871 17114
rect 42799 17024 42818 17058
rect 42852 17024 42871 17058
rect 42799 16968 42871 17024
rect 42799 16934 42818 16968
rect 42852 16934 42871 16968
rect 42799 16878 42871 16934
rect 42799 16844 42818 16878
rect 42852 16844 42871 16878
rect 42799 16788 42871 16844
rect 42799 16754 42818 16788
rect 42852 16754 42871 16788
rect 42799 16698 42871 16754
rect 42799 16664 42818 16698
rect 42852 16664 42871 16698
rect 42799 16608 42871 16664
rect 42799 16574 42818 16608
rect 42852 16574 42871 16608
rect 42799 16518 42871 16574
rect 42799 16484 42818 16518
rect 42852 16484 42871 16518
rect 42799 16428 42871 16484
rect 43689 17095 43708 17129
rect 43742 17095 43761 17129
rect 43689 17039 43761 17095
rect 43689 17005 43708 17039
rect 43742 17005 43761 17039
rect 43689 16949 43761 17005
rect 43689 16915 43708 16949
rect 43742 16915 43761 16949
rect 43689 16859 43761 16915
rect 43689 16825 43708 16859
rect 43742 16825 43761 16859
rect 43689 16769 43761 16825
rect 43689 16735 43708 16769
rect 43742 16735 43761 16769
rect 43689 16679 43761 16735
rect 43689 16645 43708 16679
rect 43742 16645 43761 16679
rect 43689 16589 43761 16645
rect 43689 16555 43708 16589
rect 43742 16555 43761 16589
rect 43689 16499 43761 16555
rect 43689 16465 43708 16499
rect 43742 16465 43761 16499
rect 42799 16394 42818 16428
rect 42852 16394 42871 16428
rect 42799 16371 42871 16394
rect 43689 16409 43761 16465
rect 43689 16375 43708 16409
rect 43742 16375 43761 16409
rect 43689 16371 43761 16375
rect 42799 16352 43761 16371
rect 42799 16318 42876 16352
rect 42910 16318 42966 16352
rect 43000 16318 43056 16352
rect 43090 16318 43146 16352
rect 43180 16318 43236 16352
rect 43270 16318 43326 16352
rect 43360 16318 43416 16352
rect 43450 16318 43506 16352
rect 43540 16318 43596 16352
rect 43630 16318 43761 16352
rect 42799 16299 43761 16318
rect 44159 17242 45121 17261
rect 44159 17208 44270 17242
rect 44304 17208 44360 17242
rect 44394 17208 44450 17242
rect 44484 17208 44540 17242
rect 44574 17208 44630 17242
rect 44664 17208 44720 17242
rect 44754 17208 44810 17242
rect 44844 17208 44900 17242
rect 44934 17208 44990 17242
rect 45024 17208 45121 17242
rect 44159 17189 45121 17208
rect 44159 17148 44231 17189
rect 44159 17114 44178 17148
rect 44212 17114 44231 17148
rect 45049 17129 45121 17189
rect 44159 17058 44231 17114
rect 44159 17024 44178 17058
rect 44212 17024 44231 17058
rect 44159 16968 44231 17024
rect 44159 16934 44178 16968
rect 44212 16934 44231 16968
rect 44159 16878 44231 16934
rect 44159 16844 44178 16878
rect 44212 16844 44231 16878
rect 44159 16788 44231 16844
rect 44159 16754 44178 16788
rect 44212 16754 44231 16788
rect 44159 16698 44231 16754
rect 44159 16664 44178 16698
rect 44212 16664 44231 16698
rect 44159 16608 44231 16664
rect 44159 16574 44178 16608
rect 44212 16574 44231 16608
rect 44159 16518 44231 16574
rect 44159 16484 44178 16518
rect 44212 16484 44231 16518
rect 44159 16428 44231 16484
rect 45049 17095 45068 17129
rect 45102 17095 45121 17129
rect 45049 17039 45121 17095
rect 45049 17005 45068 17039
rect 45102 17005 45121 17039
rect 45049 16949 45121 17005
rect 45049 16915 45068 16949
rect 45102 16915 45121 16949
rect 45049 16859 45121 16915
rect 45049 16825 45068 16859
rect 45102 16825 45121 16859
rect 45049 16769 45121 16825
rect 45049 16735 45068 16769
rect 45102 16735 45121 16769
rect 45049 16679 45121 16735
rect 45049 16645 45068 16679
rect 45102 16645 45121 16679
rect 45049 16589 45121 16645
rect 45049 16555 45068 16589
rect 45102 16555 45121 16589
rect 45049 16499 45121 16555
rect 45049 16465 45068 16499
rect 45102 16465 45121 16499
rect 44159 16394 44178 16428
rect 44212 16394 44231 16428
rect 44159 16371 44231 16394
rect 45049 16409 45121 16465
rect 45049 16375 45068 16409
rect 45102 16375 45121 16409
rect 45049 16371 45121 16375
rect 44159 16352 45121 16371
rect 44159 16318 44236 16352
rect 44270 16318 44326 16352
rect 44360 16318 44416 16352
rect 44450 16318 44506 16352
rect 44540 16318 44596 16352
rect 44630 16318 44686 16352
rect 44720 16318 44776 16352
rect 44810 16318 44866 16352
rect 44900 16318 44956 16352
rect 44990 16318 45121 16352
rect 44159 16299 45121 16318
rect 46233 18501 46267 18563
rect 45483 16181 45517 16243
rect 46233 16181 46267 16243
rect 45483 16147 45579 16181
rect 46171 16147 46267 16181
rect 46593 18561 46689 18595
rect 46949 18561 47045 18595
rect 46593 18499 46627 18561
rect 39801 14957 39835 15019
rect 39383 14923 39479 14957
rect 39739 14923 39835 14957
rect 41439 15882 42401 15901
rect 41439 15848 41550 15882
rect 41584 15848 41640 15882
rect 41674 15848 41730 15882
rect 41764 15848 41820 15882
rect 41854 15848 41910 15882
rect 41944 15848 42000 15882
rect 42034 15848 42090 15882
rect 42124 15848 42180 15882
rect 42214 15848 42270 15882
rect 42304 15848 42401 15882
rect 41439 15829 42401 15848
rect 41439 15788 41511 15829
rect 41439 15754 41458 15788
rect 41492 15754 41511 15788
rect 42329 15769 42401 15829
rect 41439 15698 41511 15754
rect 41439 15664 41458 15698
rect 41492 15664 41511 15698
rect 41439 15608 41511 15664
rect 41439 15574 41458 15608
rect 41492 15574 41511 15608
rect 41439 15518 41511 15574
rect 41439 15484 41458 15518
rect 41492 15484 41511 15518
rect 41439 15428 41511 15484
rect 41439 15394 41458 15428
rect 41492 15394 41511 15428
rect 41439 15338 41511 15394
rect 41439 15304 41458 15338
rect 41492 15304 41511 15338
rect 41439 15248 41511 15304
rect 41439 15214 41458 15248
rect 41492 15214 41511 15248
rect 41439 15158 41511 15214
rect 41439 15124 41458 15158
rect 41492 15124 41511 15158
rect 41439 15068 41511 15124
rect 42329 15735 42348 15769
rect 42382 15735 42401 15769
rect 42329 15679 42401 15735
rect 42329 15645 42348 15679
rect 42382 15645 42401 15679
rect 42329 15589 42401 15645
rect 42329 15555 42348 15589
rect 42382 15555 42401 15589
rect 42329 15499 42401 15555
rect 42329 15465 42348 15499
rect 42382 15465 42401 15499
rect 42329 15409 42401 15465
rect 42329 15375 42348 15409
rect 42382 15375 42401 15409
rect 42329 15319 42401 15375
rect 42329 15285 42348 15319
rect 42382 15285 42401 15319
rect 42329 15229 42401 15285
rect 42329 15195 42348 15229
rect 42382 15195 42401 15229
rect 42329 15139 42401 15195
rect 42329 15105 42348 15139
rect 42382 15105 42401 15139
rect 41439 15034 41458 15068
rect 41492 15034 41511 15068
rect 41439 15011 41511 15034
rect 42329 15049 42401 15105
rect 42329 15015 42348 15049
rect 42382 15015 42401 15049
rect 42329 15011 42401 15015
rect 41439 14992 42401 15011
rect 41439 14958 41516 14992
rect 41550 14958 41606 14992
rect 41640 14958 41696 14992
rect 41730 14958 41786 14992
rect 41820 14958 41876 14992
rect 41910 14958 41966 14992
rect 42000 14958 42056 14992
rect 42090 14958 42146 14992
rect 42180 14958 42236 14992
rect 42270 14958 42401 14992
rect 41439 14939 42401 14958
rect 42799 15882 43761 15901
rect 42799 15848 42910 15882
rect 42944 15848 43000 15882
rect 43034 15848 43090 15882
rect 43124 15848 43180 15882
rect 43214 15848 43270 15882
rect 43304 15848 43360 15882
rect 43394 15848 43450 15882
rect 43484 15848 43540 15882
rect 43574 15848 43630 15882
rect 43664 15848 43761 15882
rect 42799 15829 43761 15848
rect 42799 15788 42871 15829
rect 42799 15754 42818 15788
rect 42852 15754 42871 15788
rect 43689 15769 43761 15829
rect 42799 15698 42871 15754
rect 42799 15664 42818 15698
rect 42852 15664 42871 15698
rect 42799 15608 42871 15664
rect 42799 15574 42818 15608
rect 42852 15574 42871 15608
rect 42799 15518 42871 15574
rect 42799 15484 42818 15518
rect 42852 15484 42871 15518
rect 42799 15428 42871 15484
rect 42799 15394 42818 15428
rect 42852 15394 42871 15428
rect 42799 15338 42871 15394
rect 42799 15304 42818 15338
rect 42852 15304 42871 15338
rect 42799 15248 42871 15304
rect 42799 15214 42818 15248
rect 42852 15214 42871 15248
rect 42799 15158 42871 15214
rect 42799 15124 42818 15158
rect 42852 15124 42871 15158
rect 42799 15068 42871 15124
rect 43689 15735 43708 15769
rect 43742 15735 43761 15769
rect 43689 15679 43761 15735
rect 43689 15645 43708 15679
rect 43742 15645 43761 15679
rect 43689 15589 43761 15645
rect 43689 15555 43708 15589
rect 43742 15555 43761 15589
rect 43689 15499 43761 15555
rect 43689 15465 43708 15499
rect 43742 15465 43761 15499
rect 43689 15409 43761 15465
rect 43689 15375 43708 15409
rect 43742 15375 43761 15409
rect 43689 15319 43761 15375
rect 43689 15285 43708 15319
rect 43742 15285 43761 15319
rect 43689 15229 43761 15285
rect 43689 15195 43708 15229
rect 43742 15195 43761 15229
rect 43689 15139 43761 15195
rect 43689 15105 43708 15139
rect 43742 15105 43761 15139
rect 42799 15034 42818 15068
rect 42852 15034 42871 15068
rect 42799 15011 42871 15034
rect 43689 15049 43761 15105
rect 43689 15015 43708 15049
rect 43742 15015 43761 15049
rect 43689 15011 43761 15015
rect 42799 14992 43761 15011
rect 42799 14958 42876 14992
rect 42910 14958 42966 14992
rect 43000 14958 43056 14992
rect 43090 14958 43146 14992
rect 43180 14958 43236 14992
rect 43270 14958 43326 14992
rect 43360 14958 43416 14992
rect 43450 14958 43506 14992
rect 43540 14958 43596 14992
rect 43630 14958 43761 14992
rect 42799 14939 43761 14958
rect 44159 15882 45121 15901
rect 44159 15848 44270 15882
rect 44304 15848 44360 15882
rect 44394 15848 44450 15882
rect 44484 15848 44540 15882
rect 44574 15848 44630 15882
rect 44664 15848 44720 15882
rect 44754 15848 44810 15882
rect 44844 15848 44900 15882
rect 44934 15848 44990 15882
rect 45024 15848 45121 15882
rect 44159 15829 45121 15848
rect 44159 15788 44231 15829
rect 44159 15754 44178 15788
rect 44212 15754 44231 15788
rect 45049 15769 45121 15829
rect 44159 15698 44231 15754
rect 44159 15664 44178 15698
rect 44212 15664 44231 15698
rect 44159 15608 44231 15664
rect 44159 15574 44178 15608
rect 44212 15574 44231 15608
rect 44159 15518 44231 15574
rect 44159 15484 44178 15518
rect 44212 15484 44231 15518
rect 44159 15428 44231 15484
rect 44159 15394 44178 15428
rect 44212 15394 44231 15428
rect 44159 15338 44231 15394
rect 44159 15304 44178 15338
rect 44212 15304 44231 15338
rect 44159 15248 44231 15304
rect 44159 15214 44178 15248
rect 44212 15214 44231 15248
rect 44159 15158 44231 15214
rect 44159 15124 44178 15158
rect 44212 15124 44231 15158
rect 44159 15068 44231 15124
rect 45049 15735 45068 15769
rect 45102 15735 45121 15769
rect 45049 15679 45121 15735
rect 45049 15645 45068 15679
rect 45102 15645 45121 15679
rect 45049 15589 45121 15645
rect 45049 15555 45068 15589
rect 45102 15555 45121 15589
rect 45049 15499 45121 15555
rect 45049 15465 45068 15499
rect 45102 15465 45121 15499
rect 45049 15409 45121 15465
rect 45049 15375 45068 15409
rect 45102 15375 45121 15409
rect 45049 15319 45121 15375
rect 45049 15285 45068 15319
rect 45102 15285 45121 15319
rect 45049 15229 45121 15285
rect 45049 15195 45068 15229
rect 45102 15195 45121 15229
rect 45049 15139 45121 15195
rect 45049 15105 45068 15139
rect 45102 15105 45121 15139
rect 44159 15034 44178 15068
rect 44212 15034 44231 15068
rect 44159 15011 44231 15034
rect 45049 15049 45121 15105
rect 45049 15015 45068 15049
rect 45102 15015 45121 15049
rect 45049 15011 45121 15015
rect 44159 14992 45121 15011
rect 44159 14958 44236 14992
rect 44270 14958 44326 14992
rect 44360 14958 44416 14992
rect 44450 14958 44506 14992
rect 44540 14958 44596 14992
rect 44630 14958 44686 14992
rect 44720 14958 44776 14992
rect 44810 14958 44866 14992
rect 44900 14958 44956 14992
rect 44990 14958 45121 14992
rect 44159 14939 45121 14958
rect 47011 18499 47045 18561
rect 46593 15847 46627 15909
rect 47383 18555 47479 18589
rect 47739 18555 47835 18589
rect 47383 18493 47417 18555
rect 47801 18493 47835 18555
rect 47383 16527 47417 16589
rect 47801 16527 47835 16589
rect 47383 16493 47479 16527
rect 47739 16493 47835 16527
rect 47011 15847 47045 15909
rect 46593 15813 46689 15847
rect 46949 15813 47045 15847
rect 41403 14571 41499 14605
rect 45057 14571 45153 14605
rect 41403 14509 41437 14571
rect 45119 14509 45153 14571
rect 41403 14187 41437 14249
rect 45119 14187 45153 14249
rect 41403 14153 41499 14187
rect 45057 14153 45153 14187
rect 40440 11390 40520 11420
rect 40440 11350 40460 11390
rect 40500 11350 40520 11390
rect 40440 11290 40520 11350
rect 40440 11250 40460 11290
rect 40500 11250 40520 11290
rect 40440 11220 40520 11250
rect 43000 11390 43080 11420
rect 43000 11350 43020 11390
rect 43060 11350 43080 11390
rect 43000 11290 43080 11350
rect 43000 11250 43020 11290
rect 43060 11250 43080 11290
rect 43000 11220 43080 11250
rect 43480 11390 43560 11420
rect 43480 11350 43500 11390
rect 43540 11350 43560 11390
rect 43480 11290 43560 11350
rect 43480 11250 43500 11290
rect 43540 11250 43560 11290
rect 43480 11220 43560 11250
rect 46040 11390 46120 11420
rect 46040 11350 46060 11390
rect 46100 11350 46120 11390
rect 46040 11290 46120 11350
rect 46040 11250 46060 11290
rect 46100 11250 46120 11290
rect 46040 11220 46120 11250
rect 41540 10230 41620 10260
rect 41540 10190 41560 10230
rect 41600 10190 41620 10230
rect 41540 10130 41620 10190
rect 41540 10090 41560 10130
rect 41600 10090 41620 10130
rect 41540 10030 41620 10090
rect 41540 9990 41560 10030
rect 41600 9990 41620 10030
rect 41540 9930 41620 9990
rect 41540 9890 41560 9930
rect 41600 9890 41620 9930
rect 41540 9830 41620 9890
rect 41540 9790 41560 9830
rect 41600 9790 41620 9830
rect 41540 9730 41620 9790
rect 41540 9690 41560 9730
rect 41600 9690 41620 9730
rect 41540 9660 41620 9690
rect 44940 10230 45020 10260
rect 44940 10190 44960 10230
rect 45000 10190 45020 10230
rect 44940 10130 45020 10190
rect 44940 10090 44960 10130
rect 45000 10090 45020 10130
rect 44940 10030 45020 10090
rect 44940 9990 44960 10030
rect 45000 9990 45020 10030
rect 44940 9930 45020 9990
rect 44940 9890 44960 9930
rect 45000 9890 45020 9930
rect 44940 9830 45020 9890
rect 45400 10030 45480 10060
rect 45400 9990 45420 10030
rect 45460 9990 45480 10030
rect 45400 9930 45480 9990
rect 45400 9890 45420 9930
rect 45460 9890 45480 9930
rect 45400 9860 45480 9890
rect 46010 10030 46090 10060
rect 46010 9990 46030 10030
rect 46070 9990 46090 10030
rect 46010 9930 46090 9990
rect 46010 9890 46030 9930
rect 46070 9890 46090 9930
rect 46010 9860 46090 9890
rect 44940 9790 44960 9830
rect 45000 9790 45020 9830
rect 44940 9730 45020 9790
rect 44940 9690 44960 9730
rect 45000 9690 45020 9730
rect 44940 9660 45020 9690
rect 41550 9230 41630 9260
rect 41550 9190 41570 9230
rect 41610 9190 41630 9230
rect 41550 9130 41630 9190
rect 41550 9090 41570 9130
rect 41610 9090 41630 9130
rect 41550 9060 41630 9090
rect 43030 9230 43110 9260
rect 43030 9190 43050 9230
rect 43090 9190 43110 9230
rect 43030 9130 43110 9190
rect 43030 9090 43050 9130
rect 43090 9090 43110 9130
rect 43030 9060 43110 9090
rect 43450 9230 43530 9260
rect 43450 9190 43470 9230
rect 43510 9190 43530 9230
rect 43450 9130 43530 9190
rect 43450 9090 43470 9130
rect 43510 9090 43530 9130
rect 43450 9060 43530 9090
rect 44930 9230 45010 9260
rect 44930 9190 44950 9230
rect 44990 9190 45010 9230
rect 44930 9130 45010 9190
rect 44930 9090 44950 9130
rect 44990 9090 45010 9130
rect 44930 9060 45010 9090
<< psubdiffcont >>
rect 43260 19030 43300 19070
rect 43260 18950 43300 18990
rect 43260 18870 43300 18910
rect 41410 18718 41444 18752
rect 41500 18718 41534 18752
rect 41590 18718 41624 18752
rect 41680 18718 41714 18752
rect 41770 18718 41804 18752
rect 41860 18718 41894 18752
rect 41950 18718 41984 18752
rect 42040 18718 42074 18752
rect 42130 18718 42164 18752
rect 42220 18718 42254 18752
rect 42310 18718 42344 18752
rect 42400 18718 42434 18752
rect 41309 18634 41343 18668
rect 42496 18634 42530 18668
rect 41309 18544 41343 18578
rect 41309 18454 41343 18488
rect 41309 18364 41343 18398
rect 41309 18274 41343 18308
rect 41309 18184 41343 18218
rect 41309 18094 41343 18128
rect 41309 18004 41343 18038
rect 41309 17914 41343 17948
rect 41309 17824 41343 17858
rect 41309 17734 41343 17768
rect 41309 17644 41343 17678
rect 42496 18544 42530 18578
rect 42496 18454 42530 18488
rect 42496 18364 42530 18398
rect 42496 18274 42530 18308
rect 42496 18184 42530 18218
rect 42496 18094 42530 18128
rect 42496 18004 42530 18038
rect 42496 17914 42530 17948
rect 42496 17824 42530 17858
rect 42496 17734 42530 17768
rect 42496 17644 42530 17678
rect 41309 17554 41343 17588
rect 41410 17531 41444 17565
rect 41500 17531 41534 17565
rect 41590 17531 41624 17565
rect 41680 17531 41714 17565
rect 41770 17531 41804 17565
rect 41860 17531 41894 17565
rect 41950 17531 41984 17565
rect 42040 17531 42074 17565
rect 42130 17531 42164 17565
rect 42220 17531 42254 17565
rect 42310 17531 42344 17565
rect 42400 17531 42434 17565
rect 42496 17554 42530 17588
rect 42770 18718 42804 18752
rect 42860 18718 42894 18752
rect 42950 18718 42984 18752
rect 43040 18718 43074 18752
rect 43130 18718 43164 18752
rect 43220 18718 43254 18752
rect 43310 18718 43344 18752
rect 43400 18718 43434 18752
rect 43490 18718 43524 18752
rect 43580 18718 43614 18752
rect 43670 18718 43704 18752
rect 43760 18718 43794 18752
rect 42669 18634 42703 18668
rect 43856 18634 43890 18668
rect 42669 18544 42703 18578
rect 42669 18454 42703 18488
rect 42669 18364 42703 18398
rect 42669 18274 42703 18308
rect 42669 18184 42703 18218
rect 42669 18094 42703 18128
rect 42669 18004 42703 18038
rect 42669 17914 42703 17948
rect 42669 17824 42703 17858
rect 42669 17734 42703 17768
rect 42669 17644 42703 17678
rect 43856 18544 43890 18578
rect 43856 18454 43890 18488
rect 43856 18364 43890 18398
rect 43856 18274 43890 18308
rect 43856 18184 43890 18218
rect 43856 18094 43890 18128
rect 43856 18004 43890 18038
rect 43856 17914 43890 17948
rect 43856 17824 43890 17858
rect 43856 17734 43890 17768
rect 43856 17644 43890 17678
rect 42669 17554 42703 17588
rect 42770 17531 42804 17565
rect 42860 17531 42894 17565
rect 42950 17531 42984 17565
rect 43040 17531 43074 17565
rect 43130 17531 43164 17565
rect 43220 17531 43254 17565
rect 43310 17531 43344 17565
rect 43400 17531 43434 17565
rect 43490 17531 43524 17565
rect 43580 17531 43614 17565
rect 43670 17531 43704 17565
rect 43760 17531 43794 17565
rect 43856 17554 43890 17588
rect 44130 18718 44164 18752
rect 44220 18718 44254 18752
rect 44310 18718 44344 18752
rect 44400 18718 44434 18752
rect 44490 18718 44524 18752
rect 44580 18718 44614 18752
rect 44670 18718 44704 18752
rect 44760 18718 44794 18752
rect 44850 18718 44884 18752
rect 44940 18718 44974 18752
rect 45030 18718 45064 18752
rect 45120 18718 45154 18752
rect 44029 18634 44063 18668
rect 45216 18634 45250 18668
rect 44029 18544 44063 18578
rect 44029 18454 44063 18488
rect 44029 18364 44063 18398
rect 44029 18274 44063 18308
rect 44029 18184 44063 18218
rect 44029 18094 44063 18128
rect 44029 18004 44063 18038
rect 44029 17914 44063 17948
rect 44029 17824 44063 17858
rect 44029 17734 44063 17768
rect 44029 17644 44063 17678
rect 45216 18544 45250 18578
rect 45216 18454 45250 18488
rect 45216 18364 45250 18398
rect 45216 18274 45250 18308
rect 45216 18184 45250 18218
rect 45216 18094 45250 18128
rect 45216 18004 45250 18038
rect 45216 17914 45250 17948
rect 45216 17824 45250 17858
rect 45216 17734 45250 17768
rect 45216 17644 45250 17678
rect 44029 17554 44063 17588
rect 44130 17531 44164 17565
rect 44220 17531 44254 17565
rect 44310 17531 44344 17565
rect 44400 17531 44434 17565
rect 44490 17531 44524 17565
rect 44580 17531 44614 17565
rect 44670 17531 44704 17565
rect 44760 17531 44794 17565
rect 44850 17531 44884 17565
rect 44940 17531 44974 17565
rect 45030 17531 45064 17565
rect 45120 17531 45154 17565
rect 45216 17554 45250 17588
rect 41410 17358 41444 17392
rect 41500 17358 41534 17392
rect 41590 17358 41624 17392
rect 41680 17358 41714 17392
rect 41770 17358 41804 17392
rect 41860 17358 41894 17392
rect 41950 17358 41984 17392
rect 42040 17358 42074 17392
rect 42130 17358 42164 17392
rect 42220 17358 42254 17392
rect 42310 17358 42344 17392
rect 42400 17358 42434 17392
rect 41309 17274 41343 17308
rect 42496 17274 42530 17308
rect 41309 17184 41343 17218
rect 41309 17094 41343 17128
rect 41309 17004 41343 17038
rect 41309 16914 41343 16948
rect 41309 16824 41343 16858
rect 41309 16734 41343 16768
rect 41309 16644 41343 16678
rect 41309 16554 41343 16588
rect 41309 16464 41343 16498
rect 41309 16374 41343 16408
rect 41309 16284 41343 16318
rect 42496 17184 42530 17218
rect 42496 17094 42530 17128
rect 42496 17004 42530 17038
rect 42496 16914 42530 16948
rect 42496 16824 42530 16858
rect 42496 16734 42530 16768
rect 42496 16644 42530 16678
rect 42496 16554 42530 16588
rect 42496 16464 42530 16498
rect 42496 16374 42530 16408
rect 42496 16284 42530 16318
rect 41309 16194 41343 16228
rect 41410 16171 41444 16205
rect 41500 16171 41534 16205
rect 41590 16171 41624 16205
rect 41680 16171 41714 16205
rect 41770 16171 41804 16205
rect 41860 16171 41894 16205
rect 41950 16171 41984 16205
rect 42040 16171 42074 16205
rect 42130 16171 42164 16205
rect 42220 16171 42254 16205
rect 42310 16171 42344 16205
rect 42400 16171 42434 16205
rect 42496 16194 42530 16228
rect 42770 17358 42804 17392
rect 42860 17358 42894 17392
rect 42950 17358 42984 17392
rect 43040 17358 43074 17392
rect 43130 17358 43164 17392
rect 43220 17358 43254 17392
rect 43310 17358 43344 17392
rect 43400 17358 43434 17392
rect 43490 17358 43524 17392
rect 43580 17358 43614 17392
rect 43670 17358 43704 17392
rect 43760 17358 43794 17392
rect 42669 17274 42703 17308
rect 43856 17274 43890 17308
rect 42669 17184 42703 17218
rect 42669 17094 42703 17128
rect 42669 17004 42703 17038
rect 42669 16914 42703 16948
rect 42669 16824 42703 16858
rect 42669 16734 42703 16768
rect 42669 16644 42703 16678
rect 42669 16554 42703 16588
rect 42669 16464 42703 16498
rect 42669 16374 42703 16408
rect 42669 16284 42703 16318
rect 43856 17184 43890 17218
rect 43856 17094 43890 17128
rect 43856 17004 43890 17038
rect 43856 16914 43890 16948
rect 43856 16824 43890 16858
rect 43856 16734 43890 16768
rect 43856 16644 43890 16678
rect 43856 16554 43890 16588
rect 43856 16464 43890 16498
rect 43856 16374 43890 16408
rect 43856 16284 43890 16318
rect 42669 16194 42703 16228
rect 42770 16171 42804 16205
rect 42860 16171 42894 16205
rect 42950 16171 42984 16205
rect 43040 16171 43074 16205
rect 43130 16171 43164 16205
rect 43220 16171 43254 16205
rect 43310 16171 43344 16205
rect 43400 16171 43434 16205
rect 43490 16171 43524 16205
rect 43580 16171 43614 16205
rect 43670 16171 43704 16205
rect 43760 16171 43794 16205
rect 43856 16194 43890 16228
rect 44130 17358 44164 17392
rect 44220 17358 44254 17392
rect 44310 17358 44344 17392
rect 44400 17358 44434 17392
rect 44490 17358 44524 17392
rect 44580 17358 44614 17392
rect 44670 17358 44704 17392
rect 44760 17358 44794 17392
rect 44850 17358 44884 17392
rect 44940 17358 44974 17392
rect 45030 17358 45064 17392
rect 45120 17358 45154 17392
rect 44029 17274 44063 17308
rect 45216 17274 45250 17308
rect 44029 17184 44063 17218
rect 44029 17094 44063 17128
rect 44029 17004 44063 17038
rect 44029 16914 44063 16948
rect 44029 16824 44063 16858
rect 44029 16734 44063 16768
rect 44029 16644 44063 16678
rect 44029 16554 44063 16588
rect 44029 16464 44063 16498
rect 44029 16374 44063 16408
rect 44029 16284 44063 16318
rect 45216 17184 45250 17218
rect 45216 17094 45250 17128
rect 45216 17004 45250 17038
rect 45216 16914 45250 16948
rect 45216 16824 45250 16858
rect 45216 16734 45250 16768
rect 45216 16644 45250 16678
rect 45216 16554 45250 16588
rect 45216 16464 45250 16498
rect 45216 16374 45250 16408
rect 45216 16284 45250 16318
rect 44029 16194 44063 16228
rect 44130 16171 44164 16205
rect 44220 16171 44254 16205
rect 44310 16171 44344 16205
rect 44400 16171 44434 16205
rect 44490 16171 44524 16205
rect 44580 16171 44614 16205
rect 44670 16171 44704 16205
rect 44760 16171 44794 16205
rect 44850 16171 44884 16205
rect 44940 16171 44974 16205
rect 45030 16171 45064 16205
rect 45120 16171 45154 16205
rect 45216 16194 45250 16228
rect 41410 15998 41444 16032
rect 41500 15998 41534 16032
rect 41590 15998 41624 16032
rect 41680 15998 41714 16032
rect 41770 15998 41804 16032
rect 41860 15998 41894 16032
rect 41950 15998 41984 16032
rect 42040 15998 42074 16032
rect 42130 15998 42164 16032
rect 42220 15998 42254 16032
rect 42310 15998 42344 16032
rect 42400 15998 42434 16032
rect 41309 15914 41343 15948
rect 42496 15914 42530 15948
rect 41309 15824 41343 15858
rect 41309 15734 41343 15768
rect 41309 15644 41343 15678
rect 41309 15554 41343 15588
rect 41309 15464 41343 15498
rect 41309 15374 41343 15408
rect 41309 15284 41343 15318
rect 41309 15194 41343 15228
rect 41309 15104 41343 15138
rect 41309 15014 41343 15048
rect 41309 14924 41343 14958
rect 42496 15824 42530 15858
rect 42496 15734 42530 15768
rect 42496 15644 42530 15678
rect 42496 15554 42530 15588
rect 42496 15464 42530 15498
rect 42496 15374 42530 15408
rect 42496 15284 42530 15318
rect 42496 15194 42530 15228
rect 42496 15104 42530 15138
rect 42496 15014 42530 15048
rect 42496 14924 42530 14958
rect 41309 14834 41343 14868
rect 41410 14811 41444 14845
rect 41500 14811 41534 14845
rect 41590 14811 41624 14845
rect 41680 14811 41714 14845
rect 41770 14811 41804 14845
rect 41860 14811 41894 14845
rect 41950 14811 41984 14845
rect 42040 14811 42074 14845
rect 42130 14811 42164 14845
rect 42220 14811 42254 14845
rect 42310 14811 42344 14845
rect 42400 14811 42434 14845
rect 42496 14834 42530 14868
rect 42770 15998 42804 16032
rect 42860 15998 42894 16032
rect 42950 15998 42984 16032
rect 43040 15998 43074 16032
rect 43130 15998 43164 16032
rect 43220 15998 43254 16032
rect 43310 15998 43344 16032
rect 43400 15998 43434 16032
rect 43490 15998 43524 16032
rect 43580 15998 43614 16032
rect 43670 15998 43704 16032
rect 43760 15998 43794 16032
rect 42669 15914 42703 15948
rect 43856 15914 43890 15948
rect 42669 15824 42703 15858
rect 42669 15734 42703 15768
rect 42669 15644 42703 15678
rect 42669 15554 42703 15588
rect 42669 15464 42703 15498
rect 42669 15374 42703 15408
rect 42669 15284 42703 15318
rect 42669 15194 42703 15228
rect 42669 15104 42703 15138
rect 42669 15014 42703 15048
rect 42669 14924 42703 14958
rect 43856 15824 43890 15858
rect 43856 15734 43890 15768
rect 43856 15644 43890 15678
rect 43856 15554 43890 15588
rect 43856 15464 43890 15498
rect 43856 15374 43890 15408
rect 43856 15284 43890 15318
rect 43856 15194 43890 15228
rect 43856 15104 43890 15138
rect 43856 15014 43890 15048
rect 43856 14924 43890 14958
rect 42669 14834 42703 14868
rect 42770 14811 42804 14845
rect 42860 14811 42894 14845
rect 42950 14811 42984 14845
rect 43040 14811 43074 14845
rect 43130 14811 43164 14845
rect 43220 14811 43254 14845
rect 43310 14811 43344 14845
rect 43400 14811 43434 14845
rect 43490 14811 43524 14845
rect 43580 14811 43614 14845
rect 43670 14811 43704 14845
rect 43760 14811 43794 14845
rect 43856 14834 43890 14868
rect 44130 15998 44164 16032
rect 44220 15998 44254 16032
rect 44310 15998 44344 16032
rect 44400 15998 44434 16032
rect 44490 15998 44524 16032
rect 44580 15998 44614 16032
rect 44670 15998 44704 16032
rect 44760 15998 44794 16032
rect 44850 15998 44884 16032
rect 44940 15998 44974 16032
rect 45030 15998 45064 16032
rect 45120 15998 45154 16032
rect 44029 15914 44063 15948
rect 45216 15914 45250 15948
rect 44029 15824 44063 15858
rect 44029 15734 44063 15768
rect 44029 15644 44063 15678
rect 44029 15554 44063 15588
rect 44029 15464 44063 15498
rect 44029 15374 44063 15408
rect 44029 15284 44063 15318
rect 44029 15194 44063 15228
rect 44029 15104 44063 15138
rect 44029 15014 44063 15048
rect 44029 14924 44063 14958
rect 45216 15824 45250 15858
rect 45216 15734 45250 15768
rect 45216 15644 45250 15678
rect 45216 15554 45250 15588
rect 45216 15464 45250 15498
rect 45216 15374 45250 15408
rect 45216 15284 45250 15318
rect 45216 15194 45250 15228
rect 45216 15104 45250 15138
rect 45216 15014 45250 15048
rect 45216 14924 45250 14958
rect 44029 14834 44063 14868
rect 44130 14811 44164 14845
rect 44220 14811 44254 14845
rect 44310 14811 44344 14845
rect 44400 14811 44434 14845
rect 44490 14811 44524 14845
rect 44580 14811 44614 14845
rect 44670 14811 44704 14845
rect 44760 14811 44794 14845
rect 44850 14811 44884 14845
rect 44940 14811 44974 14845
rect 45030 14811 45064 14845
rect 45120 14811 45154 14845
rect 45216 14834 45250 14868
rect 45420 13810 45460 13850
rect 45420 13710 45460 13750
rect 41920 13200 41960 13240
rect 41920 13100 41960 13140
rect 41920 13000 41960 13040
rect 41920 12900 41960 12940
rect 41920 12800 41960 12840
rect 44600 13200 44640 13240
rect 44600 13100 44640 13140
rect 44600 13000 44640 13040
rect 44600 12900 44640 12940
rect 44600 12800 44640 12840
rect 42820 12280 42860 12320
rect 42820 12200 42860 12240
rect 42820 12120 42860 12160
rect 43700 12280 43740 12320
rect 43700 12200 43740 12240
rect 43700 12120 43740 12160
<< nsubdiffcont >>
rect 38699 18555 38959 18589
rect 38603 16589 38637 18493
rect 39021 16589 39055 18493
rect 38699 16493 38959 16527
rect 39479 18561 39739 18595
rect 39383 15019 39417 18499
rect 39801 15019 39835 18499
rect 40259 18563 40851 18597
rect 40163 16243 40197 18501
rect 40913 16243 40947 18501
rect 41550 18568 41584 18602
rect 41640 18568 41674 18602
rect 41730 18568 41764 18602
rect 41820 18568 41854 18602
rect 41910 18568 41944 18602
rect 42000 18568 42034 18602
rect 42090 18568 42124 18602
rect 42180 18568 42214 18602
rect 42270 18568 42304 18602
rect 41458 18474 41492 18508
rect 41458 18384 41492 18418
rect 41458 18294 41492 18328
rect 41458 18204 41492 18238
rect 41458 18114 41492 18148
rect 41458 18024 41492 18058
rect 41458 17934 41492 17968
rect 41458 17844 41492 17878
rect 42348 18455 42382 18489
rect 42348 18365 42382 18399
rect 42348 18275 42382 18309
rect 42348 18185 42382 18219
rect 42348 18095 42382 18129
rect 42348 18005 42382 18039
rect 42348 17915 42382 17949
rect 42348 17825 42382 17859
rect 41458 17754 41492 17788
rect 42348 17735 42382 17769
rect 41516 17678 41550 17712
rect 41606 17678 41640 17712
rect 41696 17678 41730 17712
rect 41786 17678 41820 17712
rect 41876 17678 41910 17712
rect 41966 17678 42000 17712
rect 42056 17678 42090 17712
rect 42146 17678 42180 17712
rect 42236 17678 42270 17712
rect 42910 18568 42944 18602
rect 43000 18568 43034 18602
rect 43090 18568 43124 18602
rect 43180 18568 43214 18602
rect 43270 18568 43304 18602
rect 43360 18568 43394 18602
rect 43450 18568 43484 18602
rect 43540 18568 43574 18602
rect 43630 18568 43664 18602
rect 42818 18474 42852 18508
rect 42818 18384 42852 18418
rect 42818 18294 42852 18328
rect 42818 18204 42852 18238
rect 42818 18114 42852 18148
rect 42818 18024 42852 18058
rect 42818 17934 42852 17968
rect 42818 17844 42852 17878
rect 43708 18455 43742 18489
rect 43708 18365 43742 18399
rect 43708 18275 43742 18309
rect 43708 18185 43742 18219
rect 43708 18095 43742 18129
rect 43708 18005 43742 18039
rect 43708 17915 43742 17949
rect 43708 17825 43742 17859
rect 42818 17754 42852 17788
rect 43708 17735 43742 17769
rect 42876 17678 42910 17712
rect 42966 17678 43000 17712
rect 43056 17678 43090 17712
rect 43146 17678 43180 17712
rect 43236 17678 43270 17712
rect 43326 17678 43360 17712
rect 43416 17678 43450 17712
rect 43506 17678 43540 17712
rect 43596 17678 43630 17712
rect 44270 18568 44304 18602
rect 44360 18568 44394 18602
rect 44450 18568 44484 18602
rect 44540 18568 44574 18602
rect 44630 18568 44664 18602
rect 44720 18568 44754 18602
rect 44810 18568 44844 18602
rect 44900 18568 44934 18602
rect 44990 18568 45024 18602
rect 44178 18474 44212 18508
rect 44178 18384 44212 18418
rect 44178 18294 44212 18328
rect 44178 18204 44212 18238
rect 44178 18114 44212 18148
rect 44178 18024 44212 18058
rect 44178 17934 44212 17968
rect 44178 17844 44212 17878
rect 45068 18455 45102 18489
rect 45068 18365 45102 18399
rect 45068 18275 45102 18309
rect 45068 18185 45102 18219
rect 45068 18095 45102 18129
rect 45068 18005 45102 18039
rect 45068 17915 45102 17949
rect 45068 17825 45102 17859
rect 44178 17754 44212 17788
rect 45068 17735 45102 17769
rect 44236 17678 44270 17712
rect 44326 17678 44360 17712
rect 44416 17678 44450 17712
rect 44506 17678 44540 17712
rect 44596 17678 44630 17712
rect 44686 17678 44720 17712
rect 44776 17678 44810 17712
rect 44866 17678 44900 17712
rect 44956 17678 44990 17712
rect 45579 18563 46171 18597
rect 40259 16147 40851 16181
rect 41550 17208 41584 17242
rect 41640 17208 41674 17242
rect 41730 17208 41764 17242
rect 41820 17208 41854 17242
rect 41910 17208 41944 17242
rect 42000 17208 42034 17242
rect 42090 17208 42124 17242
rect 42180 17208 42214 17242
rect 42270 17208 42304 17242
rect 41458 17114 41492 17148
rect 41458 17024 41492 17058
rect 41458 16934 41492 16968
rect 41458 16844 41492 16878
rect 41458 16754 41492 16788
rect 41458 16664 41492 16698
rect 41458 16574 41492 16608
rect 41458 16484 41492 16518
rect 42348 17095 42382 17129
rect 42348 17005 42382 17039
rect 42348 16915 42382 16949
rect 42348 16825 42382 16859
rect 42348 16735 42382 16769
rect 42348 16645 42382 16679
rect 42348 16555 42382 16589
rect 42348 16465 42382 16499
rect 41458 16394 41492 16428
rect 42348 16375 42382 16409
rect 41516 16318 41550 16352
rect 41606 16318 41640 16352
rect 41696 16318 41730 16352
rect 41786 16318 41820 16352
rect 41876 16318 41910 16352
rect 41966 16318 42000 16352
rect 42056 16318 42090 16352
rect 42146 16318 42180 16352
rect 42236 16318 42270 16352
rect 42910 17208 42944 17242
rect 43000 17208 43034 17242
rect 43090 17208 43124 17242
rect 43180 17208 43214 17242
rect 43270 17208 43304 17242
rect 43360 17208 43394 17242
rect 43450 17208 43484 17242
rect 43540 17208 43574 17242
rect 43630 17208 43664 17242
rect 42818 17114 42852 17148
rect 42818 17024 42852 17058
rect 42818 16934 42852 16968
rect 42818 16844 42852 16878
rect 42818 16754 42852 16788
rect 42818 16664 42852 16698
rect 42818 16574 42852 16608
rect 42818 16484 42852 16518
rect 43708 17095 43742 17129
rect 43708 17005 43742 17039
rect 43708 16915 43742 16949
rect 43708 16825 43742 16859
rect 43708 16735 43742 16769
rect 43708 16645 43742 16679
rect 43708 16555 43742 16589
rect 43708 16465 43742 16499
rect 42818 16394 42852 16428
rect 43708 16375 43742 16409
rect 42876 16318 42910 16352
rect 42966 16318 43000 16352
rect 43056 16318 43090 16352
rect 43146 16318 43180 16352
rect 43236 16318 43270 16352
rect 43326 16318 43360 16352
rect 43416 16318 43450 16352
rect 43506 16318 43540 16352
rect 43596 16318 43630 16352
rect 44270 17208 44304 17242
rect 44360 17208 44394 17242
rect 44450 17208 44484 17242
rect 44540 17208 44574 17242
rect 44630 17208 44664 17242
rect 44720 17208 44754 17242
rect 44810 17208 44844 17242
rect 44900 17208 44934 17242
rect 44990 17208 45024 17242
rect 44178 17114 44212 17148
rect 44178 17024 44212 17058
rect 44178 16934 44212 16968
rect 44178 16844 44212 16878
rect 44178 16754 44212 16788
rect 44178 16664 44212 16698
rect 44178 16574 44212 16608
rect 44178 16484 44212 16518
rect 45068 17095 45102 17129
rect 45068 17005 45102 17039
rect 45068 16915 45102 16949
rect 45068 16825 45102 16859
rect 45068 16735 45102 16769
rect 45068 16645 45102 16679
rect 45068 16555 45102 16589
rect 45068 16465 45102 16499
rect 44178 16394 44212 16428
rect 45068 16375 45102 16409
rect 44236 16318 44270 16352
rect 44326 16318 44360 16352
rect 44416 16318 44450 16352
rect 44506 16318 44540 16352
rect 44596 16318 44630 16352
rect 44686 16318 44720 16352
rect 44776 16318 44810 16352
rect 44866 16318 44900 16352
rect 44956 16318 44990 16352
rect 45483 16243 45517 18501
rect 46233 16243 46267 18501
rect 45579 16147 46171 16181
rect 46689 18561 46949 18595
rect 39479 14923 39739 14957
rect 41550 15848 41584 15882
rect 41640 15848 41674 15882
rect 41730 15848 41764 15882
rect 41820 15848 41854 15882
rect 41910 15848 41944 15882
rect 42000 15848 42034 15882
rect 42090 15848 42124 15882
rect 42180 15848 42214 15882
rect 42270 15848 42304 15882
rect 41458 15754 41492 15788
rect 41458 15664 41492 15698
rect 41458 15574 41492 15608
rect 41458 15484 41492 15518
rect 41458 15394 41492 15428
rect 41458 15304 41492 15338
rect 41458 15214 41492 15248
rect 41458 15124 41492 15158
rect 42348 15735 42382 15769
rect 42348 15645 42382 15679
rect 42348 15555 42382 15589
rect 42348 15465 42382 15499
rect 42348 15375 42382 15409
rect 42348 15285 42382 15319
rect 42348 15195 42382 15229
rect 42348 15105 42382 15139
rect 41458 15034 41492 15068
rect 42348 15015 42382 15049
rect 41516 14958 41550 14992
rect 41606 14958 41640 14992
rect 41696 14958 41730 14992
rect 41786 14958 41820 14992
rect 41876 14958 41910 14992
rect 41966 14958 42000 14992
rect 42056 14958 42090 14992
rect 42146 14958 42180 14992
rect 42236 14958 42270 14992
rect 42910 15848 42944 15882
rect 43000 15848 43034 15882
rect 43090 15848 43124 15882
rect 43180 15848 43214 15882
rect 43270 15848 43304 15882
rect 43360 15848 43394 15882
rect 43450 15848 43484 15882
rect 43540 15848 43574 15882
rect 43630 15848 43664 15882
rect 42818 15754 42852 15788
rect 42818 15664 42852 15698
rect 42818 15574 42852 15608
rect 42818 15484 42852 15518
rect 42818 15394 42852 15428
rect 42818 15304 42852 15338
rect 42818 15214 42852 15248
rect 42818 15124 42852 15158
rect 43708 15735 43742 15769
rect 43708 15645 43742 15679
rect 43708 15555 43742 15589
rect 43708 15465 43742 15499
rect 43708 15375 43742 15409
rect 43708 15285 43742 15319
rect 43708 15195 43742 15229
rect 43708 15105 43742 15139
rect 42818 15034 42852 15068
rect 43708 15015 43742 15049
rect 42876 14958 42910 14992
rect 42966 14958 43000 14992
rect 43056 14958 43090 14992
rect 43146 14958 43180 14992
rect 43236 14958 43270 14992
rect 43326 14958 43360 14992
rect 43416 14958 43450 14992
rect 43506 14958 43540 14992
rect 43596 14958 43630 14992
rect 44270 15848 44304 15882
rect 44360 15848 44394 15882
rect 44450 15848 44484 15882
rect 44540 15848 44574 15882
rect 44630 15848 44664 15882
rect 44720 15848 44754 15882
rect 44810 15848 44844 15882
rect 44900 15848 44934 15882
rect 44990 15848 45024 15882
rect 44178 15754 44212 15788
rect 44178 15664 44212 15698
rect 44178 15574 44212 15608
rect 44178 15484 44212 15518
rect 44178 15394 44212 15428
rect 44178 15304 44212 15338
rect 44178 15214 44212 15248
rect 44178 15124 44212 15158
rect 45068 15735 45102 15769
rect 45068 15645 45102 15679
rect 45068 15555 45102 15589
rect 45068 15465 45102 15499
rect 45068 15375 45102 15409
rect 45068 15285 45102 15319
rect 45068 15195 45102 15229
rect 45068 15105 45102 15139
rect 44178 15034 44212 15068
rect 45068 15015 45102 15049
rect 44236 14958 44270 14992
rect 44326 14958 44360 14992
rect 44416 14958 44450 14992
rect 44506 14958 44540 14992
rect 44596 14958 44630 14992
rect 44686 14958 44720 14992
rect 44776 14958 44810 14992
rect 44866 14958 44900 14992
rect 44956 14958 44990 14992
rect 46593 15909 46627 18499
rect 47011 15909 47045 18499
rect 47479 18555 47739 18589
rect 47383 16589 47417 18493
rect 47801 16589 47835 18493
rect 47479 16493 47739 16527
rect 46689 15813 46949 15847
rect 41499 14571 45057 14605
rect 41403 14249 41437 14509
rect 45119 14249 45153 14509
rect 41499 14153 45057 14187
rect 40460 11350 40500 11390
rect 40460 11250 40500 11290
rect 43020 11350 43060 11390
rect 43020 11250 43060 11290
rect 43500 11350 43540 11390
rect 43500 11250 43540 11290
rect 46060 11350 46100 11390
rect 46060 11250 46100 11290
rect 41560 10190 41600 10230
rect 41560 10090 41600 10130
rect 41560 9990 41600 10030
rect 41560 9890 41600 9930
rect 41560 9790 41600 9830
rect 41560 9690 41600 9730
rect 44960 10190 45000 10230
rect 44960 10090 45000 10130
rect 44960 9990 45000 10030
rect 44960 9890 45000 9930
rect 45420 9990 45460 10030
rect 45420 9890 45460 9930
rect 46030 9990 46070 10030
rect 46030 9890 46070 9930
rect 44960 9790 45000 9830
rect 44960 9690 45000 9730
rect 41570 9190 41610 9230
rect 41570 9090 41610 9130
rect 43050 9190 43090 9230
rect 43050 9090 43090 9130
rect 43470 9190 43510 9230
rect 43470 9090 43510 9130
rect 44950 9190 44990 9230
rect 44950 9090 44990 9130
<< poly >>
rect 41240 13880 43240 13910
rect 43320 13880 45320 13910
rect 41240 13650 43240 13680
rect 43320 13650 45320 13680
rect 41320 13630 41400 13650
rect 41320 13590 41340 13630
rect 41380 13590 41400 13630
rect 41320 13570 41400 13590
rect 41480 13630 41560 13650
rect 41480 13590 41500 13630
rect 41540 13590 41560 13630
rect 41480 13570 41560 13590
rect 41640 13630 41720 13650
rect 41640 13590 41660 13630
rect 41700 13590 41720 13630
rect 41640 13570 41720 13590
rect 41800 13630 41880 13650
rect 41800 13590 41820 13630
rect 41860 13590 41880 13630
rect 41800 13570 41880 13590
rect 41960 13630 42040 13650
rect 41960 13590 41980 13630
rect 42020 13590 42040 13630
rect 41960 13570 42040 13590
rect 42120 13630 42200 13650
rect 42120 13590 42140 13630
rect 42180 13590 42200 13630
rect 42120 13570 42200 13590
rect 42280 13630 42360 13650
rect 42280 13590 42300 13630
rect 42340 13590 42360 13630
rect 42280 13570 42360 13590
rect 42440 13630 42520 13650
rect 42440 13590 42460 13630
rect 42500 13590 42520 13630
rect 42440 13570 42520 13590
rect 42600 13630 42680 13650
rect 42600 13590 42620 13630
rect 42660 13590 42680 13630
rect 42600 13570 42680 13590
rect 42760 13630 42840 13650
rect 42760 13590 42780 13630
rect 42820 13590 42840 13630
rect 42760 13570 42840 13590
rect 42920 13630 43000 13650
rect 42920 13590 42940 13630
rect 42980 13590 43000 13630
rect 42920 13570 43000 13590
rect 43080 13630 43160 13650
rect 43080 13590 43100 13630
rect 43140 13590 43160 13630
rect 43080 13570 43160 13590
rect 43400 13630 43480 13650
rect 43400 13590 43420 13630
rect 43460 13590 43480 13630
rect 43400 13570 43480 13590
rect 43560 13630 43640 13650
rect 43560 13590 43580 13630
rect 43620 13590 43640 13630
rect 43560 13570 43640 13590
rect 43720 13630 43800 13650
rect 43720 13590 43740 13630
rect 43780 13590 43800 13630
rect 43720 13570 43800 13590
rect 43880 13630 43960 13650
rect 43880 13590 43900 13630
rect 43940 13590 43960 13630
rect 43880 13570 43960 13590
rect 44040 13630 44120 13650
rect 44040 13590 44060 13630
rect 44100 13590 44120 13630
rect 44040 13570 44120 13590
rect 44200 13630 44280 13650
rect 44200 13590 44220 13630
rect 44260 13590 44280 13630
rect 44200 13570 44280 13590
rect 44360 13630 44440 13650
rect 44360 13590 44380 13630
rect 44420 13590 44440 13630
rect 44360 13570 44440 13590
rect 44520 13630 44600 13650
rect 44520 13590 44540 13630
rect 44580 13590 44600 13630
rect 44520 13570 44600 13590
rect 44680 13630 44760 13650
rect 44680 13590 44700 13630
rect 44740 13590 44760 13630
rect 44680 13570 44760 13590
rect 44840 13630 44920 13650
rect 44840 13590 44860 13630
rect 44900 13590 44920 13630
rect 44840 13570 44920 13590
rect 45000 13630 45080 13650
rect 45000 13590 45020 13630
rect 45060 13590 45080 13630
rect 45000 13570 45080 13590
rect 45160 13630 45240 13650
rect 45160 13590 45180 13630
rect 45220 13590 45240 13630
rect 45160 13570 45240 13590
rect 40820 13270 41820 13300
rect 42060 13270 43060 13300
rect 43500 13270 44500 13300
rect 44740 13270 45740 13300
rect 40820 12740 41820 12770
rect 42060 12740 43060 12770
rect 43500 12740 44500 12770
rect 44740 12740 45740 12770
rect 40920 12720 41000 12740
rect 40920 12680 40940 12720
rect 40980 12680 41000 12720
rect 40920 12660 41000 12680
rect 41160 12720 41240 12740
rect 41160 12680 41180 12720
rect 41220 12680 41240 12720
rect 41160 12660 41240 12680
rect 41400 12720 41480 12740
rect 41400 12680 41420 12720
rect 41460 12680 41480 12720
rect 41400 12660 41480 12680
rect 41640 12720 41720 12740
rect 41640 12680 41660 12720
rect 41700 12680 41720 12720
rect 41640 12660 41720 12680
rect 42280 12720 42360 12740
rect 42280 12680 42300 12720
rect 42340 12680 42360 12720
rect 42280 12660 42360 12680
rect 42520 12720 42600 12740
rect 42520 12680 42540 12720
rect 42580 12680 42600 12720
rect 42520 12660 42600 12680
rect 42760 12720 42840 12740
rect 42760 12680 42780 12720
rect 42820 12680 42840 12720
rect 42760 12660 42840 12680
rect 43720 12720 43800 12740
rect 43720 12680 43740 12720
rect 43780 12680 43800 12720
rect 43720 12660 43800 12680
rect 43960 12720 44040 12740
rect 43960 12680 43980 12720
rect 44020 12680 44040 12720
rect 43960 12660 44040 12680
rect 44200 12720 44280 12740
rect 44200 12680 44220 12720
rect 44260 12680 44280 12720
rect 44200 12660 44280 12680
rect 44840 12720 44920 12740
rect 44840 12680 44860 12720
rect 44900 12680 44920 12720
rect 44840 12660 44920 12680
rect 45080 12720 45160 12740
rect 45080 12680 45100 12720
rect 45140 12680 45160 12720
rect 45080 12660 45160 12680
rect 45320 12720 45400 12740
rect 45320 12680 45340 12720
rect 45380 12680 45400 12720
rect 45320 12660 45400 12680
rect 45560 12720 45640 12740
rect 45560 12680 45580 12720
rect 45620 12680 45640 12720
rect 45560 12660 45640 12680
rect 41431 12342 41489 12360
rect 41431 12308 41443 12342
rect 41477 12308 41489 12342
rect 41431 12290 41489 12308
rect 41791 12342 41849 12360
rect 41791 12308 41803 12342
rect 41837 12308 41849 12342
rect 41791 12290 41849 12308
rect 41911 12342 41969 12360
rect 41911 12308 41923 12342
rect 41957 12308 41969 12342
rect 41911 12290 41969 12308
rect 42271 12342 42329 12360
rect 42271 12308 42283 12342
rect 42317 12308 42329 12342
rect 42271 12290 42329 12308
rect 42391 12342 42449 12360
rect 42391 12308 42403 12342
rect 42437 12308 42449 12342
rect 42391 12290 42449 12308
rect 41440 12260 41480 12290
rect 41560 12260 41600 12290
rect 41680 12260 41720 12290
rect 41800 12260 41840 12290
rect 41920 12260 41960 12290
rect 42040 12260 42080 12290
rect 42160 12260 42200 12290
rect 42280 12260 42320 12290
rect 42400 12260 42440 12290
rect 42520 12260 42560 12290
rect 41440 12130 41480 12160
rect 41560 12130 41600 12160
rect 41532 12112 41600 12130
rect 41532 12078 41544 12112
rect 41578 12078 41600 12112
rect 41532 12060 41600 12078
rect 41680 12130 41720 12160
rect 41800 12130 41840 12160
rect 41920 12130 41960 12160
rect 42040 12130 42080 12160
rect 41680 12112 41748 12130
rect 41680 12078 41702 12112
rect 41736 12078 41748 12112
rect 41680 12060 41748 12078
rect 42014 12112 42080 12130
rect 42014 12078 42026 12112
rect 42060 12078 42080 12112
rect 42014 12060 42080 12078
rect 42160 12130 42200 12160
rect 42280 12130 42320 12160
rect 42400 12130 42440 12160
rect 42520 12130 42560 12160
rect 42160 12112 42226 12130
rect 42160 12078 42180 12112
rect 42214 12078 42226 12112
rect 42160 12060 42226 12078
rect 42492 12112 42560 12130
rect 42492 12078 42504 12112
rect 42538 12078 42560 12112
rect 44111 12342 44169 12360
rect 44111 12308 44123 12342
rect 44157 12308 44169 12342
rect 44111 12290 44169 12308
rect 44231 12342 44289 12360
rect 44231 12308 44243 12342
rect 44277 12308 44289 12342
rect 44231 12290 44289 12308
rect 44591 12342 44649 12360
rect 44591 12308 44603 12342
rect 44637 12308 44649 12342
rect 44591 12290 44649 12308
rect 44711 12342 44769 12360
rect 44711 12308 44723 12342
rect 44757 12308 44769 12342
rect 44711 12290 44769 12308
rect 45071 12342 45129 12360
rect 45071 12308 45083 12342
rect 45117 12308 45129 12342
rect 45071 12290 45129 12308
rect 44000 12260 44040 12290
rect 44120 12260 44160 12290
rect 44240 12260 44280 12290
rect 44360 12260 44400 12290
rect 44480 12260 44520 12290
rect 44600 12260 44640 12290
rect 44720 12260 44760 12290
rect 44840 12260 44880 12290
rect 44960 12260 45000 12290
rect 45080 12260 45120 12290
rect 44000 12130 44040 12160
rect 44120 12130 44160 12160
rect 44240 12130 44280 12160
rect 44360 12130 44400 12160
rect 44000 12112 44068 12130
rect 42492 12060 42560 12078
rect 44000 12078 44022 12112
rect 44056 12078 44068 12112
rect 44000 12060 44068 12078
rect 44334 12112 44400 12130
rect 44334 12078 44346 12112
rect 44380 12078 44400 12112
rect 44334 12060 44400 12078
rect 44480 12130 44520 12160
rect 44600 12130 44640 12160
rect 44720 12130 44760 12160
rect 44840 12130 44880 12160
rect 44480 12112 44546 12130
rect 44480 12078 44500 12112
rect 44534 12078 44546 12112
rect 44480 12060 44546 12078
rect 44812 12112 44880 12130
rect 44812 12078 44824 12112
rect 44858 12078 44880 12112
rect 44812 12060 44880 12078
rect 44960 12130 45000 12160
rect 45080 12130 45120 12160
rect 44960 12112 45028 12130
rect 44960 12078 44982 12112
rect 45016 12078 45028 12112
rect 44960 12060 45028 12078
rect 40710 11520 40770 11540
rect 40710 11480 40720 11520
rect 40760 11480 40770 11520
rect 40710 11460 40770 11480
rect 40880 11510 40960 11530
rect 40880 11470 40900 11510
rect 40940 11470 40960 11510
rect 41370 11510 41430 11530
rect 41370 11470 41380 11510
rect 41420 11470 41430 11510
rect 41600 11510 41680 11530
rect 41600 11470 41620 11510
rect 41660 11470 41680 11510
rect 42090 11510 42150 11530
rect 42090 11470 42100 11510
rect 42140 11470 42150 11510
rect 42320 11510 42400 11530
rect 42320 11470 42340 11510
rect 42380 11470 42400 11510
rect 42750 11510 42810 11530
rect 42750 11470 42760 11510
rect 42800 11470 42810 11510
rect 40600 11420 40640 11450
rect 40720 11420 40760 11460
rect 40840 11440 41240 11470
rect 40840 11420 40880 11440
rect 40960 11420 41000 11440
rect 41080 11420 41120 11440
rect 41200 11420 41240 11440
rect 41320 11440 41480 11470
rect 41320 11420 41360 11440
rect 41440 11420 41480 11440
rect 41560 11440 41960 11470
rect 41560 11420 41600 11440
rect 41680 11420 41720 11440
rect 41800 11420 41840 11440
rect 41920 11420 41960 11440
rect 42040 11440 42200 11470
rect 42040 11420 42080 11440
rect 42160 11420 42200 11440
rect 42280 11440 42680 11470
rect 42750 11450 42810 11470
rect 43750 11510 43810 11530
rect 43750 11470 43760 11510
rect 43800 11470 43810 11510
rect 44160 11510 44240 11530
rect 44160 11470 44180 11510
rect 44220 11470 44240 11510
rect 44410 11510 44470 11530
rect 44410 11470 44420 11510
rect 44460 11470 44470 11510
rect 44880 11510 44960 11530
rect 44880 11470 44900 11510
rect 44940 11470 44960 11510
rect 45130 11510 45190 11530
rect 45130 11470 45140 11510
rect 45180 11470 45190 11510
rect 45600 11510 45680 11530
rect 45600 11470 45620 11510
rect 45660 11470 45680 11510
rect 45790 11520 45850 11540
rect 45790 11480 45800 11520
rect 45840 11480 45850 11520
rect 43750 11450 43810 11470
rect 42280 11420 42320 11440
rect 42400 11420 42440 11440
rect 42520 11420 42560 11440
rect 42640 11420 42680 11440
rect 42760 11420 42800 11450
rect 42880 11420 42920 11450
rect 43640 11420 43680 11450
rect 43760 11420 43800 11450
rect 43880 11440 44280 11470
rect 43880 11420 43920 11440
rect 44000 11420 44040 11440
rect 44120 11420 44160 11440
rect 44240 11420 44280 11440
rect 44360 11440 44520 11470
rect 44360 11420 44400 11440
rect 44480 11420 44520 11440
rect 44600 11440 45000 11470
rect 44600 11420 44640 11440
rect 44720 11420 44760 11440
rect 44840 11420 44880 11440
rect 44960 11420 45000 11440
rect 45080 11440 45240 11470
rect 45080 11420 45120 11440
rect 45200 11420 45240 11440
rect 45320 11440 45720 11470
rect 45790 11460 45850 11480
rect 45320 11420 45360 11440
rect 45440 11420 45480 11440
rect 45560 11420 45600 11440
rect 45680 11420 45720 11440
rect 45800 11420 45840 11460
rect 45920 11420 45960 11450
rect 40600 11190 40640 11220
rect 40720 11190 40760 11220
rect 40840 11190 40880 11220
rect 40960 11190 41000 11220
rect 41080 11190 41120 11220
rect 41200 11190 41240 11220
rect 41320 11190 41360 11220
rect 41440 11190 41480 11220
rect 41560 11190 41600 11220
rect 41680 11190 41720 11220
rect 41800 11190 41840 11220
rect 41920 11190 41960 11220
rect 42040 11190 42080 11220
rect 42160 11190 42200 11220
rect 42280 11190 42320 11220
rect 42400 11190 42440 11220
rect 42520 11190 42560 11220
rect 42640 11190 42680 11220
rect 42760 11190 42800 11220
rect 42880 11190 42920 11220
rect 43640 11190 43680 11220
rect 43760 11190 43800 11220
rect 43880 11190 43920 11220
rect 44000 11190 44040 11220
rect 44120 11190 44160 11220
rect 44240 11190 44280 11220
rect 44360 11190 44400 11220
rect 44480 11190 44520 11220
rect 44600 11190 44640 11220
rect 44720 11190 44760 11220
rect 44840 11190 44880 11220
rect 44960 11190 45000 11220
rect 45080 11190 45120 11220
rect 45200 11190 45240 11220
rect 45320 11190 45360 11220
rect 45440 11190 45480 11220
rect 45560 11190 45600 11220
rect 45680 11190 45720 11220
rect 45800 11190 45840 11220
rect 45920 11190 45960 11220
rect 40530 11170 40640 11190
rect 40530 11130 40540 11170
rect 40580 11160 40640 11170
rect 42880 11170 42990 11190
rect 42880 11160 42940 11170
rect 40580 11130 40590 11160
rect 40530 11110 40590 11130
rect 42930 11130 42940 11160
rect 42980 11130 42990 11170
rect 42930 11110 42990 11130
rect 43570 11170 43680 11190
rect 43570 11130 43580 11170
rect 43620 11160 43680 11170
rect 45920 11170 46030 11190
rect 45920 11160 45980 11170
rect 43620 11130 43630 11160
rect 43570 11110 43630 11130
rect 45970 11130 45980 11160
rect 46020 11130 46030 11170
rect 45970 11110 46030 11130
rect 41900 10350 41970 10370
rect 41900 10310 41910 10350
rect 41950 10310 41970 10350
rect 41900 10290 41970 10310
rect 42070 10350 42150 10370
rect 42070 10310 42090 10350
rect 42130 10310 42150 10350
rect 42070 10290 42150 10310
rect 42250 10350 42330 10370
rect 42250 10310 42270 10350
rect 42310 10310 42330 10350
rect 42250 10290 42330 10310
rect 42430 10350 42510 10370
rect 42430 10310 42450 10350
rect 42490 10310 42510 10350
rect 42430 10290 42510 10310
rect 42610 10350 42690 10370
rect 42610 10310 42630 10350
rect 42670 10310 42690 10350
rect 42610 10290 42690 10310
rect 42790 10350 42870 10370
rect 42790 10310 42810 10350
rect 42850 10310 42870 10350
rect 42790 10290 42870 10310
rect 42970 10350 43050 10370
rect 42970 10310 42990 10350
rect 43030 10310 43050 10350
rect 42970 10290 43050 10310
rect 43150 10350 43220 10370
rect 43150 10310 43170 10350
rect 43210 10310 43220 10350
rect 43150 10290 43220 10310
rect 43340 10350 43410 10370
rect 43340 10310 43350 10350
rect 43390 10310 43410 10350
rect 43340 10290 43410 10310
rect 43510 10350 43590 10370
rect 43510 10310 43530 10350
rect 43570 10310 43590 10350
rect 43510 10290 43590 10310
rect 43690 10350 43770 10370
rect 43690 10310 43710 10350
rect 43750 10310 43770 10350
rect 43690 10290 43770 10310
rect 43870 10350 43950 10370
rect 43870 10310 43890 10350
rect 43930 10310 43950 10350
rect 43870 10290 43950 10310
rect 44050 10350 44130 10370
rect 44050 10310 44070 10350
rect 44110 10310 44130 10350
rect 44050 10290 44130 10310
rect 44230 10350 44310 10370
rect 44230 10310 44250 10350
rect 44290 10310 44310 10350
rect 44230 10290 44310 10310
rect 44410 10350 44490 10370
rect 44410 10310 44430 10350
rect 44470 10310 44490 10350
rect 44410 10290 44490 10310
rect 44590 10350 44660 10370
rect 44590 10310 44610 10350
rect 44650 10310 44660 10350
rect 44590 10300 44660 10310
rect 41700 10260 41800 10290
rect 41880 10260 41980 10290
rect 42060 10260 42160 10290
rect 42240 10260 42340 10290
rect 42420 10260 42520 10290
rect 42600 10260 42700 10290
rect 42780 10260 42880 10290
rect 42960 10260 43060 10290
rect 43140 10260 43240 10290
rect 43320 10260 43420 10290
rect 43500 10260 43600 10290
rect 43680 10260 43780 10290
rect 43860 10260 43960 10290
rect 44040 10260 44140 10290
rect 44220 10260 44320 10290
rect 44400 10260 44500 10290
rect 44580 10260 44680 10300
rect 44760 10260 44860 10290
rect 45710 10150 45790 10170
rect 45710 10110 45730 10150
rect 45770 10110 45790 10150
rect 45570 10060 45600 10090
rect 45680 10080 45820 10110
rect 45680 10060 45710 10080
rect 45790 10060 45820 10080
rect 45900 10060 45930 10090
rect 45570 9840 45600 9860
rect 45500 9810 45600 9840
rect 45680 9830 45710 9860
rect 45790 9830 45820 9860
rect 45900 9840 45930 9860
rect 45900 9810 46000 9840
rect 45500 9770 45510 9810
rect 45550 9770 45560 9810
rect 45500 9750 45560 9770
rect 45940 9770 45950 9810
rect 45990 9770 46000 9810
rect 45940 9750 46000 9770
rect 41700 9630 41800 9660
rect 41880 9630 41980 9660
rect 42060 9630 42160 9660
rect 42240 9630 42340 9660
rect 42420 9630 42520 9660
rect 42600 9630 42700 9660
rect 42780 9630 42880 9660
rect 42960 9630 43060 9660
rect 43140 9630 43240 9660
rect 43320 9630 43420 9660
rect 43500 9630 43600 9660
rect 43680 9630 43780 9660
rect 43860 9630 43960 9660
rect 44040 9630 44140 9660
rect 44220 9630 44320 9660
rect 44400 9630 44500 9660
rect 44580 9630 44680 9660
rect 44760 9630 44860 9660
rect 41620 9610 41800 9630
rect 41620 9570 41640 9610
rect 41680 9600 41800 9610
rect 44760 9610 44940 9630
rect 44760 9600 44880 9610
rect 41680 9570 41700 9600
rect 41620 9550 41700 9570
rect 44860 9570 44880 9600
rect 44920 9570 44940 9610
rect 44860 9550 44940 9570
rect 41806 9342 41864 9360
rect 41806 9308 41818 9342
rect 41852 9308 41864 9342
rect 41806 9290 41864 9308
rect 41916 9342 41974 9360
rect 41916 9308 41928 9342
rect 41962 9308 41974 9342
rect 41916 9290 41974 9308
rect 42026 9342 42084 9360
rect 42026 9308 42038 9342
rect 42072 9308 42084 9342
rect 42026 9290 42084 9308
rect 42136 9342 42194 9360
rect 42136 9308 42148 9342
rect 42182 9308 42194 9342
rect 42136 9290 42194 9308
rect 42246 9342 42304 9360
rect 42246 9308 42258 9342
rect 42292 9308 42304 9342
rect 42246 9290 42304 9308
rect 42356 9342 42414 9360
rect 42356 9308 42368 9342
rect 42402 9308 42414 9342
rect 42356 9290 42414 9308
rect 42466 9342 42524 9360
rect 42466 9308 42478 9342
rect 42512 9308 42524 9342
rect 42466 9290 42524 9308
rect 42576 9342 42634 9360
rect 42576 9308 42588 9342
rect 42622 9308 42634 9342
rect 42576 9290 42634 9308
rect 42686 9342 42744 9360
rect 42686 9308 42698 9342
rect 42732 9308 42744 9342
rect 42686 9290 42744 9308
rect 42796 9342 42854 9360
rect 42796 9308 42808 9342
rect 42842 9308 42854 9342
rect 42796 9290 42854 9308
rect 43706 9342 43764 9360
rect 43706 9308 43718 9342
rect 43752 9308 43764 9342
rect 43706 9290 43764 9308
rect 43816 9342 43874 9360
rect 43816 9308 43828 9342
rect 43862 9308 43874 9342
rect 43816 9290 43874 9308
rect 43926 9342 43984 9360
rect 43926 9308 43938 9342
rect 43972 9308 43984 9342
rect 43926 9290 43984 9308
rect 44036 9342 44094 9360
rect 44036 9308 44048 9342
rect 44082 9308 44094 9342
rect 44036 9290 44094 9308
rect 44146 9342 44204 9360
rect 44146 9308 44158 9342
rect 44192 9308 44204 9342
rect 44146 9290 44204 9308
rect 44256 9342 44314 9360
rect 44256 9308 44268 9342
rect 44302 9308 44314 9342
rect 44256 9290 44314 9308
rect 44366 9342 44424 9360
rect 44366 9308 44378 9342
rect 44412 9308 44424 9342
rect 44366 9290 44424 9308
rect 44476 9342 44534 9360
rect 44476 9308 44488 9342
rect 44522 9308 44534 9342
rect 44476 9290 44534 9308
rect 44586 9342 44644 9360
rect 44586 9308 44598 9342
rect 44632 9308 44644 9342
rect 44586 9290 44644 9308
rect 44696 9342 44754 9360
rect 44696 9308 44708 9342
rect 44742 9308 44754 9342
rect 44696 9290 44754 9308
rect 41710 9260 41740 9290
rect 41820 9260 41850 9290
rect 41930 9260 41960 9290
rect 42040 9260 42070 9290
rect 42150 9260 42180 9290
rect 42260 9260 42290 9290
rect 42370 9260 42400 9290
rect 42480 9260 42510 9290
rect 42590 9260 42620 9290
rect 42700 9260 42730 9290
rect 42810 9260 42840 9290
rect 42920 9260 42950 9290
rect 43610 9260 43640 9290
rect 43720 9260 43750 9290
rect 43830 9260 43860 9290
rect 43940 9260 43970 9290
rect 44050 9260 44080 9290
rect 44160 9260 44190 9290
rect 44270 9260 44300 9290
rect 44380 9260 44410 9290
rect 44490 9260 44520 9290
rect 44600 9260 44630 9290
rect 44710 9260 44740 9290
rect 44820 9260 44850 9290
rect 41710 9030 41740 9060
rect 41820 9030 41850 9060
rect 41930 9030 41960 9060
rect 42040 9030 42070 9060
rect 42150 9030 42180 9060
rect 42260 9030 42290 9060
rect 42370 9030 42400 9060
rect 42480 9030 42510 9060
rect 42590 9030 42620 9060
rect 42700 9030 42730 9060
rect 42810 9030 42840 9060
rect 42920 9030 42950 9060
rect 43610 9030 43640 9060
rect 43720 9030 43750 9060
rect 43830 9030 43860 9060
rect 43940 9030 43970 9060
rect 44050 9030 44080 9060
rect 44160 9030 44190 9060
rect 44270 9030 44300 9060
rect 44380 9030 44410 9060
rect 44490 9030 44520 9060
rect 44600 9030 44630 9060
rect 44710 9030 44740 9060
rect 44820 9030 44850 9060
rect 41630 9010 41740 9030
rect 41630 8970 41650 9010
rect 41690 9000 41740 9010
rect 42920 9010 43030 9030
rect 42920 9000 42970 9010
rect 41690 8970 41710 9000
rect 41630 8950 41710 8970
rect 42950 8970 42970 9000
rect 43010 8970 43030 9010
rect 42950 8950 43030 8970
rect 43530 9010 43640 9030
rect 43530 8970 43550 9010
rect 43590 9000 43640 9010
rect 44820 9010 44930 9030
rect 44820 9000 44870 9010
rect 43590 8970 43610 9000
rect 43530 8950 43610 8970
rect 44850 8970 44870 9000
rect 44910 8970 44930 9010
rect 44850 8950 44930 8970
<< polycont >>
rect 41340 13590 41380 13630
rect 41500 13590 41540 13630
rect 41660 13590 41700 13630
rect 41820 13590 41860 13630
rect 41980 13590 42020 13630
rect 42140 13590 42180 13630
rect 42300 13590 42340 13630
rect 42460 13590 42500 13630
rect 42620 13590 42660 13630
rect 42780 13590 42820 13630
rect 42940 13590 42980 13630
rect 43100 13590 43140 13630
rect 43420 13590 43460 13630
rect 43580 13590 43620 13630
rect 43740 13590 43780 13630
rect 43900 13590 43940 13630
rect 44060 13590 44100 13630
rect 44220 13590 44260 13630
rect 44380 13590 44420 13630
rect 44540 13590 44580 13630
rect 44700 13590 44740 13630
rect 44860 13590 44900 13630
rect 45020 13590 45060 13630
rect 45180 13590 45220 13630
rect 40940 12680 40980 12720
rect 41180 12680 41220 12720
rect 41420 12680 41460 12720
rect 41660 12680 41700 12720
rect 42300 12680 42340 12720
rect 42540 12680 42580 12720
rect 42780 12680 42820 12720
rect 43740 12680 43780 12720
rect 43980 12680 44020 12720
rect 44220 12680 44260 12720
rect 44860 12680 44900 12720
rect 45100 12680 45140 12720
rect 45340 12680 45380 12720
rect 45580 12680 45620 12720
rect 41443 12308 41477 12342
rect 41803 12308 41837 12342
rect 41923 12308 41957 12342
rect 42283 12308 42317 12342
rect 42403 12308 42437 12342
rect 41544 12078 41578 12112
rect 41702 12078 41736 12112
rect 42026 12078 42060 12112
rect 42180 12078 42214 12112
rect 42504 12078 42538 12112
rect 44123 12308 44157 12342
rect 44243 12308 44277 12342
rect 44603 12308 44637 12342
rect 44723 12308 44757 12342
rect 45083 12308 45117 12342
rect 44022 12078 44056 12112
rect 44346 12078 44380 12112
rect 44500 12078 44534 12112
rect 44824 12078 44858 12112
rect 44982 12078 45016 12112
rect 40720 11480 40760 11520
rect 40900 11470 40940 11510
rect 41380 11470 41420 11510
rect 41620 11470 41660 11510
rect 42100 11470 42140 11510
rect 42340 11470 42380 11510
rect 42760 11470 42800 11510
rect 43760 11470 43800 11510
rect 44180 11470 44220 11510
rect 44420 11470 44460 11510
rect 44900 11470 44940 11510
rect 45140 11470 45180 11510
rect 45620 11470 45660 11510
rect 45800 11480 45840 11520
rect 40540 11130 40580 11170
rect 42940 11130 42980 11170
rect 43580 11130 43620 11170
rect 45980 11130 46020 11170
rect 41910 10310 41950 10350
rect 42090 10310 42130 10350
rect 42270 10310 42310 10350
rect 42450 10310 42490 10350
rect 42630 10310 42670 10350
rect 42810 10310 42850 10350
rect 42990 10310 43030 10350
rect 43170 10310 43210 10350
rect 43350 10310 43390 10350
rect 43530 10310 43570 10350
rect 43710 10310 43750 10350
rect 43890 10310 43930 10350
rect 44070 10310 44110 10350
rect 44250 10310 44290 10350
rect 44430 10310 44470 10350
rect 44610 10310 44650 10350
rect 45730 10110 45770 10150
rect 45510 9770 45550 9810
rect 45950 9770 45990 9810
rect 41640 9570 41680 9610
rect 44880 9570 44920 9610
rect 41818 9308 41852 9342
rect 41928 9308 41962 9342
rect 42038 9308 42072 9342
rect 42148 9308 42182 9342
rect 42258 9308 42292 9342
rect 42368 9308 42402 9342
rect 42478 9308 42512 9342
rect 42588 9308 42622 9342
rect 42698 9308 42732 9342
rect 42808 9308 42842 9342
rect 43718 9308 43752 9342
rect 43828 9308 43862 9342
rect 43938 9308 43972 9342
rect 44048 9308 44082 9342
rect 44158 9308 44192 9342
rect 44268 9308 44302 9342
rect 44378 9308 44412 9342
rect 44488 9308 44522 9342
rect 44598 9308 44632 9342
rect 44708 9308 44742 9342
rect 41650 8970 41690 9010
rect 42970 8970 43010 9010
rect 43550 8970 43590 9010
rect 44870 8970 44910 9010
<< xpolycontact >>
rect 38760 18018 38898 18450
rect 38760 16632 38898 17064
rect 39574 18024 39644 18456
rect 39574 15062 39644 15494
rect 40686 18026 40756 18458
rect 40354 16286 40424 16718
rect 45674 18026 45744 18458
rect 46006 16286 46076 16718
rect 46784 18024 46854 18456
rect 46784 15952 46854 16384
rect 47540 18018 47678 18450
rect 47540 16632 47678 17064
rect 41542 14344 41974 14414
rect 44582 14344 45014 14414
<< ppolyres >>
rect 38760 17064 38898 18018
rect 46784 16384 46854 18024
rect 47540 17064 47678 18018
rect 41974 14344 44582 14414
<< xpolyres >>
rect 39574 15494 39644 18024
rect 40354 17852 40590 17922
rect 40354 16718 40424 17852
rect 40520 16892 40590 17852
rect 40686 16892 40756 18026
rect 40520 16822 40756 16892
rect 45674 16892 45744 18026
rect 45840 17852 46076 17922
rect 45840 16892 45910 17852
rect 45674 16822 45910 16892
rect 46006 16718 46076 17852
<< locali >>
rect 43240 19070 43320 19090
rect 43240 19030 43260 19070
rect 43300 19030 43320 19070
rect 43240 18990 43320 19030
rect 43240 18950 43260 18990
rect 43300 18950 43320 18990
rect 43240 18910 43320 18950
rect 43240 18870 43260 18910
rect 43300 18870 43320 18910
rect 42560 18784 42640 18790
rect 43240 18784 43320 18870
rect 43920 18784 44000 18790
rect 41276 18752 45284 18784
rect 41276 18718 41410 18752
rect 41444 18718 41500 18752
rect 41534 18718 41590 18752
rect 41624 18718 41680 18752
rect 41714 18718 41770 18752
rect 41804 18718 41860 18752
rect 41894 18718 41950 18752
rect 41984 18718 42040 18752
rect 42074 18718 42130 18752
rect 42164 18718 42220 18752
rect 42254 18718 42310 18752
rect 42344 18718 42400 18752
rect 42434 18718 42770 18752
rect 42804 18718 42860 18752
rect 42894 18718 42950 18752
rect 42984 18718 43040 18752
rect 43074 18718 43130 18752
rect 43164 18718 43220 18752
rect 43254 18718 43310 18752
rect 43344 18718 43400 18752
rect 43434 18718 43490 18752
rect 43524 18718 43580 18752
rect 43614 18718 43670 18752
rect 43704 18718 43760 18752
rect 43794 18718 44130 18752
rect 44164 18718 44220 18752
rect 44254 18718 44310 18752
rect 44344 18718 44400 18752
rect 44434 18718 44490 18752
rect 44524 18718 44580 18752
rect 44614 18718 44670 18752
rect 44704 18718 44760 18752
rect 44794 18718 44850 18752
rect 44884 18718 44940 18752
rect 44974 18718 45030 18752
rect 45064 18718 45120 18752
rect 45154 18718 45284 18752
rect 41276 18685 45284 18718
rect 41276 18668 41375 18685
rect 41276 18634 41309 18668
rect 41343 18634 41375 18668
rect 38790 18590 38870 18610
rect 39570 18600 39650 18620
rect 39570 18595 39590 18600
rect 39630 18595 39650 18600
rect 40680 18610 40760 18630
rect 40680 18597 40700 18610
rect 40740 18597 40760 18610
rect 38790 18589 38810 18590
rect 38850 18589 38870 18590
rect 38603 18555 38699 18589
rect 38959 18555 39055 18589
rect 38603 18493 38637 18555
rect 38790 18550 38810 18555
rect 38850 18550 38870 18555
rect 38790 18530 38870 18550
rect 39021 18493 39055 18555
rect 38603 16527 38637 16589
rect 39021 16527 39055 16589
rect 38603 16493 38699 16527
rect 38959 16493 39055 16527
rect 39383 18561 39479 18595
rect 39739 18561 39835 18595
rect 39383 18499 39417 18561
rect 39570 18560 39590 18561
rect 39630 18560 39650 18561
rect 39570 18540 39650 18560
rect 39801 18499 39835 18561
rect 39383 14957 39417 15019
rect 40163 18563 40259 18597
rect 40851 18563 40947 18597
rect 40163 18501 40197 18563
rect 40680 18550 40760 18563
rect 40913 18501 40947 18563
rect 40163 16181 40197 16243
rect 41276 18578 41375 18634
rect 42465 18668 42735 18685
rect 42465 18634 42496 18668
rect 42530 18634 42669 18668
rect 42703 18634 42735 18668
rect 41276 18544 41309 18578
rect 41343 18544 41375 18578
rect 41276 18488 41375 18544
rect 41276 18454 41309 18488
rect 41343 18454 41375 18488
rect 41276 18398 41375 18454
rect 41276 18364 41309 18398
rect 41343 18364 41375 18398
rect 41276 18308 41375 18364
rect 41276 18274 41309 18308
rect 41343 18274 41375 18308
rect 41276 18218 41375 18274
rect 41276 18184 41309 18218
rect 41343 18184 41375 18218
rect 41276 18128 41375 18184
rect 41276 18094 41309 18128
rect 41343 18094 41375 18128
rect 41276 18038 41375 18094
rect 41276 18004 41309 18038
rect 41343 18004 41375 18038
rect 41276 17948 41375 18004
rect 41276 17914 41309 17948
rect 41343 17914 41375 17948
rect 41276 17858 41375 17914
rect 41276 17824 41309 17858
rect 41343 17824 41375 17858
rect 41276 17768 41375 17824
rect 41276 17740 41309 17768
rect 41270 17734 41309 17740
rect 41343 17740 41375 17768
rect 41439 18602 42401 18621
rect 41439 18568 41550 18602
rect 41584 18568 41640 18602
rect 41674 18568 41730 18602
rect 41764 18568 41820 18602
rect 41854 18568 41910 18602
rect 41944 18568 42000 18602
rect 42034 18568 42090 18602
rect 42124 18568 42180 18602
rect 42214 18568 42270 18602
rect 42304 18568 42401 18602
rect 41439 18549 42401 18568
rect 41439 18508 41511 18549
rect 41439 18474 41458 18508
rect 41492 18474 41511 18508
rect 42329 18489 42401 18549
rect 41439 18418 41511 18474
rect 41439 18384 41458 18418
rect 41492 18384 41511 18418
rect 41439 18328 41511 18384
rect 41439 18294 41458 18328
rect 41492 18294 41511 18328
rect 41439 18238 41511 18294
rect 41439 18204 41458 18238
rect 41492 18204 41511 18238
rect 41439 18148 41511 18204
rect 41439 18114 41458 18148
rect 41492 18114 41511 18148
rect 41439 18058 41511 18114
rect 41439 18024 41458 18058
rect 41492 18024 41511 18058
rect 41439 17968 41511 18024
rect 41439 17934 41458 17968
rect 41492 17934 41511 17968
rect 41439 17878 41511 17934
rect 41439 17844 41458 17878
rect 41492 17844 41511 17878
rect 41439 17788 41511 17844
rect 41573 18426 42267 18487
rect 41573 18392 41632 18426
rect 41666 18414 41722 18426
rect 41694 18392 41722 18414
rect 41756 18414 41812 18426
rect 41756 18392 41760 18414
rect 41573 18380 41660 18392
rect 41694 18380 41760 18392
rect 41794 18392 41812 18414
rect 41846 18414 41902 18426
rect 41846 18392 41860 18414
rect 41794 18380 41860 18392
rect 41894 18392 41902 18414
rect 41936 18414 41992 18426
rect 42026 18414 42082 18426
rect 42116 18414 42172 18426
rect 41936 18392 41960 18414
rect 42026 18392 42060 18414
rect 42116 18392 42160 18414
rect 42206 18392 42267 18426
rect 41894 18380 41960 18392
rect 41994 18380 42060 18392
rect 42094 18380 42160 18392
rect 42194 18380 42267 18392
rect 41573 18336 42267 18380
rect 41573 18302 41632 18336
rect 41666 18314 41722 18336
rect 41694 18302 41722 18314
rect 41756 18314 41812 18336
rect 41756 18302 41760 18314
rect 41573 18280 41660 18302
rect 41694 18280 41760 18302
rect 41794 18302 41812 18314
rect 41846 18314 41902 18336
rect 41846 18302 41860 18314
rect 41794 18280 41860 18302
rect 41894 18302 41902 18314
rect 41936 18314 41992 18336
rect 42026 18314 42082 18336
rect 42116 18314 42172 18336
rect 41936 18302 41960 18314
rect 42026 18302 42060 18314
rect 42116 18302 42160 18314
rect 42206 18302 42267 18336
rect 41894 18280 41960 18302
rect 41994 18280 42060 18302
rect 42094 18280 42160 18302
rect 42194 18280 42267 18302
rect 41573 18246 42267 18280
rect 41573 18212 41632 18246
rect 41666 18214 41722 18246
rect 41694 18212 41722 18214
rect 41756 18214 41812 18246
rect 41756 18212 41760 18214
rect 41573 18180 41660 18212
rect 41694 18180 41760 18212
rect 41794 18212 41812 18214
rect 41846 18214 41902 18246
rect 41846 18212 41860 18214
rect 41794 18180 41860 18212
rect 41894 18212 41902 18214
rect 41936 18214 41992 18246
rect 42026 18214 42082 18246
rect 42116 18214 42172 18246
rect 41936 18212 41960 18214
rect 42026 18212 42060 18214
rect 42116 18212 42160 18214
rect 42206 18212 42267 18246
rect 41894 18180 41960 18212
rect 41994 18180 42060 18212
rect 42094 18180 42160 18212
rect 42194 18180 42267 18212
rect 41573 18156 42267 18180
rect 41573 18122 41632 18156
rect 41666 18122 41722 18156
rect 41756 18122 41812 18156
rect 41846 18122 41902 18156
rect 41936 18122 41992 18156
rect 42026 18122 42082 18156
rect 42116 18122 42172 18156
rect 42206 18122 42267 18156
rect 41573 18114 42267 18122
rect 41573 18080 41660 18114
rect 41694 18080 41760 18114
rect 41794 18080 41860 18114
rect 41894 18080 41960 18114
rect 41994 18080 42060 18114
rect 42094 18080 42160 18114
rect 42194 18080 42267 18114
rect 41573 18066 42267 18080
rect 41573 18032 41632 18066
rect 41666 18032 41722 18066
rect 41756 18032 41812 18066
rect 41846 18032 41902 18066
rect 41936 18032 41992 18066
rect 42026 18032 42082 18066
rect 42116 18032 42172 18066
rect 42206 18032 42267 18066
rect 41573 18014 42267 18032
rect 41573 17980 41660 18014
rect 41694 17980 41760 18014
rect 41794 17980 41860 18014
rect 41894 17980 41960 18014
rect 41994 17980 42060 18014
rect 42094 17980 42160 18014
rect 42194 17980 42267 18014
rect 41573 17976 42267 17980
rect 41573 17942 41632 17976
rect 41666 17942 41722 17976
rect 41756 17942 41812 17976
rect 41846 17942 41902 17976
rect 41936 17942 41992 17976
rect 42026 17942 42082 17976
rect 42116 17942 42172 17976
rect 42206 17942 42267 17976
rect 41573 17914 42267 17942
rect 41573 17886 41660 17914
rect 41694 17886 41760 17914
rect 41573 17852 41632 17886
rect 41694 17880 41722 17886
rect 41666 17852 41722 17880
rect 41756 17880 41760 17886
rect 41794 17886 41860 17914
rect 41794 17880 41812 17886
rect 41756 17852 41812 17880
rect 41846 17880 41860 17886
rect 41894 17886 41960 17914
rect 41994 17886 42060 17914
rect 42094 17886 42160 17914
rect 42194 17886 42267 17914
rect 41894 17880 41902 17886
rect 41846 17852 41902 17880
rect 41936 17880 41960 17886
rect 42026 17880 42060 17886
rect 42116 17880 42160 17886
rect 41936 17852 41992 17880
rect 42026 17852 42082 17880
rect 42116 17852 42172 17880
rect 42206 17852 42267 17886
rect 41573 17793 42267 17852
rect 42329 18455 42348 18489
rect 42382 18455 42401 18489
rect 42329 18399 42401 18455
rect 42329 18365 42348 18399
rect 42382 18365 42401 18399
rect 42329 18309 42401 18365
rect 42329 18275 42348 18309
rect 42382 18275 42401 18309
rect 42329 18219 42401 18275
rect 42329 18185 42348 18219
rect 42382 18185 42401 18219
rect 42329 18129 42401 18185
rect 42329 18095 42348 18129
rect 42382 18095 42401 18129
rect 42329 18039 42401 18095
rect 42329 18005 42348 18039
rect 42382 18005 42401 18039
rect 42329 17949 42401 18005
rect 42329 17915 42348 17949
rect 42382 17915 42401 17949
rect 42329 17859 42401 17915
rect 42329 17825 42348 17859
rect 42382 17825 42401 17859
rect 41439 17754 41458 17788
rect 41492 17754 41511 17788
rect 41439 17740 41511 17754
rect 42329 17769 42401 17825
rect 42329 17740 42348 17769
rect 41343 17735 42348 17740
rect 42382 17740 42401 17769
rect 42465 18578 42735 18634
rect 43825 18668 44095 18685
rect 43825 18634 43856 18668
rect 43890 18634 44029 18668
rect 44063 18634 44095 18668
rect 42465 18544 42496 18578
rect 42530 18544 42669 18578
rect 42703 18544 42735 18578
rect 42465 18488 42735 18544
rect 42465 18454 42496 18488
rect 42530 18454 42669 18488
rect 42703 18454 42735 18488
rect 42465 18398 42735 18454
rect 42465 18364 42496 18398
rect 42530 18364 42669 18398
rect 42703 18364 42735 18398
rect 42465 18308 42735 18364
rect 42465 18274 42496 18308
rect 42530 18274 42669 18308
rect 42703 18274 42735 18308
rect 42465 18218 42735 18274
rect 42465 18184 42496 18218
rect 42530 18184 42669 18218
rect 42703 18184 42735 18218
rect 42465 18128 42735 18184
rect 42465 18094 42496 18128
rect 42530 18094 42669 18128
rect 42703 18094 42735 18128
rect 42465 18038 42735 18094
rect 42465 18004 42496 18038
rect 42530 18004 42669 18038
rect 42703 18004 42735 18038
rect 42465 17948 42735 18004
rect 42465 17914 42496 17948
rect 42530 17914 42669 17948
rect 42703 17914 42735 17948
rect 42465 17858 42735 17914
rect 42465 17824 42496 17858
rect 42530 17824 42669 17858
rect 42703 17824 42735 17858
rect 42465 17768 42735 17824
rect 42465 17740 42496 17768
rect 42382 17735 42496 17740
rect 41343 17734 42496 17735
rect 42530 17734 42669 17768
rect 42703 17740 42735 17768
rect 42799 18602 43761 18621
rect 42799 18568 42910 18602
rect 42944 18568 43000 18602
rect 43034 18568 43090 18602
rect 43124 18568 43180 18602
rect 43214 18568 43270 18602
rect 43304 18568 43360 18602
rect 43394 18568 43450 18602
rect 43484 18568 43540 18602
rect 43574 18568 43630 18602
rect 43664 18568 43761 18602
rect 42799 18549 43761 18568
rect 42799 18508 42871 18549
rect 42799 18474 42818 18508
rect 42852 18474 42871 18508
rect 43689 18489 43761 18549
rect 42799 18418 42871 18474
rect 42799 18384 42818 18418
rect 42852 18384 42871 18418
rect 42799 18328 42871 18384
rect 42799 18294 42818 18328
rect 42852 18294 42871 18328
rect 42799 18238 42871 18294
rect 42799 18204 42818 18238
rect 42852 18204 42871 18238
rect 42799 18148 42871 18204
rect 42799 18114 42818 18148
rect 42852 18114 42871 18148
rect 42799 18058 42871 18114
rect 42799 18024 42818 18058
rect 42852 18024 42871 18058
rect 42799 17968 42871 18024
rect 42799 17934 42818 17968
rect 42852 17934 42871 17968
rect 42799 17878 42871 17934
rect 42799 17844 42818 17878
rect 42852 17844 42871 17878
rect 42799 17788 42871 17844
rect 42933 18426 43627 18487
rect 42933 18392 42992 18426
rect 43026 18414 43082 18426
rect 43054 18392 43082 18414
rect 43116 18414 43172 18426
rect 43116 18392 43120 18414
rect 42933 18380 43020 18392
rect 43054 18380 43120 18392
rect 43154 18392 43172 18414
rect 43206 18414 43262 18426
rect 43206 18392 43220 18414
rect 43154 18380 43220 18392
rect 43254 18392 43262 18414
rect 43296 18414 43352 18426
rect 43386 18414 43442 18426
rect 43476 18414 43532 18426
rect 43296 18392 43320 18414
rect 43386 18392 43420 18414
rect 43476 18392 43520 18414
rect 43566 18392 43627 18426
rect 43254 18380 43320 18392
rect 43354 18380 43420 18392
rect 43454 18380 43520 18392
rect 43554 18380 43627 18392
rect 42933 18336 43627 18380
rect 42933 18302 42992 18336
rect 43026 18314 43082 18336
rect 43054 18302 43082 18314
rect 43116 18314 43172 18336
rect 43116 18302 43120 18314
rect 42933 18280 43020 18302
rect 43054 18280 43120 18302
rect 43154 18302 43172 18314
rect 43206 18314 43262 18336
rect 43206 18302 43220 18314
rect 43154 18280 43220 18302
rect 43254 18302 43262 18314
rect 43296 18314 43352 18336
rect 43386 18314 43442 18336
rect 43476 18314 43532 18336
rect 43296 18302 43320 18314
rect 43386 18302 43420 18314
rect 43476 18302 43520 18314
rect 43566 18302 43627 18336
rect 43254 18280 43320 18302
rect 43354 18280 43420 18302
rect 43454 18280 43520 18302
rect 43554 18280 43627 18302
rect 42933 18246 43627 18280
rect 42933 18212 42992 18246
rect 43026 18214 43082 18246
rect 43054 18212 43082 18214
rect 43116 18214 43172 18246
rect 43116 18212 43120 18214
rect 42933 18180 43020 18212
rect 43054 18180 43120 18212
rect 43154 18212 43172 18214
rect 43206 18214 43262 18246
rect 43206 18212 43220 18214
rect 43154 18180 43220 18212
rect 43254 18212 43262 18214
rect 43296 18214 43352 18246
rect 43386 18214 43442 18246
rect 43476 18214 43532 18246
rect 43296 18212 43320 18214
rect 43386 18212 43420 18214
rect 43476 18212 43520 18214
rect 43566 18212 43627 18246
rect 43254 18180 43320 18212
rect 43354 18180 43420 18212
rect 43454 18180 43520 18212
rect 43554 18180 43627 18212
rect 42933 18156 43627 18180
rect 42933 18122 42992 18156
rect 43026 18122 43082 18156
rect 43116 18122 43172 18156
rect 43206 18122 43262 18156
rect 43296 18122 43352 18156
rect 43386 18122 43442 18156
rect 43476 18122 43532 18156
rect 43566 18122 43627 18156
rect 42933 18114 43627 18122
rect 42933 18080 43020 18114
rect 43054 18080 43120 18114
rect 43154 18080 43220 18114
rect 43254 18080 43320 18114
rect 43354 18080 43420 18114
rect 43454 18080 43520 18114
rect 43554 18080 43627 18114
rect 42933 18066 43627 18080
rect 42933 18032 42992 18066
rect 43026 18032 43082 18066
rect 43116 18032 43172 18066
rect 43206 18032 43262 18066
rect 43296 18032 43352 18066
rect 43386 18032 43442 18066
rect 43476 18032 43532 18066
rect 43566 18032 43627 18066
rect 42933 18014 43627 18032
rect 42933 17980 43020 18014
rect 43054 17980 43120 18014
rect 43154 17980 43220 18014
rect 43254 17980 43320 18014
rect 43354 17980 43420 18014
rect 43454 17980 43520 18014
rect 43554 17980 43627 18014
rect 42933 17976 43627 17980
rect 42933 17942 42992 17976
rect 43026 17942 43082 17976
rect 43116 17942 43172 17976
rect 43206 17942 43262 17976
rect 43296 17942 43352 17976
rect 43386 17942 43442 17976
rect 43476 17942 43532 17976
rect 43566 17942 43627 17976
rect 42933 17914 43627 17942
rect 42933 17886 43020 17914
rect 43054 17886 43120 17914
rect 42933 17852 42992 17886
rect 43054 17880 43082 17886
rect 43026 17852 43082 17880
rect 43116 17880 43120 17886
rect 43154 17886 43220 17914
rect 43154 17880 43172 17886
rect 43116 17852 43172 17880
rect 43206 17880 43220 17886
rect 43254 17886 43320 17914
rect 43354 17886 43420 17914
rect 43454 17886 43520 17914
rect 43554 17886 43627 17914
rect 43254 17880 43262 17886
rect 43206 17852 43262 17880
rect 43296 17880 43320 17886
rect 43386 17880 43420 17886
rect 43476 17880 43520 17886
rect 43296 17852 43352 17880
rect 43386 17852 43442 17880
rect 43476 17852 43532 17880
rect 43566 17852 43627 17886
rect 42933 17793 43627 17852
rect 43689 18455 43708 18489
rect 43742 18455 43761 18489
rect 43689 18399 43761 18455
rect 43689 18365 43708 18399
rect 43742 18365 43761 18399
rect 43689 18309 43761 18365
rect 43689 18275 43708 18309
rect 43742 18275 43761 18309
rect 43689 18219 43761 18275
rect 43689 18185 43708 18219
rect 43742 18185 43761 18219
rect 43689 18129 43761 18185
rect 43689 18095 43708 18129
rect 43742 18095 43761 18129
rect 43689 18039 43761 18095
rect 43689 18005 43708 18039
rect 43742 18005 43761 18039
rect 43689 17949 43761 18005
rect 43689 17915 43708 17949
rect 43742 17915 43761 17949
rect 43689 17859 43761 17915
rect 43689 17825 43708 17859
rect 43742 17825 43761 17859
rect 42799 17754 42818 17788
rect 42852 17754 42871 17788
rect 42799 17740 42871 17754
rect 43689 17769 43761 17825
rect 43689 17740 43708 17769
rect 42703 17735 43708 17740
rect 43742 17740 43761 17769
rect 43825 18578 44095 18634
rect 45185 18668 45284 18685
rect 45185 18634 45216 18668
rect 45250 18634 45284 18668
rect 43825 18544 43856 18578
rect 43890 18544 44029 18578
rect 44063 18544 44095 18578
rect 43825 18488 44095 18544
rect 43825 18454 43856 18488
rect 43890 18454 44029 18488
rect 44063 18454 44095 18488
rect 43825 18398 44095 18454
rect 43825 18364 43856 18398
rect 43890 18364 44029 18398
rect 44063 18364 44095 18398
rect 43825 18308 44095 18364
rect 43825 18274 43856 18308
rect 43890 18274 44029 18308
rect 44063 18274 44095 18308
rect 43825 18218 44095 18274
rect 43825 18184 43856 18218
rect 43890 18184 44029 18218
rect 44063 18184 44095 18218
rect 43825 18128 44095 18184
rect 43825 18094 43856 18128
rect 43890 18094 44029 18128
rect 44063 18094 44095 18128
rect 43825 18038 44095 18094
rect 43825 18004 43856 18038
rect 43890 18004 44029 18038
rect 44063 18004 44095 18038
rect 43825 17948 44095 18004
rect 43825 17914 43856 17948
rect 43890 17914 44029 17948
rect 44063 17914 44095 17948
rect 43825 17858 44095 17914
rect 43825 17824 43856 17858
rect 43890 17824 44029 17858
rect 44063 17824 44095 17858
rect 43825 17768 44095 17824
rect 43825 17740 43856 17768
rect 43742 17735 43856 17740
rect 42703 17734 43856 17735
rect 43890 17734 44029 17768
rect 44063 17740 44095 17768
rect 44159 18602 45121 18621
rect 44159 18568 44270 18602
rect 44304 18568 44360 18602
rect 44394 18568 44450 18602
rect 44484 18568 44540 18602
rect 44574 18568 44630 18602
rect 44664 18568 44720 18602
rect 44754 18568 44810 18602
rect 44844 18568 44900 18602
rect 44934 18568 44990 18602
rect 45024 18568 45121 18602
rect 44159 18549 45121 18568
rect 44159 18508 44231 18549
rect 44159 18474 44178 18508
rect 44212 18474 44231 18508
rect 45049 18489 45121 18549
rect 44159 18418 44231 18474
rect 44159 18384 44178 18418
rect 44212 18384 44231 18418
rect 44159 18328 44231 18384
rect 44159 18294 44178 18328
rect 44212 18294 44231 18328
rect 44159 18238 44231 18294
rect 44159 18204 44178 18238
rect 44212 18204 44231 18238
rect 44159 18148 44231 18204
rect 44159 18114 44178 18148
rect 44212 18114 44231 18148
rect 44159 18058 44231 18114
rect 44159 18024 44178 18058
rect 44212 18024 44231 18058
rect 44159 17968 44231 18024
rect 44159 17934 44178 17968
rect 44212 17934 44231 17968
rect 44159 17878 44231 17934
rect 44159 17844 44178 17878
rect 44212 17844 44231 17878
rect 44159 17788 44231 17844
rect 44293 18426 44987 18487
rect 44293 18392 44352 18426
rect 44386 18414 44442 18426
rect 44414 18392 44442 18414
rect 44476 18414 44532 18426
rect 44476 18392 44480 18414
rect 44293 18380 44380 18392
rect 44414 18380 44480 18392
rect 44514 18392 44532 18414
rect 44566 18414 44622 18426
rect 44566 18392 44580 18414
rect 44514 18380 44580 18392
rect 44614 18392 44622 18414
rect 44656 18414 44712 18426
rect 44746 18414 44802 18426
rect 44836 18414 44892 18426
rect 44656 18392 44680 18414
rect 44746 18392 44780 18414
rect 44836 18392 44880 18414
rect 44926 18392 44987 18426
rect 44614 18380 44680 18392
rect 44714 18380 44780 18392
rect 44814 18380 44880 18392
rect 44914 18380 44987 18392
rect 44293 18336 44987 18380
rect 44293 18302 44352 18336
rect 44386 18314 44442 18336
rect 44414 18302 44442 18314
rect 44476 18314 44532 18336
rect 44476 18302 44480 18314
rect 44293 18280 44380 18302
rect 44414 18280 44480 18302
rect 44514 18302 44532 18314
rect 44566 18314 44622 18336
rect 44566 18302 44580 18314
rect 44514 18280 44580 18302
rect 44614 18302 44622 18314
rect 44656 18314 44712 18336
rect 44746 18314 44802 18336
rect 44836 18314 44892 18336
rect 44656 18302 44680 18314
rect 44746 18302 44780 18314
rect 44836 18302 44880 18314
rect 44926 18302 44987 18336
rect 44614 18280 44680 18302
rect 44714 18280 44780 18302
rect 44814 18280 44880 18302
rect 44914 18280 44987 18302
rect 44293 18246 44987 18280
rect 44293 18212 44352 18246
rect 44386 18214 44442 18246
rect 44414 18212 44442 18214
rect 44476 18214 44532 18246
rect 44476 18212 44480 18214
rect 44293 18180 44380 18212
rect 44414 18180 44480 18212
rect 44514 18212 44532 18214
rect 44566 18214 44622 18246
rect 44566 18212 44580 18214
rect 44514 18180 44580 18212
rect 44614 18212 44622 18214
rect 44656 18214 44712 18246
rect 44746 18214 44802 18246
rect 44836 18214 44892 18246
rect 44656 18212 44680 18214
rect 44746 18212 44780 18214
rect 44836 18212 44880 18214
rect 44926 18212 44987 18246
rect 44614 18180 44680 18212
rect 44714 18180 44780 18212
rect 44814 18180 44880 18212
rect 44914 18180 44987 18212
rect 44293 18156 44987 18180
rect 44293 18122 44352 18156
rect 44386 18122 44442 18156
rect 44476 18122 44532 18156
rect 44566 18122 44622 18156
rect 44656 18122 44712 18156
rect 44746 18122 44802 18156
rect 44836 18122 44892 18156
rect 44926 18122 44987 18156
rect 44293 18114 44987 18122
rect 44293 18080 44380 18114
rect 44414 18080 44480 18114
rect 44514 18080 44580 18114
rect 44614 18080 44680 18114
rect 44714 18080 44780 18114
rect 44814 18080 44880 18114
rect 44914 18080 44987 18114
rect 44293 18066 44987 18080
rect 44293 18032 44352 18066
rect 44386 18032 44442 18066
rect 44476 18032 44532 18066
rect 44566 18032 44622 18066
rect 44656 18032 44712 18066
rect 44746 18032 44802 18066
rect 44836 18032 44892 18066
rect 44926 18032 44987 18066
rect 44293 18014 44987 18032
rect 44293 17980 44380 18014
rect 44414 17980 44480 18014
rect 44514 17980 44580 18014
rect 44614 17980 44680 18014
rect 44714 17980 44780 18014
rect 44814 17980 44880 18014
rect 44914 17980 44987 18014
rect 44293 17976 44987 17980
rect 44293 17942 44352 17976
rect 44386 17942 44442 17976
rect 44476 17942 44532 17976
rect 44566 17942 44622 17976
rect 44656 17942 44712 17976
rect 44746 17942 44802 17976
rect 44836 17942 44892 17976
rect 44926 17942 44987 17976
rect 44293 17914 44987 17942
rect 44293 17886 44380 17914
rect 44414 17886 44480 17914
rect 44293 17852 44352 17886
rect 44414 17880 44442 17886
rect 44386 17852 44442 17880
rect 44476 17880 44480 17886
rect 44514 17886 44580 17914
rect 44514 17880 44532 17886
rect 44476 17852 44532 17880
rect 44566 17880 44580 17886
rect 44614 17886 44680 17914
rect 44714 17886 44780 17914
rect 44814 17886 44880 17914
rect 44914 17886 44987 17914
rect 44614 17880 44622 17886
rect 44566 17852 44622 17880
rect 44656 17880 44680 17886
rect 44746 17880 44780 17886
rect 44836 17880 44880 17886
rect 44656 17852 44712 17880
rect 44746 17852 44802 17880
rect 44836 17852 44892 17880
rect 44926 17852 44987 17886
rect 44293 17793 44987 17852
rect 45049 18455 45068 18489
rect 45102 18455 45121 18489
rect 45049 18399 45121 18455
rect 45049 18365 45068 18399
rect 45102 18365 45121 18399
rect 45049 18309 45121 18365
rect 45049 18275 45068 18309
rect 45102 18275 45121 18309
rect 45049 18219 45121 18275
rect 45049 18185 45068 18219
rect 45102 18185 45121 18219
rect 45049 18129 45121 18185
rect 45049 18095 45068 18129
rect 45102 18095 45121 18129
rect 45049 18039 45121 18095
rect 45049 18005 45068 18039
rect 45102 18005 45121 18039
rect 45049 17949 45121 18005
rect 45049 17915 45068 17949
rect 45102 17915 45121 17949
rect 45049 17859 45121 17915
rect 45049 17825 45068 17859
rect 45102 17825 45121 17859
rect 44159 17754 44178 17788
rect 44212 17754 44231 17788
rect 44159 17740 44231 17754
rect 45049 17769 45121 17825
rect 45049 17740 45068 17769
rect 44063 17735 45068 17740
rect 45102 17740 45121 17769
rect 45185 18578 45284 18634
rect 45670 18610 45750 18630
rect 45670 18597 45690 18610
rect 45730 18597 45750 18610
rect 46780 18610 46860 18630
rect 45185 18544 45216 18578
rect 45250 18544 45284 18578
rect 45185 18488 45284 18544
rect 45185 18454 45216 18488
rect 45250 18454 45284 18488
rect 45185 18398 45284 18454
rect 45185 18364 45216 18398
rect 45250 18364 45284 18398
rect 45185 18308 45284 18364
rect 45185 18274 45216 18308
rect 45250 18274 45284 18308
rect 45185 18218 45284 18274
rect 45185 18184 45216 18218
rect 45250 18184 45284 18218
rect 45185 18128 45284 18184
rect 45185 18094 45216 18128
rect 45250 18094 45284 18128
rect 45185 18038 45284 18094
rect 45185 18004 45216 18038
rect 45250 18004 45284 18038
rect 45185 17948 45284 18004
rect 45185 17914 45216 17948
rect 45250 17914 45284 17948
rect 45185 17858 45284 17914
rect 45185 17824 45216 17858
rect 45250 17824 45284 17858
rect 45185 17768 45284 17824
rect 45185 17740 45216 17768
rect 45102 17735 45216 17740
rect 44063 17734 45216 17735
rect 45250 17740 45284 17768
rect 45483 18563 45579 18597
rect 46171 18563 46267 18597
rect 46780 18595 46800 18610
rect 46840 18595 46860 18610
rect 45483 18501 45517 18563
rect 45670 18550 45750 18563
rect 45250 17734 45290 17740
rect 41270 17712 45290 17734
rect 41270 17678 41516 17712
rect 41550 17678 41606 17712
rect 41640 17678 41696 17712
rect 41730 17678 41786 17712
rect 41820 17678 41876 17712
rect 41910 17678 41966 17712
rect 42000 17678 42056 17712
rect 42090 17678 42146 17712
rect 42180 17678 42236 17712
rect 42270 17678 42876 17712
rect 42910 17678 42966 17712
rect 43000 17678 43056 17712
rect 43090 17678 43146 17712
rect 43180 17678 43236 17712
rect 43270 17678 43326 17712
rect 43360 17678 43416 17712
rect 43450 17678 43506 17712
rect 43540 17678 43596 17712
rect 43630 17678 44236 17712
rect 44270 17678 44326 17712
rect 44360 17678 44416 17712
rect 44450 17678 44506 17712
rect 44540 17678 44596 17712
rect 44630 17678 44686 17712
rect 44720 17678 44776 17712
rect 44810 17678 44866 17712
rect 44900 17678 44956 17712
rect 44990 17678 45290 17712
rect 41270 17644 41309 17678
rect 41343 17644 42496 17678
rect 42530 17644 42669 17678
rect 42703 17644 43856 17678
rect 43890 17644 44029 17678
rect 44063 17644 45216 17678
rect 45250 17644 45290 17678
rect 41270 17588 45290 17644
rect 41270 17554 41309 17588
rect 41343 17565 42496 17588
rect 41343 17554 41410 17565
rect 41270 17531 41410 17554
rect 41444 17531 41500 17565
rect 41534 17531 41590 17565
rect 41624 17531 41680 17565
rect 41714 17531 41770 17565
rect 41804 17531 41860 17565
rect 41894 17531 41950 17565
rect 41984 17531 42040 17565
rect 42074 17531 42130 17565
rect 42164 17531 42220 17565
rect 42254 17531 42310 17565
rect 42344 17531 42400 17565
rect 42434 17554 42496 17565
rect 42530 17554 42669 17588
rect 42703 17565 43856 17588
rect 42703 17554 42770 17565
rect 42434 17531 42770 17554
rect 42804 17531 42860 17565
rect 42894 17531 42950 17565
rect 42984 17531 43040 17565
rect 43074 17531 43130 17565
rect 43164 17531 43220 17565
rect 43254 17531 43310 17565
rect 43344 17531 43400 17565
rect 43434 17531 43490 17565
rect 43524 17531 43580 17565
rect 43614 17531 43670 17565
rect 43704 17531 43760 17565
rect 43794 17554 43856 17565
rect 43890 17554 44029 17588
rect 44063 17565 45216 17588
rect 44063 17554 44130 17565
rect 43794 17531 44130 17554
rect 44164 17531 44220 17565
rect 44254 17531 44310 17565
rect 44344 17531 44400 17565
rect 44434 17531 44490 17565
rect 44524 17531 44580 17565
rect 44614 17531 44670 17565
rect 44704 17531 44760 17565
rect 44794 17531 44850 17565
rect 44884 17531 44940 17565
rect 44974 17531 45030 17565
rect 45064 17531 45120 17565
rect 45154 17554 45216 17565
rect 45250 17554 45290 17588
rect 45154 17531 45290 17554
rect 41270 17490 45290 17531
rect 42560 17424 42640 17490
rect 43920 17424 44000 17490
rect 41276 17392 45284 17424
rect 41276 17358 41410 17392
rect 41444 17358 41500 17392
rect 41534 17358 41590 17392
rect 41624 17358 41680 17392
rect 41714 17358 41770 17392
rect 41804 17358 41860 17392
rect 41894 17358 41950 17392
rect 41984 17358 42040 17392
rect 42074 17358 42130 17392
rect 42164 17358 42220 17392
rect 42254 17358 42310 17392
rect 42344 17358 42400 17392
rect 42434 17358 42770 17392
rect 42804 17358 42860 17392
rect 42894 17358 42950 17392
rect 42984 17358 43040 17392
rect 43074 17358 43130 17392
rect 43164 17358 43220 17392
rect 43254 17358 43310 17392
rect 43344 17358 43400 17392
rect 43434 17358 43490 17392
rect 43524 17358 43580 17392
rect 43614 17358 43670 17392
rect 43704 17358 43760 17392
rect 43794 17358 44130 17392
rect 44164 17358 44220 17392
rect 44254 17358 44310 17392
rect 44344 17358 44400 17392
rect 44434 17358 44490 17392
rect 44524 17358 44580 17392
rect 44614 17358 44670 17392
rect 44704 17358 44760 17392
rect 44794 17358 44850 17392
rect 44884 17358 44940 17392
rect 44974 17358 45030 17392
rect 45064 17358 45120 17392
rect 45154 17358 45284 17392
rect 41276 17325 45284 17358
rect 41276 17308 41375 17325
rect 41276 17274 41309 17308
rect 41343 17274 41375 17308
rect 41276 17218 41375 17274
rect 42465 17308 42735 17325
rect 42465 17274 42496 17308
rect 42530 17274 42669 17308
rect 42703 17274 42735 17308
rect 41276 17184 41309 17218
rect 41343 17184 41375 17218
rect 41276 17128 41375 17184
rect 41276 17094 41309 17128
rect 41343 17094 41375 17128
rect 41276 17038 41375 17094
rect 41276 17004 41309 17038
rect 41343 17004 41375 17038
rect 41276 16948 41375 17004
rect 41276 16914 41309 16948
rect 41343 16914 41375 16948
rect 41276 16858 41375 16914
rect 41276 16824 41309 16858
rect 41343 16824 41375 16858
rect 41276 16768 41375 16824
rect 41276 16734 41309 16768
rect 41343 16734 41375 16768
rect 41276 16678 41375 16734
rect 41276 16644 41309 16678
rect 41343 16644 41375 16678
rect 41276 16588 41375 16644
rect 41276 16554 41309 16588
rect 41343 16554 41375 16588
rect 41276 16498 41375 16554
rect 41276 16464 41309 16498
rect 41343 16464 41375 16498
rect 41276 16408 41375 16464
rect 41276 16380 41309 16408
rect 40913 16181 40947 16243
rect 40163 16147 40259 16181
rect 40851 16147 40947 16181
rect 41270 16374 41309 16380
rect 41343 16380 41375 16408
rect 41439 17242 42401 17261
rect 41439 17208 41550 17242
rect 41584 17208 41640 17242
rect 41674 17208 41730 17242
rect 41764 17208 41820 17242
rect 41854 17208 41910 17242
rect 41944 17208 42000 17242
rect 42034 17208 42090 17242
rect 42124 17208 42180 17242
rect 42214 17208 42270 17242
rect 42304 17208 42401 17242
rect 41439 17189 42401 17208
rect 41439 17148 41511 17189
rect 41439 17114 41458 17148
rect 41492 17114 41511 17148
rect 42329 17129 42401 17189
rect 41439 17058 41511 17114
rect 41439 17024 41458 17058
rect 41492 17024 41511 17058
rect 41439 16968 41511 17024
rect 41439 16934 41458 16968
rect 41492 16934 41511 16968
rect 41439 16878 41511 16934
rect 41439 16844 41458 16878
rect 41492 16844 41511 16878
rect 41439 16788 41511 16844
rect 41439 16754 41458 16788
rect 41492 16754 41511 16788
rect 41439 16698 41511 16754
rect 41439 16664 41458 16698
rect 41492 16664 41511 16698
rect 41439 16608 41511 16664
rect 41439 16574 41458 16608
rect 41492 16574 41511 16608
rect 41439 16518 41511 16574
rect 41439 16484 41458 16518
rect 41492 16484 41511 16518
rect 41439 16428 41511 16484
rect 41573 17066 42267 17127
rect 41573 17032 41632 17066
rect 41666 17054 41722 17066
rect 41694 17032 41722 17054
rect 41756 17054 41812 17066
rect 41756 17032 41760 17054
rect 41573 17020 41660 17032
rect 41694 17020 41760 17032
rect 41794 17032 41812 17054
rect 41846 17054 41902 17066
rect 41846 17032 41860 17054
rect 41794 17020 41860 17032
rect 41894 17032 41902 17054
rect 41936 17054 41992 17066
rect 42026 17054 42082 17066
rect 42116 17054 42172 17066
rect 41936 17032 41960 17054
rect 42026 17032 42060 17054
rect 42116 17032 42160 17054
rect 42206 17032 42267 17066
rect 41894 17020 41960 17032
rect 41994 17020 42060 17032
rect 42094 17020 42160 17032
rect 42194 17020 42267 17032
rect 41573 16976 42267 17020
rect 41573 16942 41632 16976
rect 41666 16954 41722 16976
rect 41694 16942 41722 16954
rect 41756 16954 41812 16976
rect 41756 16942 41760 16954
rect 41573 16920 41660 16942
rect 41694 16920 41760 16942
rect 41794 16942 41812 16954
rect 41846 16954 41902 16976
rect 41846 16942 41860 16954
rect 41794 16920 41860 16942
rect 41894 16942 41902 16954
rect 41936 16954 41992 16976
rect 42026 16954 42082 16976
rect 42116 16954 42172 16976
rect 41936 16942 41960 16954
rect 42026 16942 42060 16954
rect 42116 16942 42160 16954
rect 42206 16942 42267 16976
rect 41894 16920 41960 16942
rect 41994 16920 42060 16942
rect 42094 16920 42160 16942
rect 42194 16920 42267 16942
rect 41573 16886 42267 16920
rect 41573 16852 41632 16886
rect 41666 16854 41722 16886
rect 41694 16852 41722 16854
rect 41756 16854 41812 16886
rect 41756 16852 41760 16854
rect 41573 16820 41660 16852
rect 41694 16820 41760 16852
rect 41794 16852 41812 16854
rect 41846 16854 41902 16886
rect 41846 16852 41860 16854
rect 41794 16820 41860 16852
rect 41894 16852 41902 16854
rect 41936 16854 41992 16886
rect 42026 16854 42082 16886
rect 42116 16854 42172 16886
rect 41936 16852 41960 16854
rect 42026 16852 42060 16854
rect 42116 16852 42160 16854
rect 42206 16852 42267 16886
rect 41894 16820 41960 16852
rect 41994 16820 42060 16852
rect 42094 16820 42160 16852
rect 42194 16820 42267 16852
rect 41573 16796 42267 16820
rect 41573 16762 41632 16796
rect 41666 16762 41722 16796
rect 41756 16762 41812 16796
rect 41846 16762 41902 16796
rect 41936 16762 41992 16796
rect 42026 16762 42082 16796
rect 42116 16762 42172 16796
rect 42206 16762 42267 16796
rect 41573 16754 42267 16762
rect 41573 16720 41660 16754
rect 41694 16720 41760 16754
rect 41794 16720 41860 16754
rect 41894 16720 41960 16754
rect 41994 16720 42060 16754
rect 42094 16720 42160 16754
rect 42194 16720 42267 16754
rect 41573 16706 42267 16720
rect 41573 16672 41632 16706
rect 41666 16672 41722 16706
rect 41756 16672 41812 16706
rect 41846 16672 41902 16706
rect 41936 16672 41992 16706
rect 42026 16672 42082 16706
rect 42116 16672 42172 16706
rect 42206 16672 42267 16706
rect 41573 16654 42267 16672
rect 41573 16620 41660 16654
rect 41694 16620 41760 16654
rect 41794 16620 41860 16654
rect 41894 16620 41960 16654
rect 41994 16620 42060 16654
rect 42094 16620 42160 16654
rect 42194 16620 42267 16654
rect 41573 16616 42267 16620
rect 41573 16582 41632 16616
rect 41666 16582 41722 16616
rect 41756 16582 41812 16616
rect 41846 16582 41902 16616
rect 41936 16582 41992 16616
rect 42026 16582 42082 16616
rect 42116 16582 42172 16616
rect 42206 16582 42267 16616
rect 41573 16554 42267 16582
rect 41573 16526 41660 16554
rect 41694 16526 41760 16554
rect 41573 16492 41632 16526
rect 41694 16520 41722 16526
rect 41666 16492 41722 16520
rect 41756 16520 41760 16526
rect 41794 16526 41860 16554
rect 41794 16520 41812 16526
rect 41756 16492 41812 16520
rect 41846 16520 41860 16526
rect 41894 16526 41960 16554
rect 41994 16526 42060 16554
rect 42094 16526 42160 16554
rect 42194 16526 42267 16554
rect 41894 16520 41902 16526
rect 41846 16492 41902 16520
rect 41936 16520 41960 16526
rect 42026 16520 42060 16526
rect 42116 16520 42160 16526
rect 41936 16492 41992 16520
rect 42026 16492 42082 16520
rect 42116 16492 42172 16520
rect 42206 16492 42267 16526
rect 41573 16433 42267 16492
rect 42329 17095 42348 17129
rect 42382 17095 42401 17129
rect 42329 17039 42401 17095
rect 42329 17005 42348 17039
rect 42382 17005 42401 17039
rect 42329 16949 42401 17005
rect 42329 16915 42348 16949
rect 42382 16915 42401 16949
rect 42329 16859 42401 16915
rect 42329 16825 42348 16859
rect 42382 16825 42401 16859
rect 42329 16769 42401 16825
rect 42329 16735 42348 16769
rect 42382 16735 42401 16769
rect 42329 16679 42401 16735
rect 42329 16645 42348 16679
rect 42382 16645 42401 16679
rect 42329 16589 42401 16645
rect 42329 16555 42348 16589
rect 42382 16555 42401 16589
rect 42329 16499 42401 16555
rect 42329 16465 42348 16499
rect 42382 16465 42401 16499
rect 41439 16394 41458 16428
rect 41492 16394 41511 16428
rect 41439 16380 41511 16394
rect 42329 16409 42401 16465
rect 42329 16380 42348 16409
rect 41343 16375 42348 16380
rect 42382 16380 42401 16409
rect 42465 17218 42735 17274
rect 43825 17308 44095 17325
rect 43825 17274 43856 17308
rect 43890 17274 44029 17308
rect 44063 17274 44095 17308
rect 42465 17184 42496 17218
rect 42530 17184 42669 17218
rect 42703 17184 42735 17218
rect 42465 17128 42735 17184
rect 42465 17094 42496 17128
rect 42530 17094 42669 17128
rect 42703 17094 42735 17128
rect 42465 17038 42735 17094
rect 42465 17004 42496 17038
rect 42530 17004 42669 17038
rect 42703 17004 42735 17038
rect 42465 16948 42735 17004
rect 42465 16914 42496 16948
rect 42530 16914 42669 16948
rect 42703 16914 42735 16948
rect 42465 16858 42735 16914
rect 42465 16824 42496 16858
rect 42530 16824 42669 16858
rect 42703 16824 42735 16858
rect 42465 16768 42735 16824
rect 42465 16734 42496 16768
rect 42530 16734 42669 16768
rect 42703 16734 42735 16768
rect 42465 16678 42735 16734
rect 42465 16644 42496 16678
rect 42530 16644 42669 16678
rect 42703 16644 42735 16678
rect 42465 16588 42735 16644
rect 42465 16554 42496 16588
rect 42530 16554 42669 16588
rect 42703 16554 42735 16588
rect 42465 16498 42735 16554
rect 42465 16464 42496 16498
rect 42530 16464 42669 16498
rect 42703 16464 42735 16498
rect 42465 16408 42735 16464
rect 42465 16380 42496 16408
rect 42382 16375 42496 16380
rect 41343 16374 42496 16375
rect 42530 16374 42669 16408
rect 42703 16380 42735 16408
rect 42799 17242 43761 17261
rect 42799 17208 42910 17242
rect 42944 17208 43000 17242
rect 43034 17208 43090 17242
rect 43124 17208 43180 17242
rect 43214 17208 43270 17242
rect 43304 17208 43360 17242
rect 43394 17208 43450 17242
rect 43484 17208 43540 17242
rect 43574 17208 43630 17242
rect 43664 17208 43761 17242
rect 42799 17189 43761 17208
rect 42799 17148 42871 17189
rect 42799 17114 42818 17148
rect 42852 17114 42871 17148
rect 43689 17129 43761 17189
rect 42799 17058 42871 17114
rect 42799 17024 42818 17058
rect 42852 17024 42871 17058
rect 42799 16968 42871 17024
rect 42799 16934 42818 16968
rect 42852 16934 42871 16968
rect 42799 16878 42871 16934
rect 42799 16844 42818 16878
rect 42852 16844 42871 16878
rect 42799 16788 42871 16844
rect 42799 16754 42818 16788
rect 42852 16754 42871 16788
rect 42799 16698 42871 16754
rect 42799 16664 42818 16698
rect 42852 16664 42871 16698
rect 42799 16608 42871 16664
rect 42799 16574 42818 16608
rect 42852 16574 42871 16608
rect 42799 16518 42871 16574
rect 42799 16484 42818 16518
rect 42852 16484 42871 16518
rect 42799 16428 42871 16484
rect 42933 17066 43627 17127
rect 42933 17032 42992 17066
rect 43026 17054 43082 17066
rect 43054 17032 43082 17054
rect 43116 17054 43172 17066
rect 43116 17032 43120 17054
rect 42933 17020 43020 17032
rect 43054 17020 43120 17032
rect 43154 17032 43172 17054
rect 43206 17054 43262 17066
rect 43206 17032 43220 17054
rect 43154 17020 43220 17032
rect 43254 17032 43262 17054
rect 43296 17054 43352 17066
rect 43386 17054 43442 17066
rect 43476 17054 43532 17066
rect 43296 17032 43320 17054
rect 43386 17032 43420 17054
rect 43476 17032 43520 17054
rect 43566 17032 43627 17066
rect 43254 17020 43320 17032
rect 43354 17020 43420 17032
rect 43454 17020 43520 17032
rect 43554 17020 43627 17032
rect 42933 16976 43627 17020
rect 42933 16942 42992 16976
rect 43026 16954 43082 16976
rect 43054 16942 43082 16954
rect 43116 16954 43172 16976
rect 43116 16942 43120 16954
rect 42933 16920 43020 16942
rect 43054 16920 43120 16942
rect 43154 16942 43172 16954
rect 43206 16954 43262 16976
rect 43206 16942 43220 16954
rect 43154 16920 43220 16942
rect 43254 16942 43262 16954
rect 43296 16954 43352 16976
rect 43386 16954 43442 16976
rect 43476 16954 43532 16976
rect 43296 16942 43320 16954
rect 43386 16942 43420 16954
rect 43476 16942 43520 16954
rect 43566 16942 43627 16976
rect 43254 16920 43320 16942
rect 43354 16920 43420 16942
rect 43454 16920 43520 16942
rect 43554 16920 43627 16942
rect 42933 16886 43627 16920
rect 42933 16852 42992 16886
rect 43026 16854 43082 16886
rect 43054 16852 43082 16854
rect 43116 16854 43172 16886
rect 43116 16852 43120 16854
rect 42933 16820 43020 16852
rect 43054 16820 43120 16852
rect 43154 16852 43172 16854
rect 43206 16854 43262 16886
rect 43206 16852 43220 16854
rect 43154 16820 43220 16852
rect 43254 16852 43262 16854
rect 43296 16854 43352 16886
rect 43386 16854 43442 16886
rect 43476 16854 43532 16886
rect 43296 16852 43320 16854
rect 43386 16852 43420 16854
rect 43476 16852 43520 16854
rect 43566 16852 43627 16886
rect 43254 16820 43320 16852
rect 43354 16820 43420 16852
rect 43454 16820 43520 16852
rect 43554 16820 43627 16852
rect 42933 16796 43627 16820
rect 42933 16762 42992 16796
rect 43026 16762 43082 16796
rect 43116 16762 43172 16796
rect 43206 16762 43262 16796
rect 43296 16762 43352 16796
rect 43386 16762 43442 16796
rect 43476 16762 43532 16796
rect 43566 16762 43627 16796
rect 42933 16754 43627 16762
rect 42933 16720 43020 16754
rect 43054 16720 43120 16754
rect 43154 16720 43220 16754
rect 43254 16720 43320 16754
rect 43354 16720 43420 16754
rect 43454 16720 43520 16754
rect 43554 16720 43627 16754
rect 42933 16706 43627 16720
rect 42933 16672 42992 16706
rect 43026 16672 43082 16706
rect 43116 16672 43172 16706
rect 43206 16672 43262 16706
rect 43296 16672 43352 16706
rect 43386 16672 43442 16706
rect 43476 16672 43532 16706
rect 43566 16672 43627 16706
rect 42933 16654 43627 16672
rect 42933 16620 43020 16654
rect 43054 16620 43120 16654
rect 43154 16620 43220 16654
rect 43254 16620 43320 16654
rect 43354 16620 43420 16654
rect 43454 16620 43520 16654
rect 43554 16620 43627 16654
rect 42933 16616 43627 16620
rect 42933 16582 42992 16616
rect 43026 16582 43082 16616
rect 43116 16582 43172 16616
rect 43206 16582 43262 16616
rect 43296 16582 43352 16616
rect 43386 16582 43442 16616
rect 43476 16582 43532 16616
rect 43566 16582 43627 16616
rect 42933 16554 43627 16582
rect 42933 16526 43020 16554
rect 43054 16526 43120 16554
rect 42933 16492 42992 16526
rect 43054 16520 43082 16526
rect 43026 16492 43082 16520
rect 43116 16520 43120 16526
rect 43154 16526 43220 16554
rect 43154 16520 43172 16526
rect 43116 16492 43172 16520
rect 43206 16520 43220 16526
rect 43254 16526 43320 16554
rect 43354 16526 43420 16554
rect 43454 16526 43520 16554
rect 43554 16526 43627 16554
rect 43254 16520 43262 16526
rect 43206 16492 43262 16520
rect 43296 16520 43320 16526
rect 43386 16520 43420 16526
rect 43476 16520 43520 16526
rect 43296 16492 43352 16520
rect 43386 16492 43442 16520
rect 43476 16492 43532 16520
rect 43566 16492 43627 16526
rect 42933 16433 43627 16492
rect 43689 17095 43708 17129
rect 43742 17095 43761 17129
rect 43689 17039 43761 17095
rect 43689 17005 43708 17039
rect 43742 17005 43761 17039
rect 43689 16949 43761 17005
rect 43689 16915 43708 16949
rect 43742 16915 43761 16949
rect 43689 16859 43761 16915
rect 43689 16825 43708 16859
rect 43742 16825 43761 16859
rect 43689 16769 43761 16825
rect 43689 16735 43708 16769
rect 43742 16735 43761 16769
rect 43689 16679 43761 16735
rect 43689 16645 43708 16679
rect 43742 16645 43761 16679
rect 43689 16589 43761 16645
rect 43689 16555 43708 16589
rect 43742 16555 43761 16589
rect 43689 16499 43761 16555
rect 43689 16465 43708 16499
rect 43742 16465 43761 16499
rect 42799 16394 42818 16428
rect 42852 16394 42871 16428
rect 42799 16380 42871 16394
rect 43689 16409 43761 16465
rect 43689 16380 43708 16409
rect 42703 16375 43708 16380
rect 43742 16380 43761 16409
rect 43825 17218 44095 17274
rect 45185 17308 45284 17325
rect 45185 17274 45216 17308
rect 45250 17274 45284 17308
rect 43825 17184 43856 17218
rect 43890 17184 44029 17218
rect 44063 17184 44095 17218
rect 43825 17128 44095 17184
rect 43825 17094 43856 17128
rect 43890 17094 44029 17128
rect 44063 17094 44095 17128
rect 43825 17038 44095 17094
rect 43825 17004 43856 17038
rect 43890 17004 44029 17038
rect 44063 17004 44095 17038
rect 43825 16948 44095 17004
rect 43825 16914 43856 16948
rect 43890 16914 44029 16948
rect 44063 16914 44095 16948
rect 43825 16858 44095 16914
rect 43825 16824 43856 16858
rect 43890 16824 44029 16858
rect 44063 16824 44095 16858
rect 43825 16768 44095 16824
rect 43825 16734 43856 16768
rect 43890 16734 44029 16768
rect 44063 16734 44095 16768
rect 43825 16678 44095 16734
rect 43825 16644 43856 16678
rect 43890 16644 44029 16678
rect 44063 16644 44095 16678
rect 43825 16588 44095 16644
rect 43825 16554 43856 16588
rect 43890 16554 44029 16588
rect 44063 16554 44095 16588
rect 43825 16498 44095 16554
rect 43825 16464 43856 16498
rect 43890 16464 44029 16498
rect 44063 16464 44095 16498
rect 43825 16408 44095 16464
rect 43825 16380 43856 16408
rect 43742 16375 43856 16380
rect 42703 16374 43856 16375
rect 43890 16374 44029 16408
rect 44063 16380 44095 16408
rect 44159 17242 45121 17261
rect 44159 17208 44270 17242
rect 44304 17208 44360 17242
rect 44394 17208 44450 17242
rect 44484 17208 44540 17242
rect 44574 17208 44630 17242
rect 44664 17208 44720 17242
rect 44754 17208 44810 17242
rect 44844 17208 44900 17242
rect 44934 17208 44990 17242
rect 45024 17208 45121 17242
rect 44159 17189 45121 17208
rect 44159 17148 44231 17189
rect 44159 17114 44178 17148
rect 44212 17114 44231 17148
rect 45049 17129 45121 17189
rect 44159 17058 44231 17114
rect 44159 17024 44178 17058
rect 44212 17024 44231 17058
rect 44159 16968 44231 17024
rect 44159 16934 44178 16968
rect 44212 16934 44231 16968
rect 44159 16878 44231 16934
rect 44159 16844 44178 16878
rect 44212 16844 44231 16878
rect 44159 16788 44231 16844
rect 44159 16754 44178 16788
rect 44212 16754 44231 16788
rect 44159 16698 44231 16754
rect 44159 16664 44178 16698
rect 44212 16664 44231 16698
rect 44159 16608 44231 16664
rect 44159 16574 44178 16608
rect 44212 16574 44231 16608
rect 44159 16518 44231 16574
rect 44159 16484 44178 16518
rect 44212 16484 44231 16518
rect 44159 16428 44231 16484
rect 44293 17066 44987 17127
rect 44293 17032 44352 17066
rect 44386 17054 44442 17066
rect 44414 17032 44442 17054
rect 44476 17054 44532 17066
rect 44476 17032 44480 17054
rect 44293 17020 44380 17032
rect 44414 17020 44480 17032
rect 44514 17032 44532 17054
rect 44566 17054 44622 17066
rect 44566 17032 44580 17054
rect 44514 17020 44580 17032
rect 44614 17032 44622 17054
rect 44656 17054 44712 17066
rect 44746 17054 44802 17066
rect 44836 17054 44892 17066
rect 44656 17032 44680 17054
rect 44746 17032 44780 17054
rect 44836 17032 44880 17054
rect 44926 17032 44987 17066
rect 44614 17020 44680 17032
rect 44714 17020 44780 17032
rect 44814 17020 44880 17032
rect 44914 17020 44987 17032
rect 44293 16976 44987 17020
rect 44293 16942 44352 16976
rect 44386 16954 44442 16976
rect 44414 16942 44442 16954
rect 44476 16954 44532 16976
rect 44476 16942 44480 16954
rect 44293 16920 44380 16942
rect 44414 16920 44480 16942
rect 44514 16942 44532 16954
rect 44566 16954 44622 16976
rect 44566 16942 44580 16954
rect 44514 16920 44580 16942
rect 44614 16942 44622 16954
rect 44656 16954 44712 16976
rect 44746 16954 44802 16976
rect 44836 16954 44892 16976
rect 44656 16942 44680 16954
rect 44746 16942 44780 16954
rect 44836 16942 44880 16954
rect 44926 16942 44987 16976
rect 44614 16920 44680 16942
rect 44714 16920 44780 16942
rect 44814 16920 44880 16942
rect 44914 16920 44987 16942
rect 44293 16886 44987 16920
rect 44293 16852 44352 16886
rect 44386 16854 44442 16886
rect 44414 16852 44442 16854
rect 44476 16854 44532 16886
rect 44476 16852 44480 16854
rect 44293 16820 44380 16852
rect 44414 16820 44480 16852
rect 44514 16852 44532 16854
rect 44566 16854 44622 16886
rect 44566 16852 44580 16854
rect 44514 16820 44580 16852
rect 44614 16852 44622 16854
rect 44656 16854 44712 16886
rect 44746 16854 44802 16886
rect 44836 16854 44892 16886
rect 44656 16852 44680 16854
rect 44746 16852 44780 16854
rect 44836 16852 44880 16854
rect 44926 16852 44987 16886
rect 44614 16820 44680 16852
rect 44714 16820 44780 16852
rect 44814 16820 44880 16852
rect 44914 16820 44987 16852
rect 44293 16796 44987 16820
rect 44293 16762 44352 16796
rect 44386 16762 44442 16796
rect 44476 16762 44532 16796
rect 44566 16762 44622 16796
rect 44656 16762 44712 16796
rect 44746 16762 44802 16796
rect 44836 16762 44892 16796
rect 44926 16762 44987 16796
rect 44293 16754 44987 16762
rect 44293 16720 44380 16754
rect 44414 16720 44480 16754
rect 44514 16720 44580 16754
rect 44614 16720 44680 16754
rect 44714 16720 44780 16754
rect 44814 16720 44880 16754
rect 44914 16720 44987 16754
rect 44293 16706 44987 16720
rect 44293 16672 44352 16706
rect 44386 16672 44442 16706
rect 44476 16672 44532 16706
rect 44566 16672 44622 16706
rect 44656 16672 44712 16706
rect 44746 16672 44802 16706
rect 44836 16672 44892 16706
rect 44926 16672 44987 16706
rect 44293 16654 44987 16672
rect 44293 16620 44380 16654
rect 44414 16620 44480 16654
rect 44514 16620 44580 16654
rect 44614 16620 44680 16654
rect 44714 16620 44780 16654
rect 44814 16620 44880 16654
rect 44914 16620 44987 16654
rect 44293 16616 44987 16620
rect 44293 16582 44352 16616
rect 44386 16582 44442 16616
rect 44476 16582 44532 16616
rect 44566 16582 44622 16616
rect 44656 16582 44712 16616
rect 44746 16582 44802 16616
rect 44836 16582 44892 16616
rect 44926 16582 44987 16616
rect 44293 16554 44987 16582
rect 44293 16526 44380 16554
rect 44414 16526 44480 16554
rect 44293 16492 44352 16526
rect 44414 16520 44442 16526
rect 44386 16492 44442 16520
rect 44476 16520 44480 16526
rect 44514 16526 44580 16554
rect 44514 16520 44532 16526
rect 44476 16492 44532 16520
rect 44566 16520 44580 16526
rect 44614 16526 44680 16554
rect 44714 16526 44780 16554
rect 44814 16526 44880 16554
rect 44914 16526 44987 16554
rect 44614 16520 44622 16526
rect 44566 16492 44622 16520
rect 44656 16520 44680 16526
rect 44746 16520 44780 16526
rect 44836 16520 44880 16526
rect 44656 16492 44712 16520
rect 44746 16492 44802 16520
rect 44836 16492 44892 16520
rect 44926 16492 44987 16526
rect 44293 16433 44987 16492
rect 45049 17095 45068 17129
rect 45102 17095 45121 17129
rect 45049 17039 45121 17095
rect 45049 17005 45068 17039
rect 45102 17005 45121 17039
rect 45049 16949 45121 17005
rect 45049 16915 45068 16949
rect 45102 16915 45121 16949
rect 45049 16859 45121 16915
rect 45049 16825 45068 16859
rect 45102 16825 45121 16859
rect 45049 16769 45121 16825
rect 45049 16735 45068 16769
rect 45102 16735 45121 16769
rect 45049 16679 45121 16735
rect 45049 16645 45068 16679
rect 45102 16645 45121 16679
rect 45049 16589 45121 16645
rect 45049 16555 45068 16589
rect 45102 16555 45121 16589
rect 45049 16499 45121 16555
rect 45049 16465 45068 16499
rect 45102 16465 45121 16499
rect 44159 16394 44178 16428
rect 44212 16394 44231 16428
rect 44159 16380 44231 16394
rect 45049 16409 45121 16465
rect 45049 16380 45068 16409
rect 44063 16375 45068 16380
rect 45102 16380 45121 16409
rect 45185 17218 45284 17274
rect 45185 17184 45216 17218
rect 45250 17184 45284 17218
rect 45185 17128 45284 17184
rect 45185 17094 45216 17128
rect 45250 17094 45284 17128
rect 45185 17038 45284 17094
rect 45185 17004 45216 17038
rect 45250 17004 45284 17038
rect 45185 16948 45284 17004
rect 45185 16914 45216 16948
rect 45250 16914 45284 16948
rect 45185 16858 45284 16914
rect 45185 16824 45216 16858
rect 45250 16824 45284 16858
rect 45185 16768 45284 16824
rect 45185 16734 45216 16768
rect 45250 16734 45284 16768
rect 45185 16678 45284 16734
rect 45185 16644 45216 16678
rect 45250 16644 45284 16678
rect 45185 16588 45284 16644
rect 45185 16554 45216 16588
rect 45250 16554 45284 16588
rect 45185 16498 45284 16554
rect 45185 16464 45216 16498
rect 45250 16464 45284 16498
rect 45185 16408 45284 16464
rect 45185 16380 45216 16408
rect 45102 16375 45216 16380
rect 44063 16374 45216 16375
rect 45250 16380 45284 16408
rect 45250 16374 45290 16380
rect 41270 16352 45290 16374
rect 41270 16318 41516 16352
rect 41550 16318 41606 16352
rect 41640 16318 41696 16352
rect 41730 16318 41786 16352
rect 41820 16318 41876 16352
rect 41910 16318 41966 16352
rect 42000 16318 42056 16352
rect 42090 16318 42146 16352
rect 42180 16318 42236 16352
rect 42270 16318 42876 16352
rect 42910 16318 42966 16352
rect 43000 16318 43056 16352
rect 43090 16318 43146 16352
rect 43180 16318 43236 16352
rect 43270 16318 43326 16352
rect 43360 16318 43416 16352
rect 43450 16318 43506 16352
rect 43540 16318 43596 16352
rect 43630 16318 44236 16352
rect 44270 16318 44326 16352
rect 44360 16318 44416 16352
rect 44450 16318 44506 16352
rect 44540 16318 44596 16352
rect 44630 16318 44686 16352
rect 44720 16318 44776 16352
rect 44810 16318 44866 16352
rect 44900 16318 44956 16352
rect 44990 16318 45290 16352
rect 41270 16284 41309 16318
rect 41343 16284 42496 16318
rect 42530 16284 42669 16318
rect 42703 16284 43856 16318
rect 43890 16284 44029 16318
rect 44063 16284 45216 16318
rect 45250 16284 45290 16318
rect 41270 16228 45290 16284
rect 41270 16194 41309 16228
rect 41343 16205 42496 16228
rect 41343 16194 41410 16205
rect 41270 16171 41410 16194
rect 41444 16171 41500 16205
rect 41534 16171 41590 16205
rect 41624 16171 41680 16205
rect 41714 16171 41770 16205
rect 41804 16171 41860 16205
rect 41894 16171 41950 16205
rect 41984 16171 42040 16205
rect 42074 16171 42130 16205
rect 42164 16171 42220 16205
rect 42254 16171 42310 16205
rect 42344 16171 42400 16205
rect 42434 16194 42496 16205
rect 42530 16194 42669 16228
rect 42703 16205 43856 16228
rect 42703 16194 42770 16205
rect 42434 16171 42770 16194
rect 42804 16171 42860 16205
rect 42894 16171 42950 16205
rect 42984 16171 43040 16205
rect 43074 16171 43130 16205
rect 43164 16171 43220 16205
rect 43254 16171 43310 16205
rect 43344 16171 43400 16205
rect 43434 16171 43490 16205
rect 43524 16171 43580 16205
rect 43614 16171 43670 16205
rect 43704 16171 43760 16205
rect 43794 16194 43856 16205
rect 43890 16194 44029 16228
rect 44063 16205 45216 16228
rect 44063 16194 44130 16205
rect 43794 16171 44130 16194
rect 44164 16171 44220 16205
rect 44254 16171 44310 16205
rect 44344 16171 44400 16205
rect 44434 16171 44490 16205
rect 44524 16171 44580 16205
rect 44614 16171 44670 16205
rect 44704 16171 44760 16205
rect 44794 16171 44850 16205
rect 44884 16171 44940 16205
rect 44974 16171 45030 16205
rect 45064 16171 45120 16205
rect 45154 16194 45216 16205
rect 45250 16194 45290 16228
rect 45154 16171 45290 16194
rect 41270 16130 45290 16171
rect 46233 18501 46267 18563
rect 45483 16181 45517 16243
rect 46233 16181 46267 16243
rect 45483 16147 45579 16181
rect 46171 16147 46267 16181
rect 46593 18561 46689 18595
rect 46949 18561 47045 18595
rect 47570 18590 47650 18610
rect 47570 18589 47590 18590
rect 47630 18589 47650 18590
rect 46593 18499 46627 18561
rect 46780 18550 46860 18561
rect 42560 16064 42640 16130
rect 43920 16064 44000 16130
rect 41276 16032 45284 16064
rect 41276 15998 41410 16032
rect 41444 15998 41500 16032
rect 41534 15998 41590 16032
rect 41624 15998 41680 16032
rect 41714 15998 41770 16032
rect 41804 15998 41860 16032
rect 41894 15998 41950 16032
rect 41984 15998 42040 16032
rect 42074 15998 42130 16032
rect 42164 15998 42220 16032
rect 42254 15998 42310 16032
rect 42344 15998 42400 16032
rect 42434 15998 42770 16032
rect 42804 15998 42860 16032
rect 42894 15998 42950 16032
rect 42984 15998 43040 16032
rect 43074 15998 43130 16032
rect 43164 15998 43220 16032
rect 43254 15998 43310 16032
rect 43344 15998 43400 16032
rect 43434 15998 43490 16032
rect 43524 15998 43580 16032
rect 43614 15998 43670 16032
rect 43704 15998 43760 16032
rect 43794 15998 44130 16032
rect 44164 15998 44220 16032
rect 44254 15998 44310 16032
rect 44344 15998 44400 16032
rect 44434 15998 44490 16032
rect 44524 15998 44580 16032
rect 44614 15998 44670 16032
rect 44704 15998 44760 16032
rect 44794 15998 44850 16032
rect 44884 15998 44940 16032
rect 44974 15998 45030 16032
rect 45064 15998 45120 16032
rect 45154 15998 45284 16032
rect 41276 15965 45284 15998
rect 41276 15948 41375 15965
rect 41276 15914 41309 15948
rect 41343 15914 41375 15948
rect 41276 15858 41375 15914
rect 42465 15948 42735 15965
rect 42465 15914 42496 15948
rect 42530 15914 42669 15948
rect 42703 15914 42735 15948
rect 41276 15824 41309 15858
rect 41343 15824 41375 15858
rect 41276 15768 41375 15824
rect 41276 15734 41309 15768
rect 41343 15734 41375 15768
rect 41276 15678 41375 15734
rect 41276 15644 41309 15678
rect 41343 15644 41375 15678
rect 41276 15588 41375 15644
rect 41276 15554 41309 15588
rect 41343 15554 41375 15588
rect 41276 15498 41375 15554
rect 41276 15464 41309 15498
rect 41343 15464 41375 15498
rect 41276 15408 41375 15464
rect 41276 15374 41309 15408
rect 41343 15374 41375 15408
rect 41276 15318 41375 15374
rect 41276 15284 41309 15318
rect 41343 15284 41375 15318
rect 41276 15228 41375 15284
rect 41276 15194 41309 15228
rect 41343 15194 41375 15228
rect 41276 15138 41375 15194
rect 41276 15104 41309 15138
rect 41343 15104 41375 15138
rect 41276 15048 41375 15104
rect 41276 15020 41309 15048
rect 39801 14957 39835 15019
rect 39383 14923 39479 14957
rect 39739 14923 39835 14957
rect 41270 15014 41309 15020
rect 41343 15020 41375 15048
rect 41439 15882 42401 15901
rect 41439 15848 41550 15882
rect 41584 15848 41640 15882
rect 41674 15848 41730 15882
rect 41764 15848 41820 15882
rect 41854 15848 41910 15882
rect 41944 15848 42000 15882
rect 42034 15848 42090 15882
rect 42124 15848 42180 15882
rect 42214 15848 42270 15882
rect 42304 15848 42401 15882
rect 41439 15829 42401 15848
rect 41439 15788 41511 15829
rect 41439 15754 41458 15788
rect 41492 15754 41511 15788
rect 42329 15769 42401 15829
rect 41439 15698 41511 15754
rect 41439 15664 41458 15698
rect 41492 15664 41511 15698
rect 41439 15608 41511 15664
rect 41439 15574 41458 15608
rect 41492 15574 41511 15608
rect 41439 15518 41511 15574
rect 41439 15484 41458 15518
rect 41492 15484 41511 15518
rect 41439 15428 41511 15484
rect 41439 15394 41458 15428
rect 41492 15394 41511 15428
rect 41439 15338 41511 15394
rect 41439 15304 41458 15338
rect 41492 15304 41511 15338
rect 41439 15248 41511 15304
rect 41439 15214 41458 15248
rect 41492 15214 41511 15248
rect 41439 15158 41511 15214
rect 41439 15124 41458 15158
rect 41492 15124 41511 15158
rect 41439 15068 41511 15124
rect 41573 15706 42267 15767
rect 41573 15672 41632 15706
rect 41666 15694 41722 15706
rect 41694 15672 41722 15694
rect 41756 15694 41812 15706
rect 41756 15672 41760 15694
rect 41573 15660 41660 15672
rect 41694 15660 41760 15672
rect 41794 15672 41812 15694
rect 41846 15694 41902 15706
rect 41846 15672 41860 15694
rect 41794 15660 41860 15672
rect 41894 15672 41902 15694
rect 41936 15694 41992 15706
rect 42026 15694 42082 15706
rect 42116 15694 42172 15706
rect 41936 15672 41960 15694
rect 42026 15672 42060 15694
rect 42116 15672 42160 15694
rect 42206 15672 42267 15706
rect 41894 15660 41960 15672
rect 41994 15660 42060 15672
rect 42094 15660 42160 15672
rect 42194 15660 42267 15672
rect 41573 15616 42267 15660
rect 41573 15582 41632 15616
rect 41666 15594 41722 15616
rect 41694 15582 41722 15594
rect 41756 15594 41812 15616
rect 41756 15582 41760 15594
rect 41573 15560 41660 15582
rect 41694 15560 41760 15582
rect 41794 15582 41812 15594
rect 41846 15594 41902 15616
rect 41846 15582 41860 15594
rect 41794 15560 41860 15582
rect 41894 15582 41902 15594
rect 41936 15594 41992 15616
rect 42026 15594 42082 15616
rect 42116 15594 42172 15616
rect 41936 15582 41960 15594
rect 42026 15582 42060 15594
rect 42116 15582 42160 15594
rect 42206 15582 42267 15616
rect 41894 15560 41960 15582
rect 41994 15560 42060 15582
rect 42094 15560 42160 15582
rect 42194 15560 42267 15582
rect 41573 15526 42267 15560
rect 41573 15492 41632 15526
rect 41666 15494 41722 15526
rect 41694 15492 41722 15494
rect 41756 15494 41812 15526
rect 41756 15492 41760 15494
rect 41573 15460 41660 15492
rect 41694 15460 41760 15492
rect 41794 15492 41812 15494
rect 41846 15494 41902 15526
rect 41846 15492 41860 15494
rect 41794 15460 41860 15492
rect 41894 15492 41902 15494
rect 41936 15494 41992 15526
rect 42026 15494 42082 15526
rect 42116 15494 42172 15526
rect 41936 15492 41960 15494
rect 42026 15492 42060 15494
rect 42116 15492 42160 15494
rect 42206 15492 42267 15526
rect 41894 15460 41960 15492
rect 41994 15460 42060 15492
rect 42094 15460 42160 15492
rect 42194 15460 42267 15492
rect 41573 15436 42267 15460
rect 41573 15402 41632 15436
rect 41666 15402 41722 15436
rect 41756 15402 41812 15436
rect 41846 15402 41902 15436
rect 41936 15402 41992 15436
rect 42026 15402 42082 15436
rect 42116 15402 42172 15436
rect 42206 15402 42267 15436
rect 41573 15394 42267 15402
rect 41573 15360 41660 15394
rect 41694 15360 41760 15394
rect 41794 15360 41860 15394
rect 41894 15360 41960 15394
rect 41994 15360 42060 15394
rect 42094 15360 42160 15394
rect 42194 15360 42267 15394
rect 41573 15346 42267 15360
rect 41573 15312 41632 15346
rect 41666 15312 41722 15346
rect 41756 15312 41812 15346
rect 41846 15312 41902 15346
rect 41936 15312 41992 15346
rect 42026 15312 42082 15346
rect 42116 15312 42172 15346
rect 42206 15312 42267 15346
rect 41573 15294 42267 15312
rect 41573 15260 41660 15294
rect 41694 15260 41760 15294
rect 41794 15260 41860 15294
rect 41894 15260 41960 15294
rect 41994 15260 42060 15294
rect 42094 15260 42160 15294
rect 42194 15260 42267 15294
rect 41573 15256 42267 15260
rect 41573 15222 41632 15256
rect 41666 15222 41722 15256
rect 41756 15222 41812 15256
rect 41846 15222 41902 15256
rect 41936 15222 41992 15256
rect 42026 15222 42082 15256
rect 42116 15222 42172 15256
rect 42206 15222 42267 15256
rect 41573 15194 42267 15222
rect 41573 15166 41660 15194
rect 41694 15166 41760 15194
rect 41573 15132 41632 15166
rect 41694 15160 41722 15166
rect 41666 15132 41722 15160
rect 41756 15160 41760 15166
rect 41794 15166 41860 15194
rect 41794 15160 41812 15166
rect 41756 15132 41812 15160
rect 41846 15160 41860 15166
rect 41894 15166 41960 15194
rect 41994 15166 42060 15194
rect 42094 15166 42160 15194
rect 42194 15166 42267 15194
rect 41894 15160 41902 15166
rect 41846 15132 41902 15160
rect 41936 15160 41960 15166
rect 42026 15160 42060 15166
rect 42116 15160 42160 15166
rect 41936 15132 41992 15160
rect 42026 15132 42082 15160
rect 42116 15132 42172 15160
rect 42206 15132 42267 15166
rect 41573 15073 42267 15132
rect 42329 15735 42348 15769
rect 42382 15735 42401 15769
rect 42329 15679 42401 15735
rect 42329 15645 42348 15679
rect 42382 15645 42401 15679
rect 42329 15589 42401 15645
rect 42329 15555 42348 15589
rect 42382 15555 42401 15589
rect 42329 15499 42401 15555
rect 42329 15465 42348 15499
rect 42382 15465 42401 15499
rect 42329 15409 42401 15465
rect 42329 15375 42348 15409
rect 42382 15375 42401 15409
rect 42329 15319 42401 15375
rect 42329 15285 42348 15319
rect 42382 15285 42401 15319
rect 42329 15229 42401 15285
rect 42329 15195 42348 15229
rect 42382 15195 42401 15229
rect 42329 15139 42401 15195
rect 42329 15105 42348 15139
rect 42382 15105 42401 15139
rect 41439 15034 41458 15068
rect 41492 15034 41511 15068
rect 41439 15020 41511 15034
rect 42329 15049 42401 15105
rect 42329 15020 42348 15049
rect 41343 15015 42348 15020
rect 42382 15020 42401 15049
rect 42465 15858 42735 15914
rect 43825 15948 44095 15965
rect 43825 15914 43856 15948
rect 43890 15914 44029 15948
rect 44063 15914 44095 15948
rect 42465 15824 42496 15858
rect 42530 15824 42669 15858
rect 42703 15824 42735 15858
rect 42465 15768 42735 15824
rect 42465 15734 42496 15768
rect 42530 15734 42669 15768
rect 42703 15734 42735 15768
rect 42465 15678 42735 15734
rect 42465 15644 42496 15678
rect 42530 15644 42669 15678
rect 42703 15644 42735 15678
rect 42465 15588 42735 15644
rect 42465 15554 42496 15588
rect 42530 15554 42669 15588
rect 42703 15554 42735 15588
rect 42465 15498 42735 15554
rect 42465 15464 42496 15498
rect 42530 15464 42669 15498
rect 42703 15464 42735 15498
rect 42465 15408 42735 15464
rect 42465 15374 42496 15408
rect 42530 15374 42669 15408
rect 42703 15374 42735 15408
rect 42465 15318 42735 15374
rect 42465 15284 42496 15318
rect 42530 15284 42669 15318
rect 42703 15284 42735 15318
rect 42465 15228 42735 15284
rect 42465 15194 42496 15228
rect 42530 15194 42669 15228
rect 42703 15194 42735 15228
rect 42465 15138 42735 15194
rect 42465 15104 42496 15138
rect 42530 15104 42669 15138
rect 42703 15104 42735 15138
rect 42465 15048 42735 15104
rect 42465 15020 42496 15048
rect 42382 15015 42496 15020
rect 41343 15014 42496 15015
rect 42530 15014 42669 15048
rect 42703 15020 42735 15048
rect 42799 15882 43761 15901
rect 42799 15848 42910 15882
rect 42944 15848 43000 15882
rect 43034 15848 43090 15882
rect 43124 15848 43180 15882
rect 43214 15848 43270 15882
rect 43304 15848 43360 15882
rect 43394 15848 43450 15882
rect 43484 15848 43540 15882
rect 43574 15848 43630 15882
rect 43664 15848 43761 15882
rect 42799 15829 43761 15848
rect 42799 15788 42871 15829
rect 42799 15754 42818 15788
rect 42852 15754 42871 15788
rect 43689 15769 43761 15829
rect 42799 15698 42871 15754
rect 42799 15664 42818 15698
rect 42852 15664 42871 15698
rect 42799 15608 42871 15664
rect 42799 15574 42818 15608
rect 42852 15574 42871 15608
rect 42799 15518 42871 15574
rect 42799 15484 42818 15518
rect 42852 15484 42871 15518
rect 42799 15428 42871 15484
rect 42799 15394 42818 15428
rect 42852 15394 42871 15428
rect 42799 15338 42871 15394
rect 42799 15304 42818 15338
rect 42852 15304 42871 15338
rect 42799 15248 42871 15304
rect 42799 15214 42818 15248
rect 42852 15214 42871 15248
rect 42799 15158 42871 15214
rect 42799 15124 42818 15158
rect 42852 15124 42871 15158
rect 42799 15068 42871 15124
rect 42933 15706 43627 15767
rect 42933 15672 42992 15706
rect 43026 15694 43082 15706
rect 43054 15672 43082 15694
rect 43116 15694 43172 15706
rect 43116 15672 43120 15694
rect 42933 15660 43020 15672
rect 43054 15660 43120 15672
rect 43154 15672 43172 15694
rect 43206 15694 43262 15706
rect 43206 15672 43220 15694
rect 43154 15660 43220 15672
rect 43254 15672 43262 15694
rect 43296 15694 43352 15706
rect 43386 15694 43442 15706
rect 43476 15694 43532 15706
rect 43296 15672 43320 15694
rect 43386 15672 43420 15694
rect 43476 15672 43520 15694
rect 43566 15672 43627 15706
rect 43254 15660 43320 15672
rect 43354 15660 43420 15672
rect 43454 15660 43520 15672
rect 43554 15660 43627 15672
rect 42933 15616 43627 15660
rect 42933 15582 42992 15616
rect 43026 15594 43082 15616
rect 43054 15582 43082 15594
rect 43116 15594 43172 15616
rect 43116 15582 43120 15594
rect 42933 15560 43020 15582
rect 43054 15560 43120 15582
rect 43154 15582 43172 15594
rect 43206 15594 43262 15616
rect 43206 15582 43220 15594
rect 43154 15560 43220 15582
rect 43254 15582 43262 15594
rect 43296 15594 43352 15616
rect 43386 15594 43442 15616
rect 43476 15594 43532 15616
rect 43296 15582 43320 15594
rect 43386 15582 43420 15594
rect 43476 15582 43520 15594
rect 43566 15582 43627 15616
rect 43254 15560 43320 15582
rect 43354 15560 43420 15582
rect 43454 15560 43520 15582
rect 43554 15560 43627 15582
rect 42933 15526 43627 15560
rect 42933 15492 42992 15526
rect 43026 15494 43082 15526
rect 43054 15492 43082 15494
rect 43116 15494 43172 15526
rect 43116 15492 43120 15494
rect 42933 15460 43020 15492
rect 43054 15460 43120 15492
rect 43154 15492 43172 15494
rect 43206 15494 43262 15526
rect 43206 15492 43220 15494
rect 43154 15460 43220 15492
rect 43254 15492 43262 15494
rect 43296 15494 43352 15526
rect 43386 15494 43442 15526
rect 43476 15494 43532 15526
rect 43296 15492 43320 15494
rect 43386 15492 43420 15494
rect 43476 15492 43520 15494
rect 43566 15492 43627 15526
rect 43254 15460 43320 15492
rect 43354 15460 43420 15492
rect 43454 15460 43520 15492
rect 43554 15460 43627 15492
rect 42933 15436 43627 15460
rect 42933 15402 42992 15436
rect 43026 15402 43082 15436
rect 43116 15402 43172 15436
rect 43206 15402 43262 15436
rect 43296 15402 43352 15436
rect 43386 15402 43442 15436
rect 43476 15402 43532 15436
rect 43566 15402 43627 15436
rect 42933 15394 43627 15402
rect 42933 15360 43020 15394
rect 43054 15360 43120 15394
rect 43154 15360 43220 15394
rect 43254 15360 43320 15394
rect 43354 15360 43420 15394
rect 43454 15360 43520 15394
rect 43554 15360 43627 15394
rect 42933 15346 43627 15360
rect 42933 15312 42992 15346
rect 43026 15312 43082 15346
rect 43116 15312 43172 15346
rect 43206 15312 43262 15346
rect 43296 15312 43352 15346
rect 43386 15312 43442 15346
rect 43476 15312 43532 15346
rect 43566 15312 43627 15346
rect 42933 15294 43627 15312
rect 42933 15260 43020 15294
rect 43054 15260 43120 15294
rect 43154 15260 43220 15294
rect 43254 15260 43320 15294
rect 43354 15260 43420 15294
rect 43454 15260 43520 15294
rect 43554 15260 43627 15294
rect 42933 15256 43627 15260
rect 42933 15222 42992 15256
rect 43026 15222 43082 15256
rect 43116 15222 43172 15256
rect 43206 15222 43262 15256
rect 43296 15222 43352 15256
rect 43386 15222 43442 15256
rect 43476 15222 43532 15256
rect 43566 15222 43627 15256
rect 42933 15194 43627 15222
rect 42933 15166 43020 15194
rect 43054 15166 43120 15194
rect 42933 15132 42992 15166
rect 43054 15160 43082 15166
rect 43026 15132 43082 15160
rect 43116 15160 43120 15166
rect 43154 15166 43220 15194
rect 43154 15160 43172 15166
rect 43116 15132 43172 15160
rect 43206 15160 43220 15166
rect 43254 15166 43320 15194
rect 43354 15166 43420 15194
rect 43454 15166 43520 15194
rect 43554 15166 43627 15194
rect 43254 15160 43262 15166
rect 43206 15132 43262 15160
rect 43296 15160 43320 15166
rect 43386 15160 43420 15166
rect 43476 15160 43520 15166
rect 43296 15132 43352 15160
rect 43386 15132 43442 15160
rect 43476 15132 43532 15160
rect 43566 15132 43627 15166
rect 42933 15073 43627 15132
rect 43689 15735 43708 15769
rect 43742 15735 43761 15769
rect 43689 15679 43761 15735
rect 43689 15645 43708 15679
rect 43742 15645 43761 15679
rect 43689 15589 43761 15645
rect 43689 15555 43708 15589
rect 43742 15555 43761 15589
rect 43689 15499 43761 15555
rect 43689 15465 43708 15499
rect 43742 15465 43761 15499
rect 43689 15409 43761 15465
rect 43689 15375 43708 15409
rect 43742 15375 43761 15409
rect 43689 15319 43761 15375
rect 43689 15285 43708 15319
rect 43742 15285 43761 15319
rect 43689 15229 43761 15285
rect 43689 15195 43708 15229
rect 43742 15195 43761 15229
rect 43689 15139 43761 15195
rect 43689 15105 43708 15139
rect 43742 15105 43761 15139
rect 42799 15034 42818 15068
rect 42852 15034 42871 15068
rect 42799 15020 42871 15034
rect 43689 15049 43761 15105
rect 43689 15020 43708 15049
rect 42703 15015 43708 15020
rect 43742 15020 43761 15049
rect 43825 15858 44095 15914
rect 45185 15948 45284 15965
rect 45185 15914 45216 15948
rect 45250 15914 45284 15948
rect 43825 15824 43856 15858
rect 43890 15824 44029 15858
rect 44063 15824 44095 15858
rect 43825 15768 44095 15824
rect 43825 15734 43856 15768
rect 43890 15734 44029 15768
rect 44063 15734 44095 15768
rect 43825 15678 44095 15734
rect 43825 15644 43856 15678
rect 43890 15644 44029 15678
rect 44063 15644 44095 15678
rect 43825 15588 44095 15644
rect 43825 15554 43856 15588
rect 43890 15554 44029 15588
rect 44063 15554 44095 15588
rect 43825 15498 44095 15554
rect 43825 15464 43856 15498
rect 43890 15464 44029 15498
rect 44063 15464 44095 15498
rect 43825 15408 44095 15464
rect 43825 15374 43856 15408
rect 43890 15374 44029 15408
rect 44063 15374 44095 15408
rect 43825 15318 44095 15374
rect 43825 15284 43856 15318
rect 43890 15284 44029 15318
rect 44063 15284 44095 15318
rect 43825 15228 44095 15284
rect 43825 15194 43856 15228
rect 43890 15194 44029 15228
rect 44063 15194 44095 15228
rect 43825 15138 44095 15194
rect 43825 15104 43856 15138
rect 43890 15104 44029 15138
rect 44063 15104 44095 15138
rect 43825 15048 44095 15104
rect 43825 15020 43856 15048
rect 43742 15015 43856 15020
rect 42703 15014 43856 15015
rect 43890 15014 44029 15048
rect 44063 15020 44095 15048
rect 44159 15882 45121 15901
rect 44159 15848 44270 15882
rect 44304 15848 44360 15882
rect 44394 15848 44450 15882
rect 44484 15848 44540 15882
rect 44574 15848 44630 15882
rect 44664 15848 44720 15882
rect 44754 15848 44810 15882
rect 44844 15848 44900 15882
rect 44934 15848 44990 15882
rect 45024 15848 45121 15882
rect 44159 15829 45121 15848
rect 44159 15788 44231 15829
rect 44159 15754 44178 15788
rect 44212 15754 44231 15788
rect 45049 15769 45121 15829
rect 44159 15698 44231 15754
rect 44159 15664 44178 15698
rect 44212 15664 44231 15698
rect 44159 15608 44231 15664
rect 44159 15574 44178 15608
rect 44212 15574 44231 15608
rect 44159 15518 44231 15574
rect 44159 15484 44178 15518
rect 44212 15484 44231 15518
rect 44159 15428 44231 15484
rect 44159 15394 44178 15428
rect 44212 15394 44231 15428
rect 44159 15338 44231 15394
rect 44159 15304 44178 15338
rect 44212 15304 44231 15338
rect 44159 15248 44231 15304
rect 44159 15214 44178 15248
rect 44212 15214 44231 15248
rect 44159 15158 44231 15214
rect 44159 15124 44178 15158
rect 44212 15124 44231 15158
rect 44159 15068 44231 15124
rect 44293 15706 44987 15767
rect 44293 15672 44352 15706
rect 44386 15694 44442 15706
rect 44414 15672 44442 15694
rect 44476 15694 44532 15706
rect 44476 15672 44480 15694
rect 44293 15660 44380 15672
rect 44414 15660 44480 15672
rect 44514 15672 44532 15694
rect 44566 15694 44622 15706
rect 44566 15672 44580 15694
rect 44514 15660 44580 15672
rect 44614 15672 44622 15694
rect 44656 15694 44712 15706
rect 44746 15694 44802 15706
rect 44836 15694 44892 15706
rect 44656 15672 44680 15694
rect 44746 15672 44780 15694
rect 44836 15672 44880 15694
rect 44926 15672 44987 15706
rect 44614 15660 44680 15672
rect 44714 15660 44780 15672
rect 44814 15660 44880 15672
rect 44914 15660 44987 15672
rect 44293 15616 44987 15660
rect 44293 15582 44352 15616
rect 44386 15594 44442 15616
rect 44414 15582 44442 15594
rect 44476 15594 44532 15616
rect 44476 15582 44480 15594
rect 44293 15560 44380 15582
rect 44414 15560 44480 15582
rect 44514 15582 44532 15594
rect 44566 15594 44622 15616
rect 44566 15582 44580 15594
rect 44514 15560 44580 15582
rect 44614 15582 44622 15594
rect 44656 15594 44712 15616
rect 44746 15594 44802 15616
rect 44836 15594 44892 15616
rect 44656 15582 44680 15594
rect 44746 15582 44780 15594
rect 44836 15582 44880 15594
rect 44926 15582 44987 15616
rect 44614 15560 44680 15582
rect 44714 15560 44780 15582
rect 44814 15560 44880 15582
rect 44914 15560 44987 15582
rect 44293 15526 44987 15560
rect 44293 15492 44352 15526
rect 44386 15494 44442 15526
rect 44414 15492 44442 15494
rect 44476 15494 44532 15526
rect 44476 15492 44480 15494
rect 44293 15460 44380 15492
rect 44414 15460 44480 15492
rect 44514 15492 44532 15494
rect 44566 15494 44622 15526
rect 44566 15492 44580 15494
rect 44514 15460 44580 15492
rect 44614 15492 44622 15494
rect 44656 15494 44712 15526
rect 44746 15494 44802 15526
rect 44836 15494 44892 15526
rect 44656 15492 44680 15494
rect 44746 15492 44780 15494
rect 44836 15492 44880 15494
rect 44926 15492 44987 15526
rect 44614 15460 44680 15492
rect 44714 15460 44780 15492
rect 44814 15460 44880 15492
rect 44914 15460 44987 15492
rect 44293 15436 44987 15460
rect 44293 15402 44352 15436
rect 44386 15402 44442 15436
rect 44476 15402 44532 15436
rect 44566 15402 44622 15436
rect 44656 15402 44712 15436
rect 44746 15402 44802 15436
rect 44836 15402 44892 15436
rect 44926 15402 44987 15436
rect 44293 15394 44987 15402
rect 44293 15360 44380 15394
rect 44414 15360 44480 15394
rect 44514 15360 44580 15394
rect 44614 15360 44680 15394
rect 44714 15360 44780 15394
rect 44814 15360 44880 15394
rect 44914 15360 44987 15394
rect 44293 15346 44987 15360
rect 44293 15312 44352 15346
rect 44386 15312 44442 15346
rect 44476 15312 44532 15346
rect 44566 15312 44622 15346
rect 44656 15312 44712 15346
rect 44746 15312 44802 15346
rect 44836 15312 44892 15346
rect 44926 15312 44987 15346
rect 44293 15294 44987 15312
rect 44293 15260 44380 15294
rect 44414 15260 44480 15294
rect 44514 15260 44580 15294
rect 44614 15260 44680 15294
rect 44714 15260 44780 15294
rect 44814 15260 44880 15294
rect 44914 15260 44987 15294
rect 44293 15256 44987 15260
rect 44293 15222 44352 15256
rect 44386 15222 44442 15256
rect 44476 15222 44532 15256
rect 44566 15222 44622 15256
rect 44656 15222 44712 15256
rect 44746 15222 44802 15256
rect 44836 15222 44892 15256
rect 44926 15222 44987 15256
rect 44293 15194 44987 15222
rect 44293 15166 44380 15194
rect 44414 15166 44480 15194
rect 44293 15132 44352 15166
rect 44414 15160 44442 15166
rect 44386 15132 44442 15160
rect 44476 15160 44480 15166
rect 44514 15166 44580 15194
rect 44514 15160 44532 15166
rect 44476 15132 44532 15160
rect 44566 15160 44580 15166
rect 44614 15166 44680 15194
rect 44714 15166 44780 15194
rect 44814 15166 44880 15194
rect 44914 15166 44987 15194
rect 44614 15160 44622 15166
rect 44566 15132 44622 15160
rect 44656 15160 44680 15166
rect 44746 15160 44780 15166
rect 44836 15160 44880 15166
rect 44656 15132 44712 15160
rect 44746 15132 44802 15160
rect 44836 15132 44892 15160
rect 44926 15132 44987 15166
rect 44293 15073 44987 15132
rect 45049 15735 45068 15769
rect 45102 15735 45121 15769
rect 45049 15679 45121 15735
rect 45049 15645 45068 15679
rect 45102 15645 45121 15679
rect 45049 15589 45121 15645
rect 45049 15555 45068 15589
rect 45102 15555 45121 15589
rect 45049 15499 45121 15555
rect 45049 15465 45068 15499
rect 45102 15465 45121 15499
rect 45049 15409 45121 15465
rect 45049 15375 45068 15409
rect 45102 15375 45121 15409
rect 45049 15319 45121 15375
rect 45049 15285 45068 15319
rect 45102 15285 45121 15319
rect 45049 15229 45121 15285
rect 45049 15195 45068 15229
rect 45102 15195 45121 15229
rect 45049 15139 45121 15195
rect 45049 15105 45068 15139
rect 45102 15105 45121 15139
rect 44159 15034 44178 15068
rect 44212 15034 44231 15068
rect 44159 15020 44231 15034
rect 45049 15049 45121 15105
rect 45049 15020 45068 15049
rect 44063 15015 45068 15020
rect 45102 15020 45121 15049
rect 45185 15858 45284 15914
rect 45185 15824 45216 15858
rect 45250 15824 45284 15858
rect 45185 15768 45284 15824
rect 47011 18499 47045 18561
rect 46593 15847 46627 15909
rect 47383 18555 47479 18589
rect 47739 18555 47835 18589
rect 47383 18493 47417 18555
rect 47570 18550 47590 18555
rect 47630 18550 47650 18555
rect 47570 18530 47650 18550
rect 47801 18493 47835 18555
rect 47383 16527 47417 16589
rect 47801 16527 47835 16589
rect 47383 16493 47479 16527
rect 47739 16493 47835 16527
rect 47011 15847 47045 15909
rect 46593 15813 46689 15847
rect 46949 15813 47045 15847
rect 45185 15734 45216 15768
rect 45250 15734 45284 15768
rect 45185 15678 45284 15734
rect 45185 15644 45216 15678
rect 45250 15644 45284 15678
rect 45185 15588 45284 15644
rect 45185 15554 45216 15588
rect 45250 15554 45284 15588
rect 45185 15498 45284 15554
rect 45185 15464 45216 15498
rect 45250 15464 45284 15498
rect 45185 15408 45284 15464
rect 45185 15374 45216 15408
rect 45250 15374 45284 15408
rect 45185 15318 45284 15374
rect 45185 15284 45216 15318
rect 45250 15284 45284 15318
rect 45185 15228 45284 15284
rect 45185 15194 45216 15228
rect 45250 15194 45284 15228
rect 45185 15138 45284 15194
rect 45185 15104 45216 15138
rect 45250 15104 45284 15138
rect 45185 15048 45284 15104
rect 45185 15020 45216 15048
rect 45102 15015 45216 15020
rect 44063 15014 45216 15015
rect 45250 15020 45284 15048
rect 45250 15014 45290 15020
rect 41270 14992 45290 15014
rect 41270 14958 41516 14992
rect 41550 14958 41606 14992
rect 41640 14958 41696 14992
rect 41730 14958 41786 14992
rect 41820 14958 41876 14992
rect 41910 14958 41966 14992
rect 42000 14958 42056 14992
rect 42090 14958 42146 14992
rect 42180 14958 42236 14992
rect 42270 14958 42876 14992
rect 42910 14958 42966 14992
rect 43000 14958 43056 14992
rect 43090 14958 43146 14992
rect 43180 14958 43236 14992
rect 43270 14958 43326 14992
rect 43360 14958 43416 14992
rect 43450 14958 43506 14992
rect 43540 14958 43596 14992
rect 43630 14958 44236 14992
rect 44270 14958 44326 14992
rect 44360 14958 44416 14992
rect 44450 14958 44506 14992
rect 44540 14958 44596 14992
rect 44630 14958 44686 14992
rect 44720 14958 44776 14992
rect 44810 14958 44866 14992
rect 44900 14958 44956 14992
rect 44990 14958 45290 14992
rect 41270 14924 41309 14958
rect 41343 14924 42496 14958
rect 42530 14924 42669 14958
rect 42703 14924 43856 14958
rect 43890 14924 44029 14958
rect 44063 14924 45216 14958
rect 45250 14924 45290 14958
rect 41270 14868 45290 14924
rect 41270 14834 41309 14868
rect 41343 14845 42496 14868
rect 41343 14834 41410 14845
rect 41270 14811 41410 14834
rect 41444 14811 41500 14845
rect 41534 14811 41590 14845
rect 41624 14811 41680 14845
rect 41714 14811 41770 14845
rect 41804 14811 41860 14845
rect 41894 14811 41950 14845
rect 41984 14811 42040 14845
rect 42074 14811 42130 14845
rect 42164 14811 42220 14845
rect 42254 14811 42310 14845
rect 42344 14811 42400 14845
rect 42434 14834 42496 14845
rect 42530 14834 42669 14868
rect 42703 14845 43856 14868
rect 42703 14834 42770 14845
rect 42434 14811 42770 14834
rect 42804 14811 42860 14845
rect 42894 14811 42950 14845
rect 42984 14811 43040 14845
rect 43074 14811 43130 14845
rect 43164 14811 43220 14845
rect 43254 14811 43310 14845
rect 43344 14811 43400 14845
rect 43434 14811 43490 14845
rect 43524 14811 43580 14845
rect 43614 14811 43670 14845
rect 43704 14811 43760 14845
rect 43794 14834 43856 14845
rect 43890 14834 44029 14868
rect 44063 14845 45216 14868
rect 44063 14834 44130 14845
rect 43794 14811 44130 14834
rect 44164 14811 44220 14845
rect 44254 14811 44310 14845
rect 44344 14811 44400 14845
rect 44434 14811 44490 14845
rect 44524 14811 44580 14845
rect 44614 14811 44670 14845
rect 44704 14811 44760 14845
rect 44794 14811 44850 14845
rect 44884 14811 44940 14845
rect 44974 14811 45030 14845
rect 45064 14811 45120 14845
rect 45154 14834 45216 14845
rect 45250 14834 45290 14868
rect 45154 14811 45290 14834
rect 41270 14770 45290 14811
rect 41403 14571 41499 14605
rect 45057 14571 45153 14605
rect 41403 14509 41437 14571
rect 45119 14509 45153 14571
rect 41403 14187 41437 14249
rect 45119 14187 45153 14249
rect 41403 14153 41499 14187
rect 45057 14153 45153 14187
rect 41170 13850 41230 13870
rect 41170 13820 41180 13850
rect 41080 13810 41180 13820
rect 41220 13810 41230 13850
rect 41080 13800 41230 13810
rect 41080 13760 41100 13800
rect 41140 13760 41230 13800
rect 41080 13750 41230 13760
rect 41080 13740 41180 13750
rect 41170 13710 41180 13740
rect 41220 13710 41230 13750
rect 41170 13690 41230 13710
rect 43250 13850 43310 13870
rect 43250 13810 43260 13850
rect 43300 13810 43310 13850
rect 43250 13750 43310 13810
rect 43250 13710 43260 13750
rect 43300 13710 43310 13750
rect 43250 13690 43310 13710
rect 45330 13860 45470 13870
rect 45330 13850 45550 13860
rect 45330 13810 45340 13850
rect 45380 13810 45420 13850
rect 45460 13840 45550 13850
rect 45460 13810 45490 13840
rect 45330 13800 45490 13810
rect 45530 13800 45550 13840
rect 45330 13760 45550 13800
rect 45330 13750 45490 13760
rect 45330 13710 45340 13750
rect 45380 13710 45420 13750
rect 45460 13720 45490 13750
rect 45530 13720 45550 13760
rect 45460 13710 45550 13720
rect 45330 13700 45550 13710
rect 45330 13690 45470 13700
rect 41180 13650 41220 13690
rect 43260 13650 43300 13690
rect 41160 13630 41240 13650
rect 41160 13590 41180 13630
rect 41220 13590 41240 13630
rect 41160 13570 41240 13590
rect 41320 13630 41400 13650
rect 41320 13590 41340 13630
rect 41380 13590 41400 13630
rect 41320 13570 41400 13590
rect 41480 13630 41560 13650
rect 41480 13590 41500 13630
rect 41540 13590 41560 13630
rect 41480 13570 41560 13590
rect 41640 13630 41720 13650
rect 41640 13590 41660 13630
rect 41700 13590 41720 13630
rect 41640 13570 41720 13590
rect 41800 13630 41880 13650
rect 41800 13590 41820 13630
rect 41860 13590 41880 13630
rect 41800 13570 41880 13590
rect 41960 13630 42040 13650
rect 41960 13590 41980 13630
rect 42020 13590 42040 13630
rect 41960 13570 42040 13590
rect 42120 13630 42200 13650
rect 42120 13590 42140 13630
rect 42180 13590 42200 13630
rect 42120 13570 42200 13590
rect 42280 13630 42360 13650
rect 42280 13590 42300 13630
rect 42340 13590 42360 13630
rect 42280 13570 42360 13590
rect 42440 13630 42520 13650
rect 42440 13590 42460 13630
rect 42500 13590 42520 13630
rect 42440 13570 42520 13590
rect 42600 13630 42680 13650
rect 42600 13590 42620 13630
rect 42660 13590 42680 13630
rect 42600 13570 42680 13590
rect 42760 13630 42840 13650
rect 42760 13590 42780 13630
rect 42820 13590 42840 13630
rect 42760 13570 42840 13590
rect 42920 13630 43000 13650
rect 42920 13590 42940 13630
rect 42980 13590 43000 13630
rect 42920 13570 43000 13590
rect 43080 13630 43160 13650
rect 43080 13590 43100 13630
rect 43140 13590 43160 13630
rect 43080 13570 43160 13590
rect 43240 13630 43320 13650
rect 43240 13590 43260 13630
rect 43300 13590 43320 13630
rect 43240 13570 43320 13590
rect 43400 13630 43480 13650
rect 43400 13590 43420 13630
rect 43460 13590 43480 13630
rect 43400 13570 43480 13590
rect 43560 13630 43640 13650
rect 43560 13590 43580 13630
rect 43620 13590 43640 13630
rect 43560 13570 43640 13590
rect 43720 13630 43800 13650
rect 43720 13590 43740 13630
rect 43780 13590 43800 13630
rect 43720 13570 43800 13590
rect 43880 13630 43960 13650
rect 43880 13590 43900 13630
rect 43940 13590 43960 13630
rect 43880 13570 43960 13590
rect 44040 13630 44120 13650
rect 44040 13590 44060 13630
rect 44100 13590 44120 13630
rect 44040 13570 44120 13590
rect 44200 13630 44280 13650
rect 44200 13590 44220 13630
rect 44260 13590 44280 13630
rect 44200 13570 44280 13590
rect 44360 13630 44440 13650
rect 44360 13590 44380 13630
rect 44420 13590 44440 13630
rect 44360 13570 44440 13590
rect 44520 13630 44600 13650
rect 44520 13590 44540 13630
rect 44580 13590 44600 13630
rect 44520 13570 44600 13590
rect 44680 13630 44760 13650
rect 44680 13590 44700 13630
rect 44740 13590 44760 13630
rect 44680 13570 44760 13590
rect 44840 13630 44920 13650
rect 44840 13590 44860 13630
rect 44900 13590 44920 13630
rect 44840 13570 44920 13590
rect 45000 13630 45080 13650
rect 45000 13590 45020 13630
rect 45060 13590 45080 13630
rect 45000 13570 45080 13590
rect 45160 13630 45240 13650
rect 45160 13590 45180 13630
rect 45220 13590 45240 13630
rect 45160 13570 45240 13590
rect 41900 13360 41980 13380
rect 41900 13320 41920 13360
rect 41960 13320 41980 13360
rect 41900 13260 41980 13320
rect 44580 13360 44660 13380
rect 44580 13320 44600 13360
rect 44640 13320 44660 13360
rect 44580 13260 44660 13320
rect 40750 13240 40810 13260
rect 40750 13200 40760 13240
rect 40800 13200 40810 13240
rect 40750 13140 40810 13200
rect 40750 13100 40760 13140
rect 40800 13100 40810 13140
rect 40750 13040 40810 13100
rect 40750 13000 40760 13040
rect 40800 13000 40810 13040
rect 40750 12940 40810 13000
rect 40750 12900 40760 12940
rect 40800 12900 40810 12940
rect 40750 12840 40810 12900
rect 40750 12800 40760 12840
rect 40800 12800 40810 12840
rect 40750 12780 40810 12800
rect 41830 13240 42050 13260
rect 41830 13200 41840 13240
rect 41880 13200 41920 13240
rect 41960 13200 42000 13240
rect 42040 13200 42050 13240
rect 41830 13140 42050 13200
rect 41830 13100 41840 13140
rect 41880 13100 41920 13140
rect 41960 13100 42000 13140
rect 42040 13100 42050 13140
rect 41830 13040 42050 13100
rect 41830 13000 41840 13040
rect 41880 13000 41920 13040
rect 41960 13000 42000 13040
rect 42040 13000 42050 13040
rect 41830 12940 42050 13000
rect 41830 12900 41840 12940
rect 41880 12900 41920 12940
rect 41960 12900 42000 12940
rect 42040 12900 42050 12940
rect 41830 12840 42050 12900
rect 41830 12800 41840 12840
rect 41880 12800 41920 12840
rect 41960 12800 42000 12840
rect 42040 12800 42050 12840
rect 41830 12780 42050 12800
rect 43070 13240 43130 13260
rect 43070 13200 43080 13240
rect 43120 13200 43130 13240
rect 43070 13140 43130 13200
rect 43070 13100 43080 13140
rect 43120 13100 43130 13140
rect 43070 13040 43130 13100
rect 43070 13000 43080 13040
rect 43120 13000 43130 13040
rect 43070 12940 43130 13000
rect 43070 12900 43080 12940
rect 43120 12900 43130 12940
rect 43070 12840 43130 12900
rect 43070 12800 43080 12840
rect 43120 12800 43130 12840
rect 40740 12760 40820 12780
rect 40740 12720 40760 12760
rect 40800 12720 40820 12760
rect 43070 12750 43130 12800
rect 40740 12700 40820 12720
rect 40920 12720 41000 12740
rect 40920 12680 40940 12720
rect 40980 12680 41000 12720
rect 40920 12660 41000 12680
rect 41160 12720 41240 12740
rect 41160 12680 41180 12720
rect 41220 12680 41240 12720
rect 41160 12660 41240 12680
rect 41400 12720 41480 12740
rect 41400 12680 41420 12720
rect 41460 12680 41480 12720
rect 41400 12660 41480 12680
rect 41640 12720 41720 12740
rect 41640 12680 41660 12720
rect 41700 12680 41720 12720
rect 41640 12660 41720 12680
rect 42280 12720 42360 12740
rect 42280 12680 42300 12720
rect 42340 12680 42360 12720
rect 42280 12660 42360 12680
rect 42520 12720 42600 12740
rect 42520 12680 42540 12720
rect 42580 12680 42600 12720
rect 42520 12660 42600 12680
rect 42760 12720 42840 12740
rect 42760 12680 42780 12720
rect 42820 12680 42840 12720
rect 43070 12710 43080 12750
rect 43120 12710 43130 12750
rect 43070 12690 43130 12710
rect 43430 13240 43490 13260
rect 43430 13200 43440 13240
rect 43480 13200 43490 13240
rect 43430 13140 43490 13200
rect 43430 13100 43440 13140
rect 43480 13100 43490 13140
rect 43430 13040 43490 13100
rect 43430 13000 43440 13040
rect 43480 13000 43490 13040
rect 43430 12940 43490 13000
rect 43430 12900 43440 12940
rect 43480 12900 43490 12940
rect 43430 12840 43490 12900
rect 43430 12800 43440 12840
rect 43480 12800 43490 12840
rect 43430 12750 43490 12800
rect 44510 13240 44730 13260
rect 44510 13200 44520 13240
rect 44560 13200 44600 13240
rect 44640 13200 44680 13240
rect 44720 13200 44730 13240
rect 44510 13140 44730 13200
rect 44510 13100 44520 13140
rect 44560 13100 44600 13140
rect 44640 13100 44680 13140
rect 44720 13100 44730 13140
rect 44510 13040 44730 13100
rect 44510 13000 44520 13040
rect 44560 13000 44600 13040
rect 44640 13000 44680 13040
rect 44720 13000 44730 13040
rect 44510 12940 44730 13000
rect 44510 12900 44520 12940
rect 44560 12900 44600 12940
rect 44640 12900 44680 12940
rect 44720 12900 44730 12940
rect 44510 12840 44730 12900
rect 44510 12800 44520 12840
rect 44560 12800 44600 12840
rect 44640 12800 44680 12840
rect 44720 12800 44730 12840
rect 44510 12780 44730 12800
rect 45750 13240 45810 13260
rect 45750 13200 45760 13240
rect 45800 13200 45810 13240
rect 45750 13140 45810 13200
rect 45750 13100 45760 13140
rect 45800 13100 45810 13140
rect 45750 13040 45810 13100
rect 45750 13000 45760 13040
rect 45800 13000 45810 13040
rect 45750 12940 45810 13000
rect 45750 12900 45760 12940
rect 45800 12900 45810 12940
rect 45750 12840 45810 12900
rect 45750 12800 45760 12840
rect 45800 12800 45810 12840
rect 45750 12780 45810 12800
rect 43430 12710 43440 12750
rect 43480 12710 43490 12750
rect 43430 12690 43490 12710
rect 43720 12720 43800 12740
rect 42760 12660 42840 12680
rect 43720 12680 43740 12720
rect 43780 12680 43800 12720
rect 43720 12660 43800 12680
rect 43960 12720 44040 12740
rect 43960 12680 43980 12720
rect 44020 12680 44040 12720
rect 43960 12660 44040 12680
rect 44200 12720 44280 12740
rect 44200 12680 44220 12720
rect 44260 12680 44280 12720
rect 44200 12660 44280 12680
rect 44840 12720 44920 12740
rect 44840 12680 44860 12720
rect 44900 12680 44920 12720
rect 44840 12660 44920 12680
rect 45080 12720 45160 12740
rect 45080 12680 45100 12720
rect 45140 12680 45160 12720
rect 45080 12660 45160 12680
rect 45320 12720 45400 12740
rect 45320 12680 45340 12720
rect 45380 12680 45400 12720
rect 45320 12660 45400 12680
rect 45560 12720 45640 12740
rect 45560 12680 45580 12720
rect 45620 12680 45640 12720
rect 45560 12660 45640 12680
rect 41431 12342 41489 12360
rect 41431 12308 41443 12342
rect 41477 12308 41489 12342
rect 41431 12290 41489 12308
rect 41791 12342 41849 12360
rect 41791 12308 41803 12342
rect 41837 12308 41849 12342
rect 41791 12290 41849 12308
rect 41911 12342 41969 12360
rect 41911 12308 41923 12342
rect 41957 12308 41969 12342
rect 41911 12290 41969 12308
rect 42271 12342 42329 12360
rect 42271 12308 42283 12342
rect 42317 12308 42329 12342
rect 42271 12290 42329 12308
rect 42391 12342 42449 12360
rect 42391 12308 42403 12342
rect 42437 12308 42449 12342
rect 44111 12342 44169 12360
rect 42391 12290 42449 12308
rect 42800 12320 42880 12340
rect 42800 12280 42820 12320
rect 42860 12280 42880 12320
rect 41370 12230 41430 12250
rect 41370 12190 41380 12230
rect 41420 12190 41430 12230
rect 41370 12170 41430 12190
rect 41490 12230 41550 12250
rect 41490 12190 41500 12230
rect 41540 12190 41550 12230
rect 41490 12170 41550 12190
rect 41610 12230 41670 12250
rect 41610 12190 41620 12230
rect 41660 12190 41670 12230
rect 41610 12170 41670 12190
rect 41730 12230 41790 12250
rect 41730 12190 41740 12230
rect 41780 12190 41790 12230
rect 41730 12170 41790 12190
rect 41850 12230 41910 12250
rect 41850 12190 41860 12230
rect 41900 12190 41910 12230
rect 41850 12170 41910 12190
rect 41970 12230 42030 12250
rect 41970 12190 41980 12230
rect 42020 12190 42030 12230
rect 41970 12170 42030 12190
rect 42090 12230 42150 12250
rect 42090 12190 42100 12230
rect 42140 12190 42150 12230
rect 42090 12170 42150 12190
rect 42210 12230 42270 12250
rect 42210 12190 42220 12230
rect 42260 12190 42270 12230
rect 42210 12170 42270 12190
rect 42330 12230 42390 12250
rect 42330 12190 42340 12230
rect 42380 12190 42390 12230
rect 42330 12170 42390 12190
rect 42450 12230 42510 12250
rect 42450 12190 42460 12230
rect 42500 12190 42510 12230
rect 42450 12170 42510 12190
rect 42570 12230 42630 12250
rect 42570 12190 42580 12230
rect 42620 12190 42630 12230
rect 42570 12170 42630 12190
rect 42800 12240 42880 12280
rect 42800 12200 42820 12240
rect 42860 12200 42880 12240
rect 42800 12160 42880 12200
rect 41532 12112 41590 12130
rect 41532 12078 41544 12112
rect 41578 12078 41590 12112
rect 41532 12060 41590 12078
rect 41690 12112 41748 12130
rect 41690 12078 41702 12112
rect 41736 12078 41748 12112
rect 41690 12060 41748 12078
rect 42014 12112 42072 12130
rect 42014 12078 42026 12112
rect 42060 12078 42072 12112
rect 42014 12060 42072 12078
rect 42168 12112 42226 12130
rect 42168 12078 42180 12112
rect 42214 12078 42226 12112
rect 42168 12060 42226 12078
rect 42492 12112 42550 12130
rect 42492 12078 42504 12112
rect 42538 12078 42550 12112
rect 42800 12120 42820 12160
rect 42860 12120 42880 12160
rect 42800 12100 42880 12120
rect 43680 12320 43760 12340
rect 43680 12280 43700 12320
rect 43740 12280 43760 12320
rect 44111 12308 44123 12342
rect 44157 12308 44169 12342
rect 44111 12290 44169 12308
rect 44231 12342 44289 12360
rect 44231 12308 44243 12342
rect 44277 12308 44289 12342
rect 44231 12290 44289 12308
rect 44591 12342 44649 12360
rect 44591 12308 44603 12342
rect 44637 12308 44649 12342
rect 44591 12290 44649 12308
rect 44711 12342 44769 12360
rect 44711 12308 44723 12342
rect 44757 12308 44769 12342
rect 44711 12290 44769 12308
rect 45071 12342 45129 12360
rect 45071 12308 45083 12342
rect 45117 12308 45129 12342
rect 45071 12290 45129 12308
rect 43680 12240 43760 12280
rect 43680 12200 43700 12240
rect 43740 12200 43760 12240
rect 43680 12160 43760 12200
rect 43930 12230 43990 12250
rect 43930 12190 43940 12230
rect 43980 12190 43990 12230
rect 43930 12170 43990 12190
rect 44050 12230 44110 12250
rect 44050 12190 44060 12230
rect 44100 12190 44110 12230
rect 44050 12170 44110 12190
rect 44170 12230 44230 12250
rect 44170 12190 44180 12230
rect 44220 12190 44230 12230
rect 44170 12170 44230 12190
rect 44290 12230 44350 12250
rect 44290 12190 44300 12230
rect 44340 12190 44350 12230
rect 44290 12170 44350 12190
rect 44410 12230 44470 12250
rect 44410 12190 44420 12230
rect 44460 12190 44470 12230
rect 44410 12170 44470 12190
rect 44530 12230 44590 12250
rect 44530 12190 44540 12230
rect 44580 12190 44590 12230
rect 44530 12170 44590 12190
rect 44650 12230 44710 12250
rect 44650 12190 44660 12230
rect 44700 12190 44710 12230
rect 44650 12170 44710 12190
rect 44770 12230 44830 12250
rect 44770 12190 44780 12230
rect 44820 12190 44830 12230
rect 44770 12170 44830 12190
rect 44890 12230 44950 12250
rect 44890 12190 44900 12230
rect 44940 12190 44950 12230
rect 44890 12170 44950 12190
rect 45010 12230 45070 12250
rect 45010 12190 45020 12230
rect 45060 12190 45070 12230
rect 45010 12170 45070 12190
rect 45130 12230 45190 12250
rect 45130 12190 45140 12230
rect 45180 12190 45190 12230
rect 45130 12170 45190 12190
rect 43680 12120 43700 12160
rect 43740 12120 43760 12160
rect 43680 12100 43760 12120
rect 44010 12112 44068 12130
rect 42492 12060 42550 12078
rect 44010 12078 44022 12112
rect 44056 12078 44068 12112
rect 44010 12060 44068 12078
rect 44334 12112 44392 12130
rect 44334 12078 44346 12112
rect 44380 12078 44392 12112
rect 44334 12060 44392 12078
rect 44488 12112 44546 12130
rect 44488 12078 44500 12112
rect 44534 12078 44546 12112
rect 44488 12060 44546 12078
rect 44812 12112 44870 12130
rect 44812 12078 44824 12112
rect 44858 12078 44870 12112
rect 44812 12060 44870 12078
rect 44970 12112 45028 12130
rect 44970 12078 44982 12112
rect 45016 12078 45028 12112
rect 44970 12060 45028 12078
rect 40710 11520 40770 11540
rect 40710 11480 40720 11520
rect 40760 11480 40770 11520
rect 40710 11460 40770 11480
rect 40880 11510 40960 11530
rect 40880 11470 40900 11510
rect 40940 11470 40960 11510
rect 40880 11450 40960 11470
rect 41370 11510 41430 11530
rect 41370 11470 41380 11510
rect 41420 11470 41430 11510
rect 41370 11450 41430 11470
rect 41600 11510 41680 11530
rect 41600 11470 41620 11510
rect 41660 11470 41680 11510
rect 41600 11450 41680 11470
rect 42090 11510 42150 11530
rect 42090 11470 42100 11510
rect 42140 11470 42150 11510
rect 42090 11450 42150 11470
rect 42320 11510 42400 11530
rect 42320 11470 42340 11510
rect 42380 11470 42400 11510
rect 42320 11450 42400 11470
rect 42750 11510 42810 11530
rect 42750 11470 42760 11510
rect 42800 11470 42810 11510
rect 42750 11450 42810 11470
rect 43750 11510 43810 11530
rect 43750 11470 43760 11510
rect 43800 11470 43810 11510
rect 43750 11450 43810 11470
rect 44160 11510 44240 11530
rect 44160 11470 44180 11510
rect 44220 11470 44240 11510
rect 44160 11450 44240 11470
rect 44410 11510 44470 11530
rect 44410 11470 44420 11510
rect 44460 11470 44470 11510
rect 44410 11450 44470 11470
rect 44880 11510 44960 11530
rect 44880 11470 44900 11510
rect 44940 11470 44960 11510
rect 44880 11450 44960 11470
rect 45130 11510 45190 11530
rect 45130 11470 45140 11510
rect 45180 11470 45190 11510
rect 45130 11450 45190 11470
rect 45600 11510 45680 11530
rect 45600 11470 45620 11510
rect 45660 11470 45680 11510
rect 45600 11450 45680 11470
rect 45790 11520 45850 11540
rect 45790 11480 45800 11520
rect 45840 11480 45850 11520
rect 45790 11460 45850 11480
rect 40450 11390 40590 11410
rect 40450 11350 40460 11390
rect 40500 11350 40540 11390
rect 40580 11350 40590 11390
rect 40450 11290 40590 11350
rect 40450 11250 40460 11290
rect 40500 11250 40540 11290
rect 40580 11250 40590 11290
rect 40450 11230 40590 11250
rect 40650 11390 40710 11410
rect 40650 11350 40660 11390
rect 40700 11350 40710 11390
rect 40650 11290 40710 11350
rect 40650 11250 40660 11290
rect 40700 11250 40710 11290
rect 40650 11230 40710 11250
rect 40770 11390 40830 11410
rect 40770 11350 40780 11390
rect 40820 11350 40830 11390
rect 40770 11290 40830 11350
rect 40770 11250 40780 11290
rect 40820 11250 40830 11290
rect 40770 11230 40830 11250
rect 40890 11390 40950 11410
rect 40890 11350 40900 11390
rect 40940 11350 40950 11390
rect 40890 11290 40950 11350
rect 40890 11250 40900 11290
rect 40940 11250 40950 11290
rect 40890 11230 40950 11250
rect 41010 11390 41070 11410
rect 41010 11350 41020 11390
rect 41060 11350 41070 11390
rect 41010 11290 41070 11350
rect 41010 11250 41020 11290
rect 41060 11250 41070 11290
rect 41010 11230 41070 11250
rect 41130 11390 41190 11410
rect 41130 11350 41140 11390
rect 41180 11350 41190 11390
rect 41130 11290 41190 11350
rect 41130 11250 41140 11290
rect 41180 11250 41190 11290
rect 41130 11230 41190 11250
rect 41250 11390 41310 11410
rect 41250 11350 41260 11390
rect 41300 11350 41310 11390
rect 41250 11290 41310 11350
rect 41250 11250 41260 11290
rect 41300 11250 41310 11290
rect 41250 11230 41310 11250
rect 41370 11390 41430 11410
rect 41370 11350 41380 11390
rect 41420 11350 41430 11390
rect 41370 11290 41430 11350
rect 41370 11250 41380 11290
rect 41420 11250 41430 11290
rect 41370 11230 41430 11250
rect 41490 11390 41550 11410
rect 41490 11350 41500 11390
rect 41540 11350 41550 11390
rect 41490 11290 41550 11350
rect 41490 11250 41500 11290
rect 41540 11250 41550 11290
rect 41490 11230 41550 11250
rect 41610 11390 41670 11410
rect 41610 11350 41620 11390
rect 41660 11350 41670 11390
rect 41610 11290 41670 11350
rect 41610 11250 41620 11290
rect 41660 11250 41670 11290
rect 41610 11230 41670 11250
rect 41730 11390 41790 11410
rect 41730 11350 41740 11390
rect 41780 11350 41790 11390
rect 41730 11290 41790 11350
rect 41730 11250 41740 11290
rect 41780 11250 41790 11290
rect 41730 11230 41790 11250
rect 41850 11390 41910 11410
rect 41850 11350 41860 11390
rect 41900 11350 41910 11390
rect 41850 11290 41910 11350
rect 41850 11250 41860 11290
rect 41900 11250 41910 11290
rect 41850 11230 41910 11250
rect 41970 11390 42030 11410
rect 41970 11350 41980 11390
rect 42020 11350 42030 11390
rect 41970 11290 42030 11350
rect 41970 11250 41980 11290
rect 42020 11250 42030 11290
rect 41970 11230 42030 11250
rect 42090 11390 42150 11410
rect 42090 11350 42100 11390
rect 42140 11350 42150 11390
rect 42090 11290 42150 11350
rect 42090 11250 42100 11290
rect 42140 11250 42150 11290
rect 42090 11230 42150 11250
rect 42210 11390 42270 11410
rect 42210 11350 42220 11390
rect 42260 11350 42270 11390
rect 42210 11290 42270 11350
rect 42210 11250 42220 11290
rect 42260 11250 42270 11290
rect 42210 11230 42270 11250
rect 42330 11390 42390 11410
rect 42330 11350 42340 11390
rect 42380 11350 42390 11390
rect 42330 11290 42390 11350
rect 42330 11250 42340 11290
rect 42380 11250 42390 11290
rect 42330 11230 42390 11250
rect 42450 11390 42510 11410
rect 42450 11350 42460 11390
rect 42500 11350 42510 11390
rect 42450 11290 42510 11350
rect 42450 11250 42460 11290
rect 42500 11250 42510 11290
rect 42450 11230 42510 11250
rect 42570 11390 42630 11410
rect 42570 11350 42580 11390
rect 42620 11350 42630 11390
rect 42570 11290 42630 11350
rect 42570 11250 42580 11290
rect 42620 11250 42630 11290
rect 42570 11230 42630 11250
rect 42690 11390 42750 11410
rect 42690 11350 42700 11390
rect 42740 11350 42750 11390
rect 42690 11290 42750 11350
rect 42690 11250 42700 11290
rect 42740 11250 42750 11290
rect 42690 11230 42750 11250
rect 42810 11390 42870 11410
rect 42810 11350 42820 11390
rect 42860 11350 42870 11390
rect 42810 11290 42870 11350
rect 42810 11250 42820 11290
rect 42860 11250 42870 11290
rect 42810 11230 42870 11250
rect 42930 11390 43070 11410
rect 42930 11350 42940 11390
rect 42980 11350 43020 11390
rect 43060 11350 43070 11390
rect 42930 11290 43070 11350
rect 42930 11250 42940 11290
rect 42980 11250 43020 11290
rect 43060 11250 43070 11290
rect 42930 11230 43070 11250
rect 43490 11390 43630 11410
rect 43490 11350 43500 11390
rect 43540 11350 43580 11390
rect 43620 11350 43630 11390
rect 43490 11290 43630 11350
rect 43490 11250 43500 11290
rect 43540 11250 43580 11290
rect 43620 11250 43630 11290
rect 43490 11230 43630 11250
rect 43690 11390 43750 11410
rect 43690 11350 43700 11390
rect 43740 11350 43750 11390
rect 43690 11290 43750 11350
rect 43690 11250 43700 11290
rect 43740 11250 43750 11290
rect 43690 11230 43750 11250
rect 43810 11390 43870 11410
rect 43810 11350 43820 11390
rect 43860 11350 43870 11390
rect 43810 11290 43870 11350
rect 43810 11250 43820 11290
rect 43860 11250 43870 11290
rect 43810 11230 43870 11250
rect 43930 11390 43990 11410
rect 43930 11350 43940 11390
rect 43980 11350 43990 11390
rect 43930 11290 43990 11350
rect 43930 11250 43940 11290
rect 43980 11250 43990 11290
rect 43930 11230 43990 11250
rect 44050 11390 44110 11410
rect 44050 11350 44060 11390
rect 44100 11350 44110 11390
rect 44050 11290 44110 11350
rect 44050 11250 44060 11290
rect 44100 11250 44110 11290
rect 44050 11230 44110 11250
rect 44170 11390 44230 11410
rect 44170 11350 44180 11390
rect 44220 11350 44230 11390
rect 44170 11290 44230 11350
rect 44170 11250 44180 11290
rect 44220 11250 44230 11290
rect 44170 11230 44230 11250
rect 44290 11390 44350 11410
rect 44290 11350 44300 11390
rect 44340 11350 44350 11390
rect 44290 11290 44350 11350
rect 44290 11250 44300 11290
rect 44340 11250 44350 11290
rect 44290 11230 44350 11250
rect 44410 11390 44470 11410
rect 44410 11350 44420 11390
rect 44460 11350 44470 11390
rect 44410 11290 44470 11350
rect 44410 11250 44420 11290
rect 44460 11250 44470 11290
rect 44410 11230 44470 11250
rect 44530 11390 44590 11410
rect 44530 11350 44540 11390
rect 44580 11350 44590 11390
rect 44530 11290 44590 11350
rect 44530 11250 44540 11290
rect 44580 11250 44590 11290
rect 44530 11230 44590 11250
rect 44650 11390 44710 11410
rect 44650 11350 44660 11390
rect 44700 11350 44710 11390
rect 44650 11290 44710 11350
rect 44650 11250 44660 11290
rect 44700 11250 44710 11290
rect 44650 11230 44710 11250
rect 44770 11390 44830 11410
rect 44770 11350 44780 11390
rect 44820 11350 44830 11390
rect 44770 11290 44830 11350
rect 44770 11250 44780 11290
rect 44820 11250 44830 11290
rect 44770 11230 44830 11250
rect 44890 11390 44950 11410
rect 44890 11350 44900 11390
rect 44940 11350 44950 11390
rect 44890 11290 44950 11350
rect 44890 11250 44900 11290
rect 44940 11250 44950 11290
rect 44890 11230 44950 11250
rect 45010 11390 45070 11410
rect 45010 11350 45020 11390
rect 45060 11350 45070 11390
rect 45010 11290 45070 11350
rect 45010 11250 45020 11290
rect 45060 11250 45070 11290
rect 45010 11230 45070 11250
rect 45130 11390 45190 11410
rect 45130 11350 45140 11390
rect 45180 11350 45190 11390
rect 45130 11290 45190 11350
rect 45130 11250 45140 11290
rect 45180 11250 45190 11290
rect 45130 11230 45190 11250
rect 45250 11390 45310 11410
rect 45250 11350 45260 11390
rect 45300 11350 45310 11390
rect 45250 11290 45310 11350
rect 45250 11250 45260 11290
rect 45300 11250 45310 11290
rect 45250 11230 45310 11250
rect 45370 11390 45430 11410
rect 45370 11350 45380 11390
rect 45420 11350 45430 11390
rect 45370 11290 45430 11350
rect 45370 11250 45380 11290
rect 45420 11250 45430 11290
rect 45370 11230 45430 11250
rect 45490 11390 45550 11410
rect 45490 11350 45500 11390
rect 45540 11350 45550 11390
rect 45490 11290 45550 11350
rect 45490 11250 45500 11290
rect 45540 11250 45550 11290
rect 45490 11230 45550 11250
rect 45610 11390 45670 11410
rect 45610 11350 45620 11390
rect 45660 11350 45670 11390
rect 45610 11290 45670 11350
rect 45610 11250 45620 11290
rect 45660 11250 45670 11290
rect 45610 11230 45670 11250
rect 45730 11390 45790 11410
rect 45730 11350 45740 11390
rect 45780 11350 45790 11390
rect 45730 11290 45790 11350
rect 45730 11250 45740 11290
rect 45780 11250 45790 11290
rect 45730 11230 45790 11250
rect 45850 11390 45910 11410
rect 45850 11350 45860 11390
rect 45900 11350 45910 11390
rect 45850 11290 45910 11350
rect 45850 11250 45860 11290
rect 45900 11250 45910 11290
rect 45850 11230 45910 11250
rect 45970 11390 46110 11410
rect 45970 11350 45980 11390
rect 46020 11350 46060 11390
rect 46100 11350 46110 11390
rect 45970 11290 46110 11350
rect 45970 11250 45980 11290
rect 46020 11250 46060 11290
rect 46100 11250 46110 11290
rect 45970 11230 46110 11250
rect 40530 11170 40590 11190
rect 40530 11130 40540 11170
rect 40580 11130 40590 11170
rect 40530 11110 40590 11130
rect 42930 11170 42990 11190
rect 42930 11130 42940 11170
rect 42980 11130 42990 11170
rect 42930 11110 42990 11130
rect 43570 11170 43630 11190
rect 43570 11130 43580 11170
rect 43620 11130 43630 11170
rect 43570 11110 43630 11130
rect 45970 11170 46030 11190
rect 45970 11130 45980 11170
rect 46020 11130 46030 11170
rect 45970 11110 46030 11130
rect 41900 10350 41970 10370
rect 41900 10310 41910 10350
rect 41950 10310 41970 10350
rect 41900 10290 41970 10310
rect 42070 10350 42150 10370
rect 42070 10310 42090 10350
rect 42130 10310 42150 10350
rect 42070 10290 42150 10310
rect 42250 10350 42330 10370
rect 42250 10310 42270 10350
rect 42310 10310 42330 10350
rect 42250 10290 42330 10310
rect 42430 10350 42510 10370
rect 42430 10310 42450 10350
rect 42490 10310 42510 10350
rect 42430 10290 42510 10310
rect 42610 10350 42690 10370
rect 42610 10310 42630 10350
rect 42670 10310 42690 10350
rect 42610 10290 42690 10310
rect 42790 10350 42870 10370
rect 42790 10310 42810 10350
rect 42850 10310 42870 10350
rect 42790 10290 42870 10310
rect 42970 10350 43050 10370
rect 42970 10310 42990 10350
rect 43030 10310 43050 10350
rect 42970 10290 43050 10310
rect 43150 10350 43220 10370
rect 43150 10310 43170 10350
rect 43210 10310 43220 10350
rect 43150 10290 43220 10310
rect 43340 10350 43410 10370
rect 43340 10310 43350 10350
rect 43390 10310 43410 10350
rect 43340 10290 43410 10310
rect 43510 10350 43590 10370
rect 43510 10310 43530 10350
rect 43570 10310 43590 10350
rect 43510 10290 43590 10310
rect 43690 10350 43770 10370
rect 43690 10310 43710 10350
rect 43750 10310 43770 10350
rect 43690 10290 43770 10310
rect 43870 10350 43950 10370
rect 43870 10310 43890 10350
rect 43930 10310 43950 10350
rect 43870 10290 43950 10310
rect 44050 10350 44130 10370
rect 44050 10310 44070 10350
rect 44110 10310 44130 10350
rect 44050 10290 44130 10310
rect 44230 10350 44310 10370
rect 44230 10310 44250 10350
rect 44290 10310 44310 10350
rect 44230 10290 44310 10310
rect 44410 10350 44490 10370
rect 44410 10310 44430 10350
rect 44470 10310 44490 10350
rect 44410 10290 44490 10310
rect 44590 10350 44660 10370
rect 44590 10310 44610 10350
rect 44650 10310 44660 10350
rect 44590 10290 44660 10310
rect 41550 10230 41690 10250
rect 41550 10190 41560 10230
rect 41600 10190 41640 10230
rect 41680 10190 41690 10230
rect 41550 10130 41690 10190
rect 41550 10090 41560 10130
rect 41600 10090 41640 10130
rect 41680 10090 41690 10130
rect 41550 10030 41690 10090
rect 41550 9990 41560 10030
rect 41600 9990 41640 10030
rect 41680 9990 41690 10030
rect 41550 9930 41690 9990
rect 41550 9890 41560 9930
rect 41600 9890 41640 9930
rect 41680 9890 41690 9930
rect 41550 9830 41690 9890
rect 41550 9790 41560 9830
rect 41600 9790 41640 9830
rect 41680 9790 41690 9830
rect 41550 9730 41690 9790
rect 41550 9690 41560 9730
rect 41600 9690 41640 9730
rect 41680 9690 41690 9730
rect 41550 9670 41690 9690
rect 41810 10230 41870 10250
rect 41810 10190 41820 10230
rect 41860 10190 41870 10230
rect 41810 10130 41870 10190
rect 41810 10090 41820 10130
rect 41860 10090 41870 10130
rect 41810 10030 41870 10090
rect 41810 9990 41820 10030
rect 41860 9990 41870 10030
rect 41810 9930 41870 9990
rect 41810 9890 41820 9930
rect 41860 9890 41870 9930
rect 41810 9830 41870 9890
rect 41810 9790 41820 9830
rect 41860 9790 41870 9830
rect 41810 9730 41870 9790
rect 41810 9690 41820 9730
rect 41860 9690 41870 9730
rect 41810 9670 41870 9690
rect 41990 10230 42050 10250
rect 41990 10190 42000 10230
rect 42040 10190 42050 10230
rect 41990 10130 42050 10190
rect 41990 10090 42000 10130
rect 42040 10090 42050 10130
rect 41990 10030 42050 10090
rect 41990 9990 42000 10030
rect 42040 9990 42050 10030
rect 41990 9930 42050 9990
rect 41990 9890 42000 9930
rect 42040 9890 42050 9930
rect 41990 9830 42050 9890
rect 41990 9790 42000 9830
rect 42040 9790 42050 9830
rect 41990 9730 42050 9790
rect 41990 9690 42000 9730
rect 42040 9690 42050 9730
rect 41990 9670 42050 9690
rect 42170 10230 42230 10250
rect 42170 10190 42180 10230
rect 42220 10190 42230 10230
rect 42170 10130 42230 10190
rect 42170 10090 42180 10130
rect 42220 10090 42230 10130
rect 42170 10030 42230 10090
rect 42170 9990 42180 10030
rect 42220 9990 42230 10030
rect 42170 9930 42230 9990
rect 42170 9890 42180 9930
rect 42220 9890 42230 9930
rect 42170 9830 42230 9890
rect 42170 9790 42180 9830
rect 42220 9790 42230 9830
rect 42170 9730 42230 9790
rect 42170 9690 42180 9730
rect 42220 9690 42230 9730
rect 42170 9670 42230 9690
rect 42350 10230 42410 10250
rect 42350 10190 42360 10230
rect 42400 10190 42410 10230
rect 42350 10130 42410 10190
rect 42350 10090 42360 10130
rect 42400 10090 42410 10130
rect 42350 10030 42410 10090
rect 42350 9990 42360 10030
rect 42400 9990 42410 10030
rect 42350 9930 42410 9990
rect 42350 9890 42360 9930
rect 42400 9890 42410 9930
rect 42350 9830 42410 9890
rect 42350 9790 42360 9830
rect 42400 9790 42410 9830
rect 42350 9730 42410 9790
rect 42350 9690 42360 9730
rect 42400 9690 42410 9730
rect 42350 9670 42410 9690
rect 42530 10230 42590 10250
rect 42530 10190 42540 10230
rect 42580 10190 42590 10230
rect 42530 10130 42590 10190
rect 42530 10090 42540 10130
rect 42580 10090 42590 10130
rect 42530 10030 42590 10090
rect 42530 9990 42540 10030
rect 42580 9990 42590 10030
rect 42530 9930 42590 9990
rect 42530 9890 42540 9930
rect 42580 9890 42590 9930
rect 42530 9830 42590 9890
rect 42530 9790 42540 9830
rect 42580 9790 42590 9830
rect 42530 9730 42590 9790
rect 42530 9690 42540 9730
rect 42580 9690 42590 9730
rect 42530 9670 42590 9690
rect 42710 10230 42770 10250
rect 42710 10190 42720 10230
rect 42760 10190 42770 10230
rect 42710 10130 42770 10190
rect 42710 10090 42720 10130
rect 42760 10090 42770 10130
rect 42710 10030 42770 10090
rect 42710 9990 42720 10030
rect 42760 9990 42770 10030
rect 42710 9930 42770 9990
rect 42710 9890 42720 9930
rect 42760 9890 42770 9930
rect 42710 9830 42770 9890
rect 42710 9790 42720 9830
rect 42760 9790 42770 9830
rect 42710 9730 42770 9790
rect 42710 9690 42720 9730
rect 42760 9690 42770 9730
rect 42710 9670 42770 9690
rect 42890 10230 42950 10250
rect 42890 10190 42900 10230
rect 42940 10190 42950 10230
rect 42890 10130 42950 10190
rect 42890 10090 42900 10130
rect 42940 10090 42950 10130
rect 42890 10030 42950 10090
rect 42890 9990 42900 10030
rect 42940 9990 42950 10030
rect 42890 9930 42950 9990
rect 42890 9890 42900 9930
rect 42940 9890 42950 9930
rect 42890 9830 42950 9890
rect 42890 9790 42900 9830
rect 42940 9790 42950 9830
rect 42890 9730 42950 9790
rect 42890 9690 42900 9730
rect 42940 9690 42950 9730
rect 42890 9670 42950 9690
rect 43070 10230 43130 10250
rect 43070 10190 43080 10230
rect 43120 10190 43130 10230
rect 43070 10130 43130 10190
rect 43070 10090 43080 10130
rect 43120 10090 43130 10130
rect 43070 10030 43130 10090
rect 43070 9990 43080 10030
rect 43120 9990 43130 10030
rect 43070 9930 43130 9990
rect 43070 9890 43080 9930
rect 43120 9890 43130 9930
rect 43070 9830 43130 9890
rect 43070 9790 43080 9830
rect 43120 9790 43130 9830
rect 43070 9730 43130 9790
rect 43070 9690 43080 9730
rect 43120 9690 43130 9730
rect 43070 9670 43130 9690
rect 43250 10230 43310 10250
rect 43250 10190 43260 10230
rect 43300 10190 43310 10230
rect 43250 10130 43310 10190
rect 43250 10090 43260 10130
rect 43300 10090 43310 10130
rect 43250 10030 43310 10090
rect 43250 9990 43260 10030
rect 43300 9990 43310 10030
rect 43250 9930 43310 9990
rect 43250 9890 43260 9930
rect 43300 9890 43310 9930
rect 43250 9830 43310 9890
rect 43250 9790 43260 9830
rect 43300 9790 43310 9830
rect 43250 9730 43310 9790
rect 43250 9690 43260 9730
rect 43300 9690 43310 9730
rect 43250 9670 43310 9690
rect 43430 10230 43490 10250
rect 43430 10190 43440 10230
rect 43480 10190 43490 10230
rect 43430 10130 43490 10190
rect 43430 10090 43440 10130
rect 43480 10090 43490 10130
rect 43430 10030 43490 10090
rect 43430 9990 43440 10030
rect 43480 9990 43490 10030
rect 43430 9930 43490 9990
rect 43430 9890 43440 9930
rect 43480 9890 43490 9930
rect 43430 9830 43490 9890
rect 43430 9790 43440 9830
rect 43480 9790 43490 9830
rect 43430 9730 43490 9790
rect 43430 9690 43440 9730
rect 43480 9690 43490 9730
rect 43430 9670 43490 9690
rect 43610 10230 43670 10250
rect 43610 10190 43620 10230
rect 43660 10190 43670 10230
rect 43610 10130 43670 10190
rect 43610 10090 43620 10130
rect 43660 10090 43670 10130
rect 43610 10030 43670 10090
rect 43610 9990 43620 10030
rect 43660 9990 43670 10030
rect 43610 9930 43670 9990
rect 43610 9890 43620 9930
rect 43660 9890 43670 9930
rect 43610 9830 43670 9890
rect 43610 9790 43620 9830
rect 43660 9790 43670 9830
rect 43610 9730 43670 9790
rect 43610 9690 43620 9730
rect 43660 9690 43670 9730
rect 43610 9670 43670 9690
rect 43790 10230 43850 10250
rect 43790 10190 43800 10230
rect 43840 10190 43850 10230
rect 43790 10130 43850 10190
rect 43790 10090 43800 10130
rect 43840 10090 43850 10130
rect 43790 10030 43850 10090
rect 43790 9990 43800 10030
rect 43840 9990 43850 10030
rect 43790 9930 43850 9990
rect 43790 9890 43800 9930
rect 43840 9890 43850 9930
rect 43790 9830 43850 9890
rect 43790 9790 43800 9830
rect 43840 9790 43850 9830
rect 43790 9730 43850 9790
rect 43790 9690 43800 9730
rect 43840 9690 43850 9730
rect 43790 9670 43850 9690
rect 43970 10230 44030 10250
rect 43970 10190 43980 10230
rect 44020 10190 44030 10230
rect 43970 10130 44030 10190
rect 43970 10090 43980 10130
rect 44020 10090 44030 10130
rect 43970 10030 44030 10090
rect 43970 9990 43980 10030
rect 44020 9990 44030 10030
rect 43970 9930 44030 9990
rect 43970 9890 43980 9930
rect 44020 9890 44030 9930
rect 43970 9830 44030 9890
rect 43970 9790 43980 9830
rect 44020 9790 44030 9830
rect 43970 9730 44030 9790
rect 43970 9690 43980 9730
rect 44020 9690 44030 9730
rect 43970 9670 44030 9690
rect 44150 10230 44210 10250
rect 44150 10190 44160 10230
rect 44200 10190 44210 10230
rect 44150 10130 44210 10190
rect 44150 10090 44160 10130
rect 44200 10090 44210 10130
rect 44150 10030 44210 10090
rect 44150 9990 44160 10030
rect 44200 9990 44210 10030
rect 44150 9930 44210 9990
rect 44150 9890 44160 9930
rect 44200 9890 44210 9930
rect 44150 9830 44210 9890
rect 44150 9790 44160 9830
rect 44200 9790 44210 9830
rect 44150 9730 44210 9790
rect 44150 9690 44160 9730
rect 44200 9690 44210 9730
rect 44150 9670 44210 9690
rect 44330 10230 44390 10250
rect 44330 10190 44340 10230
rect 44380 10190 44390 10230
rect 44330 10130 44390 10190
rect 44330 10090 44340 10130
rect 44380 10090 44390 10130
rect 44330 10030 44390 10090
rect 44330 9990 44340 10030
rect 44380 9990 44390 10030
rect 44330 9930 44390 9990
rect 44330 9890 44340 9930
rect 44380 9890 44390 9930
rect 44330 9830 44390 9890
rect 44330 9790 44340 9830
rect 44380 9790 44390 9830
rect 44330 9730 44390 9790
rect 44330 9690 44340 9730
rect 44380 9690 44390 9730
rect 44330 9670 44390 9690
rect 44510 10230 44570 10250
rect 44510 10190 44520 10230
rect 44560 10190 44570 10230
rect 44510 10130 44570 10190
rect 44510 10090 44520 10130
rect 44560 10090 44570 10130
rect 44510 10030 44570 10090
rect 44510 9990 44520 10030
rect 44560 9990 44570 10030
rect 44510 9930 44570 9990
rect 44510 9890 44520 9930
rect 44560 9890 44570 9930
rect 44510 9830 44570 9890
rect 44510 9790 44520 9830
rect 44560 9790 44570 9830
rect 44510 9730 44570 9790
rect 44510 9690 44520 9730
rect 44560 9690 44570 9730
rect 44510 9670 44570 9690
rect 44690 10230 44750 10250
rect 44690 10190 44700 10230
rect 44740 10190 44750 10230
rect 44690 10130 44750 10190
rect 44690 10090 44700 10130
rect 44740 10090 44750 10130
rect 44690 10030 44750 10090
rect 44690 9990 44700 10030
rect 44740 9990 44750 10030
rect 44690 9930 44750 9990
rect 44690 9890 44700 9930
rect 44740 9890 44750 9930
rect 44690 9830 44750 9890
rect 44690 9790 44700 9830
rect 44740 9790 44750 9830
rect 44690 9730 44750 9790
rect 44690 9690 44700 9730
rect 44740 9690 44750 9730
rect 44690 9670 44750 9690
rect 44870 10230 45010 10250
rect 44870 10190 44880 10230
rect 44920 10190 44960 10230
rect 45000 10190 45010 10230
rect 44870 10130 45010 10190
rect 44870 10090 44880 10130
rect 44920 10090 44960 10130
rect 45000 10090 45010 10130
rect 45590 10150 45670 10170
rect 45590 10110 45610 10150
rect 45650 10110 45670 10150
rect 45590 10090 45670 10110
rect 45710 10150 45790 10170
rect 45710 10110 45730 10150
rect 45770 10110 45790 10150
rect 45710 10090 45790 10110
rect 45830 10150 45910 10170
rect 45830 10110 45850 10150
rect 45890 10110 45910 10150
rect 45830 10090 45910 10110
rect 44870 10030 45010 10090
rect 44870 9990 44880 10030
rect 44920 9990 44960 10030
rect 45000 9990 45010 10030
rect 44870 9930 45010 9990
rect 44870 9890 44880 9930
rect 44920 9890 44960 9930
rect 45000 9890 45010 9930
rect 44870 9830 45010 9890
rect 45410 10030 45560 10050
rect 45410 9990 45420 10030
rect 45460 9990 45510 10030
rect 45550 9990 45560 10030
rect 45410 9930 45560 9990
rect 45410 9890 45420 9930
rect 45460 9890 45510 9930
rect 45550 9890 45560 9930
rect 45410 9870 45560 9890
rect 45610 10030 45670 10050
rect 45610 9990 45620 10030
rect 45660 9990 45670 10030
rect 45610 9930 45670 9990
rect 45610 9890 45620 9930
rect 45660 9890 45670 9930
rect 45610 9870 45670 9890
rect 45720 10030 45780 10050
rect 45720 9990 45730 10030
rect 45770 9990 45780 10030
rect 45720 9930 45780 9990
rect 45720 9890 45730 9930
rect 45770 9890 45780 9930
rect 45720 9870 45780 9890
rect 45830 10030 45890 10050
rect 45830 9990 45840 10030
rect 45880 9990 45890 10030
rect 45830 9930 45890 9990
rect 45830 9890 45840 9930
rect 45880 9890 45890 9930
rect 45830 9870 45890 9890
rect 45940 10030 46080 10050
rect 45940 9990 45950 10030
rect 45990 9990 46030 10030
rect 46070 9990 46080 10030
rect 45940 9930 46080 9990
rect 45940 9890 45950 9930
rect 45990 9890 46030 9930
rect 46070 9890 46080 9930
rect 45940 9870 46080 9890
rect 44870 9790 44880 9830
rect 44920 9790 44960 9830
rect 45000 9790 45010 9830
rect 44870 9730 45010 9790
rect 45490 9810 45570 9830
rect 45490 9770 45510 9810
rect 45550 9770 45570 9810
rect 45490 9750 45570 9770
rect 45710 9810 45790 9830
rect 45710 9770 45730 9810
rect 45770 9770 45790 9810
rect 45710 9750 45790 9770
rect 45940 9810 46000 9830
rect 45940 9770 45950 9810
rect 45990 9770 46000 9810
rect 45940 9750 46000 9770
rect 44870 9690 44880 9730
rect 44920 9690 44960 9730
rect 45000 9690 45010 9730
rect 44870 9670 45010 9690
rect 41640 9630 41680 9670
rect 42000 9630 42040 9670
rect 42360 9630 42400 9670
rect 42720 9630 42760 9670
rect 43080 9630 43120 9670
rect 43440 9630 43480 9670
rect 43800 9630 43840 9670
rect 44160 9630 44200 9670
rect 44520 9630 44560 9670
rect 44880 9630 44920 9670
rect 41620 9610 41700 9630
rect 41620 9570 41640 9610
rect 41680 9570 41700 9610
rect 41620 9550 41700 9570
rect 41980 9610 42060 9630
rect 41980 9570 42000 9610
rect 42040 9570 42060 9610
rect 41980 9550 42060 9570
rect 42340 9610 42420 9630
rect 42340 9570 42360 9610
rect 42400 9570 42420 9610
rect 42340 9550 42420 9570
rect 42700 9610 42780 9630
rect 42700 9570 42720 9610
rect 42760 9570 42780 9610
rect 42700 9550 42780 9570
rect 43060 9610 43140 9630
rect 43060 9570 43080 9610
rect 43120 9570 43140 9610
rect 43060 9550 43140 9570
rect 43420 9610 43500 9630
rect 43420 9570 43440 9610
rect 43480 9570 43500 9610
rect 43420 9550 43500 9570
rect 43780 9610 43860 9630
rect 43780 9570 43800 9610
rect 43840 9570 43860 9610
rect 43780 9550 43860 9570
rect 44140 9610 44220 9630
rect 44140 9570 44160 9610
rect 44200 9570 44220 9610
rect 44140 9550 44220 9570
rect 44500 9610 44580 9630
rect 44500 9570 44520 9610
rect 44560 9570 44580 9610
rect 44500 9550 44580 9570
rect 44860 9610 44940 9630
rect 44860 9570 44880 9610
rect 44920 9570 44940 9610
rect 44860 9550 44940 9570
rect 41806 9342 41864 9360
rect 41806 9308 41818 9342
rect 41852 9308 41864 9342
rect 41806 9290 41864 9308
rect 41916 9342 41974 9360
rect 41916 9308 41928 9342
rect 41962 9308 41974 9342
rect 41916 9290 41974 9308
rect 42026 9342 42084 9360
rect 42026 9308 42038 9342
rect 42072 9308 42084 9342
rect 42026 9290 42084 9308
rect 42136 9342 42194 9360
rect 42136 9308 42148 9342
rect 42182 9308 42194 9342
rect 42136 9290 42194 9308
rect 42246 9342 42304 9360
rect 42246 9308 42258 9342
rect 42292 9308 42304 9342
rect 42246 9290 42304 9308
rect 42356 9342 42414 9360
rect 42356 9308 42368 9342
rect 42402 9308 42414 9342
rect 42356 9290 42414 9308
rect 42466 9342 42524 9360
rect 42466 9308 42478 9342
rect 42512 9308 42524 9342
rect 42466 9290 42524 9308
rect 42576 9342 42634 9360
rect 42576 9308 42588 9342
rect 42622 9308 42634 9342
rect 42576 9290 42634 9308
rect 42686 9342 42744 9360
rect 42686 9308 42698 9342
rect 42732 9308 42744 9342
rect 42686 9290 42744 9308
rect 42796 9342 42854 9360
rect 42796 9308 42808 9342
rect 42842 9308 42854 9342
rect 42796 9290 42854 9308
rect 43706 9342 43764 9360
rect 43706 9308 43718 9342
rect 43752 9308 43764 9342
rect 43706 9290 43764 9308
rect 43816 9342 43874 9360
rect 43816 9308 43828 9342
rect 43862 9308 43874 9342
rect 43816 9290 43874 9308
rect 43926 9342 43984 9360
rect 43926 9308 43938 9342
rect 43972 9308 43984 9342
rect 43926 9290 43984 9308
rect 44036 9342 44094 9360
rect 44036 9308 44048 9342
rect 44082 9308 44094 9342
rect 44036 9290 44094 9308
rect 44146 9342 44204 9360
rect 44146 9308 44158 9342
rect 44192 9308 44204 9342
rect 44146 9290 44204 9308
rect 44256 9342 44314 9360
rect 44256 9308 44268 9342
rect 44302 9308 44314 9342
rect 44256 9290 44314 9308
rect 44366 9342 44424 9360
rect 44366 9308 44378 9342
rect 44412 9308 44424 9342
rect 44366 9290 44424 9308
rect 44476 9342 44534 9360
rect 44476 9308 44488 9342
rect 44522 9308 44534 9342
rect 44476 9290 44534 9308
rect 44586 9342 44644 9360
rect 44586 9308 44598 9342
rect 44632 9308 44644 9342
rect 44586 9290 44644 9308
rect 44696 9342 44754 9360
rect 44696 9308 44708 9342
rect 44742 9308 44754 9342
rect 44696 9290 44754 9308
rect 41560 9230 41700 9250
rect 41560 9190 41570 9230
rect 41610 9190 41650 9230
rect 41690 9190 41700 9230
rect 41560 9130 41700 9190
rect 41560 9090 41570 9130
rect 41610 9090 41650 9130
rect 41690 9090 41700 9130
rect 41560 9070 41700 9090
rect 41750 9230 41810 9250
rect 41750 9190 41760 9230
rect 41800 9190 41810 9230
rect 41750 9130 41810 9190
rect 41750 9090 41760 9130
rect 41800 9090 41810 9130
rect 41750 9070 41810 9090
rect 41860 9230 41920 9250
rect 41860 9190 41870 9230
rect 41910 9190 41920 9230
rect 41860 9130 41920 9190
rect 41860 9090 41870 9130
rect 41910 9090 41920 9130
rect 41860 9070 41920 9090
rect 41970 9230 42030 9250
rect 41970 9190 41980 9230
rect 42020 9190 42030 9230
rect 41970 9130 42030 9190
rect 41970 9090 41980 9130
rect 42020 9090 42030 9130
rect 41970 9070 42030 9090
rect 42080 9230 42140 9250
rect 42080 9190 42090 9230
rect 42130 9190 42140 9230
rect 42080 9130 42140 9190
rect 42080 9090 42090 9130
rect 42130 9090 42140 9130
rect 42080 9070 42140 9090
rect 42190 9230 42250 9250
rect 42190 9190 42200 9230
rect 42240 9190 42250 9230
rect 42190 9130 42250 9190
rect 42190 9090 42200 9130
rect 42240 9090 42250 9130
rect 42190 9070 42250 9090
rect 42300 9230 42360 9250
rect 42300 9190 42310 9230
rect 42350 9190 42360 9230
rect 42300 9130 42360 9190
rect 42300 9090 42310 9130
rect 42350 9090 42360 9130
rect 42300 9070 42360 9090
rect 42410 9230 42470 9250
rect 42410 9190 42420 9230
rect 42460 9190 42470 9230
rect 42410 9130 42470 9190
rect 42410 9090 42420 9130
rect 42460 9090 42470 9130
rect 42410 9070 42470 9090
rect 42520 9230 42580 9250
rect 42520 9190 42530 9230
rect 42570 9190 42580 9230
rect 42520 9130 42580 9190
rect 42520 9090 42530 9130
rect 42570 9090 42580 9130
rect 42520 9070 42580 9090
rect 42630 9230 42690 9250
rect 42630 9190 42640 9230
rect 42680 9190 42690 9230
rect 42630 9130 42690 9190
rect 42630 9090 42640 9130
rect 42680 9090 42690 9130
rect 42630 9070 42690 9090
rect 42740 9230 42800 9250
rect 42740 9190 42750 9230
rect 42790 9190 42800 9230
rect 42740 9130 42800 9190
rect 42740 9090 42750 9130
rect 42790 9090 42800 9130
rect 42740 9070 42800 9090
rect 42850 9230 42910 9250
rect 42850 9190 42860 9230
rect 42900 9190 42910 9230
rect 42850 9130 42910 9190
rect 42850 9090 42860 9130
rect 42900 9090 42910 9130
rect 42850 9070 42910 9090
rect 42960 9230 43100 9250
rect 42960 9190 42970 9230
rect 43010 9190 43050 9230
rect 43090 9190 43100 9230
rect 42960 9130 43100 9190
rect 42960 9090 42970 9130
rect 43010 9090 43050 9130
rect 43090 9090 43100 9130
rect 42960 9070 43100 9090
rect 43460 9230 43600 9250
rect 43460 9190 43470 9230
rect 43510 9190 43550 9230
rect 43590 9190 43600 9230
rect 43460 9130 43600 9190
rect 43460 9090 43470 9130
rect 43510 9090 43550 9130
rect 43590 9090 43600 9130
rect 43460 9070 43600 9090
rect 43650 9230 43710 9250
rect 43650 9190 43660 9230
rect 43700 9190 43710 9230
rect 43650 9130 43710 9190
rect 43650 9090 43660 9130
rect 43700 9090 43710 9130
rect 43650 9070 43710 9090
rect 43760 9230 43820 9250
rect 43760 9190 43770 9230
rect 43810 9190 43820 9230
rect 43760 9130 43820 9190
rect 43760 9090 43770 9130
rect 43810 9090 43820 9130
rect 43760 9070 43820 9090
rect 43870 9230 43930 9250
rect 43870 9190 43880 9230
rect 43920 9190 43930 9230
rect 43870 9130 43930 9190
rect 43870 9090 43880 9130
rect 43920 9090 43930 9130
rect 43870 9070 43930 9090
rect 43980 9230 44040 9250
rect 43980 9190 43990 9230
rect 44030 9190 44040 9230
rect 43980 9130 44040 9190
rect 43980 9090 43990 9130
rect 44030 9090 44040 9130
rect 43980 9070 44040 9090
rect 44090 9230 44150 9250
rect 44090 9190 44100 9230
rect 44140 9190 44150 9230
rect 44090 9130 44150 9190
rect 44090 9090 44100 9130
rect 44140 9090 44150 9130
rect 44090 9070 44150 9090
rect 44200 9230 44260 9250
rect 44200 9190 44210 9230
rect 44250 9190 44260 9230
rect 44200 9130 44260 9190
rect 44200 9090 44210 9130
rect 44250 9090 44260 9130
rect 44200 9070 44260 9090
rect 44310 9230 44370 9250
rect 44310 9190 44320 9230
rect 44360 9190 44370 9230
rect 44310 9130 44370 9190
rect 44310 9090 44320 9130
rect 44360 9090 44370 9130
rect 44310 9070 44370 9090
rect 44420 9230 44480 9250
rect 44420 9190 44430 9230
rect 44470 9190 44480 9230
rect 44420 9130 44480 9190
rect 44420 9090 44430 9130
rect 44470 9090 44480 9130
rect 44420 9070 44480 9090
rect 44530 9230 44590 9250
rect 44530 9190 44540 9230
rect 44580 9190 44590 9230
rect 44530 9130 44590 9190
rect 44530 9090 44540 9130
rect 44580 9090 44590 9130
rect 44530 9070 44590 9090
rect 44640 9230 44700 9250
rect 44640 9190 44650 9230
rect 44690 9190 44700 9230
rect 44640 9130 44700 9190
rect 44640 9090 44650 9130
rect 44690 9090 44700 9130
rect 44640 9070 44700 9090
rect 44750 9230 44810 9250
rect 44750 9190 44760 9230
rect 44800 9190 44810 9230
rect 44750 9130 44810 9190
rect 44750 9090 44760 9130
rect 44800 9090 44810 9130
rect 44750 9070 44810 9090
rect 44860 9230 45000 9250
rect 44860 9190 44870 9230
rect 44910 9190 44950 9230
rect 44990 9190 45000 9230
rect 44860 9130 45000 9190
rect 44860 9090 44870 9130
rect 44910 9090 44950 9130
rect 44990 9090 45000 9130
rect 44860 9070 45000 9090
rect 41630 9010 41710 9030
rect 41630 8970 41650 9010
rect 41690 8970 41710 9010
rect 41630 8950 41710 8970
rect 42950 9010 43030 9030
rect 42950 8970 42970 9010
rect 43010 8970 43030 9010
rect 42950 8950 43030 8970
rect 43530 9010 43610 9030
rect 43530 8970 43550 9010
rect 43590 8970 43610 9010
rect 43530 8950 43610 8970
rect 44850 9010 44930 9030
rect 44850 8970 44870 9010
rect 44910 8970 44930 9010
rect 44850 8950 44930 8970
<< viali >>
rect 43260 19030 43300 19070
rect 43260 18950 43300 18990
rect 43260 18870 43300 18910
rect 39590 18595 39630 18600
rect 40700 18597 40740 18610
rect 38810 18589 38850 18590
rect 38810 18555 38850 18589
rect 38810 18550 38850 18555
rect 38776 18035 38882 18432
rect 38776 16650 38882 17047
rect 39590 18561 39630 18595
rect 39590 18560 39630 18561
rect 39590 18041 39628 18438
rect 39590 15080 39628 15477
rect 40700 18570 40740 18597
rect 40700 18050 40740 18440
rect 40370 16310 40410 16700
rect 41660 18392 41666 18414
rect 41666 18392 41694 18414
rect 41660 18380 41694 18392
rect 41760 18380 41794 18414
rect 41860 18380 41894 18414
rect 41960 18392 41992 18414
rect 41992 18392 41994 18414
rect 42060 18392 42082 18414
rect 42082 18392 42094 18414
rect 42160 18392 42172 18414
rect 42172 18392 42194 18414
rect 41960 18380 41994 18392
rect 42060 18380 42094 18392
rect 42160 18380 42194 18392
rect 41660 18302 41666 18314
rect 41666 18302 41694 18314
rect 41660 18280 41694 18302
rect 41760 18280 41794 18314
rect 41860 18280 41894 18314
rect 41960 18302 41992 18314
rect 41992 18302 41994 18314
rect 42060 18302 42082 18314
rect 42082 18302 42094 18314
rect 42160 18302 42172 18314
rect 42172 18302 42194 18314
rect 41960 18280 41994 18302
rect 42060 18280 42094 18302
rect 42160 18280 42194 18302
rect 41660 18212 41666 18214
rect 41666 18212 41694 18214
rect 41660 18180 41694 18212
rect 41760 18180 41794 18214
rect 41860 18180 41894 18214
rect 41960 18212 41992 18214
rect 41992 18212 41994 18214
rect 42060 18212 42082 18214
rect 42082 18212 42094 18214
rect 42160 18212 42172 18214
rect 42172 18212 42194 18214
rect 41960 18180 41994 18212
rect 42060 18180 42094 18212
rect 42160 18180 42194 18212
rect 41660 18080 41694 18114
rect 41760 18080 41794 18114
rect 41860 18080 41894 18114
rect 41960 18080 41994 18114
rect 42060 18080 42094 18114
rect 42160 18080 42194 18114
rect 41660 17980 41694 18014
rect 41760 17980 41794 18014
rect 41860 17980 41894 18014
rect 41960 17980 41994 18014
rect 42060 17980 42094 18014
rect 42160 17980 42194 18014
rect 41660 17886 41694 17914
rect 41660 17880 41666 17886
rect 41666 17880 41694 17886
rect 41760 17880 41794 17914
rect 41860 17880 41894 17914
rect 41960 17886 41994 17914
rect 42060 17886 42094 17914
rect 42160 17886 42194 17914
rect 41960 17880 41992 17886
rect 41992 17880 41994 17886
rect 42060 17880 42082 17886
rect 42082 17880 42094 17886
rect 42160 17880 42172 17886
rect 42172 17880 42194 17886
rect 43020 18392 43026 18414
rect 43026 18392 43054 18414
rect 43020 18380 43054 18392
rect 43120 18380 43154 18414
rect 43220 18380 43254 18414
rect 43320 18392 43352 18414
rect 43352 18392 43354 18414
rect 43420 18392 43442 18414
rect 43442 18392 43454 18414
rect 43520 18392 43532 18414
rect 43532 18392 43554 18414
rect 43320 18380 43354 18392
rect 43420 18380 43454 18392
rect 43520 18380 43554 18392
rect 43020 18302 43026 18314
rect 43026 18302 43054 18314
rect 43020 18280 43054 18302
rect 43120 18280 43154 18314
rect 43220 18280 43254 18314
rect 43320 18302 43352 18314
rect 43352 18302 43354 18314
rect 43420 18302 43442 18314
rect 43442 18302 43454 18314
rect 43520 18302 43532 18314
rect 43532 18302 43554 18314
rect 43320 18280 43354 18302
rect 43420 18280 43454 18302
rect 43520 18280 43554 18302
rect 43020 18212 43026 18214
rect 43026 18212 43054 18214
rect 43020 18180 43054 18212
rect 43120 18180 43154 18214
rect 43220 18180 43254 18214
rect 43320 18212 43352 18214
rect 43352 18212 43354 18214
rect 43420 18212 43442 18214
rect 43442 18212 43454 18214
rect 43520 18212 43532 18214
rect 43532 18212 43554 18214
rect 43320 18180 43354 18212
rect 43420 18180 43454 18212
rect 43520 18180 43554 18212
rect 43020 18080 43054 18114
rect 43120 18080 43154 18114
rect 43220 18080 43254 18114
rect 43320 18080 43354 18114
rect 43420 18080 43454 18114
rect 43520 18080 43554 18114
rect 43020 17980 43054 18014
rect 43120 17980 43154 18014
rect 43220 17980 43254 18014
rect 43320 17980 43354 18014
rect 43420 17980 43454 18014
rect 43520 17980 43554 18014
rect 43020 17886 43054 17914
rect 43020 17880 43026 17886
rect 43026 17880 43054 17886
rect 43120 17880 43154 17914
rect 43220 17880 43254 17914
rect 43320 17886 43354 17914
rect 43420 17886 43454 17914
rect 43520 17886 43554 17914
rect 43320 17880 43352 17886
rect 43352 17880 43354 17886
rect 43420 17880 43442 17886
rect 43442 17880 43454 17886
rect 43520 17880 43532 17886
rect 43532 17880 43554 17886
rect 44380 18392 44386 18414
rect 44386 18392 44414 18414
rect 44380 18380 44414 18392
rect 44480 18380 44514 18414
rect 44580 18380 44614 18414
rect 44680 18392 44712 18414
rect 44712 18392 44714 18414
rect 44780 18392 44802 18414
rect 44802 18392 44814 18414
rect 44880 18392 44892 18414
rect 44892 18392 44914 18414
rect 44680 18380 44714 18392
rect 44780 18380 44814 18392
rect 44880 18380 44914 18392
rect 44380 18302 44386 18314
rect 44386 18302 44414 18314
rect 44380 18280 44414 18302
rect 44480 18280 44514 18314
rect 44580 18280 44614 18314
rect 44680 18302 44712 18314
rect 44712 18302 44714 18314
rect 44780 18302 44802 18314
rect 44802 18302 44814 18314
rect 44880 18302 44892 18314
rect 44892 18302 44914 18314
rect 44680 18280 44714 18302
rect 44780 18280 44814 18302
rect 44880 18280 44914 18302
rect 44380 18212 44386 18214
rect 44386 18212 44414 18214
rect 44380 18180 44414 18212
rect 44480 18180 44514 18214
rect 44580 18180 44614 18214
rect 44680 18212 44712 18214
rect 44712 18212 44714 18214
rect 44780 18212 44802 18214
rect 44802 18212 44814 18214
rect 44880 18212 44892 18214
rect 44892 18212 44914 18214
rect 44680 18180 44714 18212
rect 44780 18180 44814 18212
rect 44880 18180 44914 18212
rect 44380 18080 44414 18114
rect 44480 18080 44514 18114
rect 44580 18080 44614 18114
rect 44680 18080 44714 18114
rect 44780 18080 44814 18114
rect 44880 18080 44914 18114
rect 44380 17980 44414 18014
rect 44480 17980 44514 18014
rect 44580 17980 44614 18014
rect 44680 17980 44714 18014
rect 44780 17980 44814 18014
rect 44880 17980 44914 18014
rect 44380 17886 44414 17914
rect 44380 17880 44386 17886
rect 44386 17880 44414 17886
rect 44480 17880 44514 17914
rect 44580 17880 44614 17914
rect 44680 17886 44714 17914
rect 44780 17886 44814 17914
rect 44880 17886 44914 17914
rect 44680 17880 44712 17886
rect 44712 17880 44714 17886
rect 44780 17880 44802 17886
rect 44802 17880 44814 17886
rect 44880 17880 44892 17886
rect 44892 17880 44914 17886
rect 45690 18597 45730 18610
rect 45690 18570 45730 18597
rect 46800 18595 46840 18610
rect 41660 17032 41666 17054
rect 41666 17032 41694 17054
rect 41660 17020 41694 17032
rect 41760 17020 41794 17054
rect 41860 17020 41894 17054
rect 41960 17032 41992 17054
rect 41992 17032 41994 17054
rect 42060 17032 42082 17054
rect 42082 17032 42094 17054
rect 42160 17032 42172 17054
rect 42172 17032 42194 17054
rect 41960 17020 41994 17032
rect 42060 17020 42094 17032
rect 42160 17020 42194 17032
rect 41660 16942 41666 16954
rect 41666 16942 41694 16954
rect 41660 16920 41694 16942
rect 41760 16920 41794 16954
rect 41860 16920 41894 16954
rect 41960 16942 41992 16954
rect 41992 16942 41994 16954
rect 42060 16942 42082 16954
rect 42082 16942 42094 16954
rect 42160 16942 42172 16954
rect 42172 16942 42194 16954
rect 41960 16920 41994 16942
rect 42060 16920 42094 16942
rect 42160 16920 42194 16942
rect 41660 16852 41666 16854
rect 41666 16852 41694 16854
rect 41660 16820 41694 16852
rect 41760 16820 41794 16854
rect 41860 16820 41894 16854
rect 41960 16852 41992 16854
rect 41992 16852 41994 16854
rect 42060 16852 42082 16854
rect 42082 16852 42094 16854
rect 42160 16852 42172 16854
rect 42172 16852 42194 16854
rect 41960 16820 41994 16852
rect 42060 16820 42094 16852
rect 42160 16820 42194 16852
rect 41660 16720 41694 16754
rect 41760 16720 41794 16754
rect 41860 16720 41894 16754
rect 41960 16720 41994 16754
rect 42060 16720 42094 16754
rect 42160 16720 42194 16754
rect 41660 16620 41694 16654
rect 41760 16620 41794 16654
rect 41860 16620 41894 16654
rect 41960 16620 41994 16654
rect 42060 16620 42094 16654
rect 42160 16620 42194 16654
rect 41660 16526 41694 16554
rect 41660 16520 41666 16526
rect 41666 16520 41694 16526
rect 41760 16520 41794 16554
rect 41860 16520 41894 16554
rect 41960 16526 41994 16554
rect 42060 16526 42094 16554
rect 42160 16526 42194 16554
rect 41960 16520 41992 16526
rect 41992 16520 41994 16526
rect 42060 16520 42082 16526
rect 42082 16520 42094 16526
rect 42160 16520 42172 16526
rect 42172 16520 42194 16526
rect 43020 17032 43026 17054
rect 43026 17032 43054 17054
rect 43020 17020 43054 17032
rect 43120 17020 43154 17054
rect 43220 17020 43254 17054
rect 43320 17032 43352 17054
rect 43352 17032 43354 17054
rect 43420 17032 43442 17054
rect 43442 17032 43454 17054
rect 43520 17032 43532 17054
rect 43532 17032 43554 17054
rect 43320 17020 43354 17032
rect 43420 17020 43454 17032
rect 43520 17020 43554 17032
rect 43020 16942 43026 16954
rect 43026 16942 43054 16954
rect 43020 16920 43054 16942
rect 43120 16920 43154 16954
rect 43220 16920 43254 16954
rect 43320 16942 43352 16954
rect 43352 16942 43354 16954
rect 43420 16942 43442 16954
rect 43442 16942 43454 16954
rect 43520 16942 43532 16954
rect 43532 16942 43554 16954
rect 43320 16920 43354 16942
rect 43420 16920 43454 16942
rect 43520 16920 43554 16942
rect 43020 16852 43026 16854
rect 43026 16852 43054 16854
rect 43020 16820 43054 16852
rect 43120 16820 43154 16854
rect 43220 16820 43254 16854
rect 43320 16852 43352 16854
rect 43352 16852 43354 16854
rect 43420 16852 43442 16854
rect 43442 16852 43454 16854
rect 43520 16852 43532 16854
rect 43532 16852 43554 16854
rect 43320 16820 43354 16852
rect 43420 16820 43454 16852
rect 43520 16820 43554 16852
rect 43020 16720 43054 16754
rect 43120 16720 43154 16754
rect 43220 16720 43254 16754
rect 43320 16720 43354 16754
rect 43420 16720 43454 16754
rect 43520 16720 43554 16754
rect 43020 16620 43054 16654
rect 43120 16620 43154 16654
rect 43220 16620 43254 16654
rect 43320 16620 43354 16654
rect 43420 16620 43454 16654
rect 43520 16620 43554 16654
rect 43020 16526 43054 16554
rect 43020 16520 43026 16526
rect 43026 16520 43054 16526
rect 43120 16520 43154 16554
rect 43220 16520 43254 16554
rect 43320 16526 43354 16554
rect 43420 16526 43454 16554
rect 43520 16526 43554 16554
rect 43320 16520 43352 16526
rect 43352 16520 43354 16526
rect 43420 16520 43442 16526
rect 43442 16520 43454 16526
rect 43520 16520 43532 16526
rect 43532 16520 43554 16526
rect 44380 17032 44386 17054
rect 44386 17032 44414 17054
rect 44380 17020 44414 17032
rect 44480 17020 44514 17054
rect 44580 17020 44614 17054
rect 44680 17032 44712 17054
rect 44712 17032 44714 17054
rect 44780 17032 44802 17054
rect 44802 17032 44814 17054
rect 44880 17032 44892 17054
rect 44892 17032 44914 17054
rect 44680 17020 44714 17032
rect 44780 17020 44814 17032
rect 44880 17020 44914 17032
rect 44380 16942 44386 16954
rect 44386 16942 44414 16954
rect 44380 16920 44414 16942
rect 44480 16920 44514 16954
rect 44580 16920 44614 16954
rect 44680 16942 44712 16954
rect 44712 16942 44714 16954
rect 44780 16942 44802 16954
rect 44802 16942 44814 16954
rect 44880 16942 44892 16954
rect 44892 16942 44914 16954
rect 44680 16920 44714 16942
rect 44780 16920 44814 16942
rect 44880 16920 44914 16942
rect 44380 16852 44386 16854
rect 44386 16852 44414 16854
rect 44380 16820 44414 16852
rect 44480 16820 44514 16854
rect 44580 16820 44614 16854
rect 44680 16852 44712 16854
rect 44712 16852 44714 16854
rect 44780 16852 44802 16854
rect 44802 16852 44814 16854
rect 44880 16852 44892 16854
rect 44892 16852 44914 16854
rect 44680 16820 44714 16852
rect 44780 16820 44814 16852
rect 44880 16820 44914 16852
rect 44380 16720 44414 16754
rect 44480 16720 44514 16754
rect 44580 16720 44614 16754
rect 44680 16720 44714 16754
rect 44780 16720 44814 16754
rect 44880 16720 44914 16754
rect 44380 16620 44414 16654
rect 44480 16620 44514 16654
rect 44580 16620 44614 16654
rect 44680 16620 44714 16654
rect 44780 16620 44814 16654
rect 44880 16620 44914 16654
rect 44380 16526 44414 16554
rect 44380 16520 44386 16526
rect 44386 16520 44414 16526
rect 44480 16520 44514 16554
rect 44580 16520 44614 16554
rect 44680 16526 44714 16554
rect 44780 16526 44814 16554
rect 44880 16526 44914 16554
rect 44680 16520 44712 16526
rect 44712 16520 44714 16526
rect 44780 16520 44802 16526
rect 44802 16520 44814 16526
rect 44880 16520 44892 16526
rect 44892 16520 44914 16526
rect 45690 18050 45730 18440
rect 46020 16310 46060 16700
rect 46800 18570 46840 18595
rect 47590 18589 47630 18590
rect 41660 15672 41666 15694
rect 41666 15672 41694 15694
rect 41660 15660 41694 15672
rect 41760 15660 41794 15694
rect 41860 15660 41894 15694
rect 41960 15672 41992 15694
rect 41992 15672 41994 15694
rect 42060 15672 42082 15694
rect 42082 15672 42094 15694
rect 42160 15672 42172 15694
rect 42172 15672 42194 15694
rect 41960 15660 41994 15672
rect 42060 15660 42094 15672
rect 42160 15660 42194 15672
rect 41660 15582 41666 15594
rect 41666 15582 41694 15594
rect 41660 15560 41694 15582
rect 41760 15560 41794 15594
rect 41860 15560 41894 15594
rect 41960 15582 41992 15594
rect 41992 15582 41994 15594
rect 42060 15582 42082 15594
rect 42082 15582 42094 15594
rect 42160 15582 42172 15594
rect 42172 15582 42194 15594
rect 41960 15560 41994 15582
rect 42060 15560 42094 15582
rect 42160 15560 42194 15582
rect 41660 15492 41666 15494
rect 41666 15492 41694 15494
rect 41660 15460 41694 15492
rect 41760 15460 41794 15494
rect 41860 15460 41894 15494
rect 41960 15492 41992 15494
rect 41992 15492 41994 15494
rect 42060 15492 42082 15494
rect 42082 15492 42094 15494
rect 42160 15492 42172 15494
rect 42172 15492 42194 15494
rect 41960 15460 41994 15492
rect 42060 15460 42094 15492
rect 42160 15460 42194 15492
rect 41660 15360 41694 15394
rect 41760 15360 41794 15394
rect 41860 15360 41894 15394
rect 41960 15360 41994 15394
rect 42060 15360 42094 15394
rect 42160 15360 42194 15394
rect 41660 15260 41694 15294
rect 41760 15260 41794 15294
rect 41860 15260 41894 15294
rect 41960 15260 41994 15294
rect 42060 15260 42094 15294
rect 42160 15260 42194 15294
rect 41660 15166 41694 15194
rect 41660 15160 41666 15166
rect 41666 15160 41694 15166
rect 41760 15160 41794 15194
rect 41860 15160 41894 15194
rect 41960 15166 41994 15194
rect 42060 15166 42094 15194
rect 42160 15166 42194 15194
rect 41960 15160 41992 15166
rect 41992 15160 41994 15166
rect 42060 15160 42082 15166
rect 42082 15160 42094 15166
rect 42160 15160 42172 15166
rect 42172 15160 42194 15166
rect 43020 15672 43026 15694
rect 43026 15672 43054 15694
rect 43020 15660 43054 15672
rect 43120 15660 43154 15694
rect 43220 15660 43254 15694
rect 43320 15672 43352 15694
rect 43352 15672 43354 15694
rect 43420 15672 43442 15694
rect 43442 15672 43454 15694
rect 43520 15672 43532 15694
rect 43532 15672 43554 15694
rect 43320 15660 43354 15672
rect 43420 15660 43454 15672
rect 43520 15660 43554 15672
rect 43020 15582 43026 15594
rect 43026 15582 43054 15594
rect 43020 15560 43054 15582
rect 43120 15560 43154 15594
rect 43220 15560 43254 15594
rect 43320 15582 43352 15594
rect 43352 15582 43354 15594
rect 43420 15582 43442 15594
rect 43442 15582 43454 15594
rect 43520 15582 43532 15594
rect 43532 15582 43554 15594
rect 43320 15560 43354 15582
rect 43420 15560 43454 15582
rect 43520 15560 43554 15582
rect 43020 15492 43026 15494
rect 43026 15492 43054 15494
rect 43020 15460 43054 15492
rect 43120 15460 43154 15494
rect 43220 15460 43254 15494
rect 43320 15492 43352 15494
rect 43352 15492 43354 15494
rect 43420 15492 43442 15494
rect 43442 15492 43454 15494
rect 43520 15492 43532 15494
rect 43532 15492 43554 15494
rect 43320 15460 43354 15492
rect 43420 15460 43454 15492
rect 43520 15460 43554 15492
rect 43020 15360 43054 15394
rect 43120 15360 43154 15394
rect 43220 15360 43254 15394
rect 43320 15360 43354 15394
rect 43420 15360 43454 15394
rect 43520 15360 43554 15394
rect 43020 15260 43054 15294
rect 43120 15260 43154 15294
rect 43220 15260 43254 15294
rect 43320 15260 43354 15294
rect 43420 15260 43454 15294
rect 43520 15260 43554 15294
rect 43020 15166 43054 15194
rect 43020 15160 43026 15166
rect 43026 15160 43054 15166
rect 43120 15160 43154 15194
rect 43220 15160 43254 15194
rect 43320 15166 43354 15194
rect 43420 15166 43454 15194
rect 43520 15166 43554 15194
rect 43320 15160 43352 15166
rect 43352 15160 43354 15166
rect 43420 15160 43442 15166
rect 43442 15160 43454 15166
rect 43520 15160 43532 15166
rect 43532 15160 43554 15166
rect 44380 15672 44386 15694
rect 44386 15672 44414 15694
rect 44380 15660 44414 15672
rect 44480 15660 44514 15694
rect 44580 15660 44614 15694
rect 44680 15672 44712 15694
rect 44712 15672 44714 15694
rect 44780 15672 44802 15694
rect 44802 15672 44814 15694
rect 44880 15672 44892 15694
rect 44892 15672 44914 15694
rect 44680 15660 44714 15672
rect 44780 15660 44814 15672
rect 44880 15660 44914 15672
rect 44380 15582 44386 15594
rect 44386 15582 44414 15594
rect 44380 15560 44414 15582
rect 44480 15560 44514 15594
rect 44580 15560 44614 15594
rect 44680 15582 44712 15594
rect 44712 15582 44714 15594
rect 44780 15582 44802 15594
rect 44802 15582 44814 15594
rect 44880 15582 44892 15594
rect 44892 15582 44914 15594
rect 44680 15560 44714 15582
rect 44780 15560 44814 15582
rect 44880 15560 44914 15582
rect 44380 15492 44386 15494
rect 44386 15492 44414 15494
rect 44380 15460 44414 15492
rect 44480 15460 44514 15494
rect 44580 15460 44614 15494
rect 44680 15492 44712 15494
rect 44712 15492 44714 15494
rect 44780 15492 44802 15494
rect 44802 15492 44814 15494
rect 44880 15492 44892 15494
rect 44892 15492 44914 15494
rect 44680 15460 44714 15492
rect 44780 15460 44814 15492
rect 44880 15460 44914 15492
rect 44380 15360 44414 15394
rect 44480 15360 44514 15394
rect 44580 15360 44614 15394
rect 44680 15360 44714 15394
rect 44780 15360 44814 15394
rect 44880 15360 44914 15394
rect 44380 15260 44414 15294
rect 44480 15260 44514 15294
rect 44580 15260 44614 15294
rect 44680 15260 44714 15294
rect 44780 15260 44814 15294
rect 44880 15260 44914 15294
rect 44380 15166 44414 15194
rect 44380 15160 44386 15166
rect 44386 15160 44414 15166
rect 44480 15160 44514 15194
rect 44580 15160 44614 15194
rect 44680 15166 44714 15194
rect 44780 15166 44814 15194
rect 44880 15166 44914 15194
rect 44680 15160 44712 15166
rect 44712 15160 44714 15166
rect 44780 15160 44802 15166
rect 44802 15160 44814 15166
rect 44880 15160 44892 15166
rect 44892 15160 44914 15166
rect 46800 18041 46838 18438
rect 46800 15970 46838 16367
rect 47590 18555 47630 18589
rect 47590 18550 47630 18555
rect 47556 18035 47662 18432
rect 47556 16650 47662 17047
rect 41560 14350 41960 14402
rect 44599 14360 44996 14398
rect 41100 13760 41140 13800
rect 45490 13800 45530 13840
rect 45490 13720 45530 13760
rect 41180 13590 41220 13630
rect 41340 13590 41380 13630
rect 41500 13590 41540 13630
rect 41660 13590 41700 13630
rect 41820 13590 41860 13630
rect 41980 13590 42020 13630
rect 42140 13590 42180 13630
rect 42300 13590 42340 13630
rect 42460 13590 42500 13630
rect 42620 13590 42660 13630
rect 42780 13590 42820 13630
rect 42940 13590 42980 13630
rect 43100 13590 43140 13630
rect 43260 13590 43300 13630
rect 43420 13590 43460 13630
rect 43580 13590 43620 13630
rect 43740 13590 43780 13630
rect 43900 13590 43940 13630
rect 44060 13590 44100 13630
rect 44220 13590 44260 13630
rect 44380 13590 44420 13630
rect 44540 13590 44580 13630
rect 44700 13590 44740 13630
rect 44860 13590 44900 13630
rect 45020 13590 45060 13630
rect 45180 13590 45220 13630
rect 41920 13320 41960 13360
rect 44600 13320 44640 13360
rect 40760 12720 40800 12760
rect 40940 12680 40980 12720
rect 41180 12680 41220 12720
rect 41420 12680 41460 12720
rect 41660 12680 41700 12720
rect 42300 12680 42340 12720
rect 42540 12680 42580 12720
rect 42780 12680 42820 12720
rect 43080 12710 43120 12750
rect 45760 13200 45800 13240
rect 45760 13100 45800 13140
rect 45760 13000 45800 13040
rect 45760 12900 45800 12940
rect 45760 12800 45800 12840
rect 43440 12710 43480 12750
rect 43740 12680 43780 12720
rect 43980 12680 44020 12720
rect 44220 12680 44260 12720
rect 44860 12680 44900 12720
rect 45100 12680 45140 12720
rect 45340 12680 45380 12720
rect 45580 12680 45620 12720
rect 41443 12308 41477 12342
rect 41803 12308 41837 12342
rect 41923 12308 41957 12342
rect 42283 12308 42317 12342
rect 42403 12308 42437 12342
rect 42820 12280 42860 12320
rect 41380 12190 41420 12230
rect 41500 12190 41540 12230
rect 41620 12190 41660 12230
rect 41740 12190 41780 12230
rect 41860 12190 41900 12230
rect 41980 12190 42020 12230
rect 42100 12190 42140 12230
rect 42220 12190 42260 12230
rect 42340 12190 42380 12230
rect 42460 12190 42500 12230
rect 42580 12190 42620 12230
rect 42820 12200 42860 12240
rect 41544 12078 41578 12112
rect 41702 12078 41736 12112
rect 42026 12078 42060 12112
rect 42180 12078 42214 12112
rect 42504 12078 42538 12112
rect 42820 12120 42860 12160
rect 43700 12280 43740 12320
rect 44123 12308 44157 12342
rect 44243 12308 44277 12342
rect 44603 12308 44637 12342
rect 44723 12308 44757 12342
rect 45083 12308 45117 12342
rect 43700 12200 43740 12240
rect 43940 12190 43980 12230
rect 44060 12190 44100 12230
rect 44180 12190 44220 12230
rect 44300 12190 44340 12230
rect 44420 12190 44460 12230
rect 44540 12190 44580 12230
rect 44660 12190 44700 12230
rect 44780 12190 44820 12230
rect 44900 12190 44940 12230
rect 45020 12190 45060 12230
rect 45140 12190 45180 12230
rect 43700 12120 43740 12160
rect 44022 12078 44056 12112
rect 44346 12078 44380 12112
rect 44500 12078 44534 12112
rect 44824 12078 44858 12112
rect 44982 12078 45016 12112
rect 40720 11480 40760 11520
rect 40900 11470 40940 11510
rect 41380 11470 41420 11510
rect 41620 11470 41660 11510
rect 42100 11470 42140 11510
rect 42340 11470 42380 11510
rect 42760 11470 42800 11510
rect 43760 11470 43800 11510
rect 44180 11470 44220 11510
rect 44420 11470 44460 11510
rect 44900 11470 44940 11510
rect 45140 11470 45180 11510
rect 45620 11470 45660 11510
rect 45800 11480 45840 11520
rect 40540 11350 40580 11390
rect 40540 11250 40580 11290
rect 40660 11350 40700 11390
rect 40660 11250 40700 11290
rect 40780 11350 40820 11390
rect 40780 11250 40820 11290
rect 40900 11350 40940 11390
rect 40900 11250 40940 11290
rect 41020 11350 41060 11390
rect 41020 11250 41060 11290
rect 41140 11350 41180 11390
rect 41140 11250 41180 11290
rect 41260 11350 41300 11390
rect 41260 11250 41300 11290
rect 41380 11350 41420 11390
rect 41380 11250 41420 11290
rect 41500 11350 41540 11390
rect 41500 11250 41540 11290
rect 41620 11350 41660 11390
rect 41620 11250 41660 11290
rect 41740 11350 41780 11390
rect 41740 11250 41780 11290
rect 41860 11350 41900 11390
rect 41860 11250 41900 11290
rect 41980 11350 42020 11390
rect 41980 11250 42020 11290
rect 42100 11350 42140 11390
rect 42100 11250 42140 11290
rect 42220 11350 42260 11390
rect 42220 11250 42260 11290
rect 42340 11350 42380 11390
rect 42340 11250 42380 11290
rect 42460 11350 42500 11390
rect 42460 11250 42500 11290
rect 42580 11350 42620 11390
rect 42580 11250 42620 11290
rect 42700 11350 42740 11390
rect 42700 11250 42740 11290
rect 42820 11350 42860 11390
rect 42820 11250 42860 11290
rect 42940 11350 42980 11390
rect 42940 11250 42980 11290
rect 43580 11350 43620 11390
rect 43580 11250 43620 11290
rect 43700 11350 43740 11390
rect 43700 11250 43740 11290
rect 43820 11350 43860 11390
rect 43820 11250 43860 11290
rect 43940 11350 43980 11390
rect 43940 11250 43980 11290
rect 44060 11350 44100 11390
rect 44060 11250 44100 11290
rect 44180 11350 44220 11390
rect 44180 11250 44220 11290
rect 44300 11350 44340 11390
rect 44300 11250 44340 11290
rect 44420 11350 44460 11390
rect 44420 11250 44460 11290
rect 44540 11350 44580 11390
rect 44540 11250 44580 11290
rect 44660 11350 44700 11390
rect 44660 11250 44700 11290
rect 44780 11350 44820 11390
rect 44780 11250 44820 11290
rect 44900 11350 44940 11390
rect 44900 11250 44940 11290
rect 45020 11350 45060 11390
rect 45020 11250 45060 11290
rect 45140 11350 45180 11390
rect 45140 11250 45180 11290
rect 45260 11350 45300 11390
rect 45260 11250 45300 11290
rect 45380 11350 45420 11390
rect 45380 11250 45420 11290
rect 45500 11350 45540 11390
rect 45500 11250 45540 11290
rect 45620 11350 45660 11390
rect 45620 11250 45660 11290
rect 45740 11350 45780 11390
rect 45740 11250 45780 11290
rect 45860 11350 45900 11390
rect 45860 11250 45900 11290
rect 45980 11350 46020 11390
rect 45980 11250 46020 11290
rect 40540 11130 40580 11170
rect 42940 11130 42980 11170
rect 43580 11130 43620 11170
rect 45980 11130 46020 11170
rect 41910 10310 41950 10350
rect 42090 10310 42130 10350
rect 42270 10310 42310 10350
rect 42450 10310 42490 10350
rect 42630 10310 42670 10350
rect 42810 10310 42850 10350
rect 42990 10310 43030 10350
rect 43170 10310 43210 10350
rect 43350 10310 43390 10350
rect 43530 10310 43570 10350
rect 43710 10310 43750 10350
rect 43890 10310 43930 10350
rect 44070 10310 44110 10350
rect 44250 10310 44290 10350
rect 44430 10310 44470 10350
rect 44610 10310 44650 10350
rect 41640 10190 41680 10230
rect 41640 10090 41680 10130
rect 41640 9990 41680 10030
rect 41640 9890 41680 9930
rect 41640 9790 41680 9830
rect 41640 9690 41680 9730
rect 41820 10190 41860 10230
rect 41820 10090 41860 10130
rect 41820 9990 41860 10030
rect 41820 9890 41860 9930
rect 41820 9790 41860 9830
rect 41820 9690 41860 9730
rect 42000 10190 42040 10230
rect 42000 10090 42040 10130
rect 42000 9990 42040 10030
rect 42000 9890 42040 9930
rect 42000 9790 42040 9830
rect 42000 9690 42040 9730
rect 42180 10190 42220 10230
rect 42180 10090 42220 10130
rect 42180 9990 42220 10030
rect 42180 9890 42220 9930
rect 42180 9790 42220 9830
rect 42180 9690 42220 9730
rect 42360 10190 42400 10230
rect 42360 10090 42400 10130
rect 42360 9990 42400 10030
rect 42360 9890 42400 9930
rect 42360 9790 42400 9830
rect 42360 9690 42400 9730
rect 42540 10190 42580 10230
rect 42540 10090 42580 10130
rect 42540 9990 42580 10030
rect 42540 9890 42580 9930
rect 42540 9790 42580 9830
rect 42540 9690 42580 9730
rect 42720 10190 42760 10230
rect 42720 10090 42760 10130
rect 42720 9990 42760 10030
rect 42720 9890 42760 9930
rect 42720 9790 42760 9830
rect 42720 9690 42760 9730
rect 42900 10190 42940 10230
rect 42900 10090 42940 10130
rect 42900 9990 42940 10030
rect 42900 9890 42940 9930
rect 42900 9790 42940 9830
rect 42900 9690 42940 9730
rect 43080 10190 43120 10230
rect 43080 10090 43120 10130
rect 43080 9990 43120 10030
rect 43080 9890 43120 9930
rect 43080 9790 43120 9830
rect 43080 9690 43120 9730
rect 43260 10190 43300 10230
rect 43260 10090 43300 10130
rect 43260 9990 43300 10030
rect 43260 9890 43300 9930
rect 43260 9790 43300 9830
rect 43260 9690 43300 9730
rect 43440 10190 43480 10230
rect 43440 10090 43480 10130
rect 43440 9990 43480 10030
rect 43440 9890 43480 9930
rect 43440 9790 43480 9830
rect 43440 9690 43480 9730
rect 43620 10190 43660 10230
rect 43620 10090 43660 10130
rect 43620 9990 43660 10030
rect 43620 9890 43660 9930
rect 43620 9790 43660 9830
rect 43620 9690 43660 9730
rect 43800 10190 43840 10230
rect 43800 10090 43840 10130
rect 43800 9990 43840 10030
rect 43800 9890 43840 9930
rect 43800 9790 43840 9830
rect 43800 9690 43840 9730
rect 43980 10190 44020 10230
rect 43980 10090 44020 10130
rect 43980 9990 44020 10030
rect 43980 9890 44020 9930
rect 43980 9790 44020 9830
rect 43980 9690 44020 9730
rect 44160 10190 44200 10230
rect 44160 10090 44200 10130
rect 44160 9990 44200 10030
rect 44160 9890 44200 9930
rect 44160 9790 44200 9830
rect 44160 9690 44200 9730
rect 44340 10190 44380 10230
rect 44340 10090 44380 10130
rect 44340 9990 44380 10030
rect 44340 9890 44380 9930
rect 44340 9790 44380 9830
rect 44340 9690 44380 9730
rect 44520 10190 44560 10230
rect 44520 10090 44560 10130
rect 44520 9990 44560 10030
rect 44520 9890 44560 9930
rect 44520 9790 44560 9830
rect 44520 9690 44560 9730
rect 44700 10190 44740 10230
rect 44700 10090 44740 10130
rect 44700 9990 44740 10030
rect 44700 9890 44740 9930
rect 44700 9790 44740 9830
rect 44700 9690 44740 9730
rect 44880 10190 44920 10230
rect 44880 10090 44920 10130
rect 45610 10110 45650 10150
rect 45730 10110 45770 10150
rect 45850 10110 45890 10150
rect 44880 9990 44920 10030
rect 44880 9890 44920 9930
rect 45510 9990 45550 10030
rect 45510 9890 45550 9930
rect 45620 9990 45660 10030
rect 45620 9890 45660 9930
rect 45730 9990 45770 10030
rect 45730 9890 45770 9930
rect 45840 9990 45880 10030
rect 45840 9890 45880 9930
rect 45950 9990 45990 10030
rect 45950 9890 45990 9930
rect 44880 9790 44920 9830
rect 45510 9770 45550 9810
rect 45730 9770 45770 9810
rect 45950 9770 45990 9810
rect 44880 9690 44920 9730
rect 41640 9570 41680 9610
rect 42000 9570 42040 9610
rect 42360 9570 42400 9610
rect 42720 9570 42760 9610
rect 43080 9570 43120 9610
rect 43440 9570 43480 9610
rect 43800 9570 43840 9610
rect 44160 9570 44200 9610
rect 44520 9570 44560 9610
rect 44880 9570 44920 9610
rect 41818 9308 41852 9342
rect 41928 9308 41962 9342
rect 42038 9308 42072 9342
rect 42148 9308 42182 9342
rect 42258 9308 42292 9342
rect 42368 9308 42402 9342
rect 42478 9308 42512 9342
rect 42588 9308 42622 9342
rect 42698 9308 42732 9342
rect 42808 9308 42842 9342
rect 43718 9308 43752 9342
rect 43828 9308 43862 9342
rect 43938 9308 43972 9342
rect 44048 9308 44082 9342
rect 44158 9308 44192 9342
rect 44268 9308 44302 9342
rect 44378 9308 44412 9342
rect 44488 9308 44522 9342
rect 44598 9308 44632 9342
rect 44708 9308 44742 9342
rect 41570 9190 41610 9230
rect 41650 9190 41690 9230
rect 41570 9090 41610 9130
rect 41650 9090 41690 9130
rect 41760 9190 41800 9230
rect 41760 9090 41800 9130
rect 41870 9190 41910 9230
rect 41870 9090 41910 9130
rect 41980 9190 42020 9230
rect 41980 9090 42020 9130
rect 42090 9190 42130 9230
rect 42090 9090 42130 9130
rect 42200 9190 42240 9230
rect 42200 9090 42240 9130
rect 42310 9190 42350 9230
rect 42310 9090 42350 9130
rect 42420 9190 42460 9230
rect 42420 9090 42460 9130
rect 42530 9190 42570 9230
rect 42530 9090 42570 9130
rect 42640 9190 42680 9230
rect 42640 9090 42680 9130
rect 42750 9190 42790 9230
rect 42750 9090 42790 9130
rect 42860 9190 42900 9230
rect 42860 9090 42900 9130
rect 42970 9190 43010 9230
rect 43050 9190 43090 9230
rect 42970 9090 43010 9130
rect 43050 9090 43090 9130
rect 43470 9190 43510 9230
rect 43550 9190 43590 9230
rect 43470 9090 43510 9130
rect 43550 9090 43590 9130
rect 43660 9190 43700 9230
rect 43660 9090 43700 9130
rect 43770 9190 43810 9230
rect 43770 9090 43810 9130
rect 43880 9190 43920 9230
rect 43880 9090 43920 9130
rect 43990 9190 44030 9230
rect 43990 9090 44030 9130
rect 44100 9190 44140 9230
rect 44100 9090 44140 9130
rect 44210 9190 44250 9230
rect 44210 9090 44250 9130
rect 44320 9190 44360 9230
rect 44320 9090 44360 9130
rect 44430 9190 44470 9230
rect 44430 9090 44470 9130
rect 44540 9190 44580 9230
rect 44540 9090 44580 9130
rect 44650 9190 44690 9230
rect 44650 9090 44690 9130
rect 44760 9190 44800 9230
rect 44760 9090 44800 9130
rect 44870 9190 44910 9230
rect 44950 9190 44990 9230
rect 44870 9090 44910 9130
rect 44950 9090 44990 9130
rect 41650 8970 41690 9010
rect 42970 8970 43010 9010
rect 43550 8970 43590 9010
rect 44870 8970 44910 9010
<< metal1 >>
rect 39170 19190 39250 19200
rect 39170 19130 39180 19190
rect 39240 19130 39250 19190
rect 38790 19080 38870 19090
rect 38790 19020 38800 19080
rect 38860 19020 38870 19080
rect 38790 19000 38870 19020
rect 38790 18940 38800 19000
rect 38860 18940 38870 19000
rect 38790 18920 38870 18940
rect 38790 18860 38800 18920
rect 38860 18860 38870 18920
rect 38790 18590 38870 18860
rect 38790 18550 38810 18590
rect 38850 18550 38870 18590
rect 38790 18530 38870 18550
rect 39170 18450 39250 19130
rect 38770 18432 38888 18444
rect 38770 18035 38776 18432
rect 38882 18035 38888 18432
rect 38770 18023 38888 18035
rect 39170 18390 39180 18450
rect 39240 18390 39250 18450
rect 39170 18370 39250 18390
rect 39170 18310 39180 18370
rect 39240 18310 39250 18370
rect 39170 18280 39250 18310
rect 39170 18220 39180 18280
rect 39240 18220 39250 18280
rect 39170 18190 39250 18220
rect 39170 18130 39180 18190
rect 39240 18130 39250 18190
rect 39170 18110 39250 18130
rect 39170 18050 39180 18110
rect 39240 18050 39250 18110
rect 39170 18030 39250 18050
rect 39570 19080 39650 19090
rect 39570 19020 39580 19080
rect 39640 19020 39650 19080
rect 39570 19000 39650 19020
rect 39570 18940 39580 19000
rect 39640 18940 39650 19000
rect 39570 18920 39650 18940
rect 39570 18860 39580 18920
rect 39640 18860 39650 18920
rect 39570 18600 39650 18860
rect 39570 18560 39590 18600
rect 39630 18560 39650 18600
rect 39570 18438 39650 18560
rect 39570 18041 39590 18438
rect 39628 18041 39650 18438
rect 39570 18020 39650 18041
rect 40680 19080 40760 19090
rect 40680 19020 40690 19080
rect 40750 19020 40760 19080
rect 40680 19000 40760 19020
rect 40680 18940 40690 19000
rect 40750 18940 40760 19000
rect 40680 18920 40760 18940
rect 40680 18860 40690 18920
rect 40750 18860 40760 18920
rect 40680 18610 40760 18860
rect 40680 18570 40700 18610
rect 40740 18570 40760 18610
rect 40680 18440 40760 18570
rect 40680 18050 40700 18440
rect 40740 18050 40760 18440
rect 40680 18030 40760 18050
rect 38770 17047 38888 17059
rect 38770 16650 38776 17047
rect 38882 16650 38888 17047
rect 38770 16638 38888 16650
rect 40350 16700 40430 16720
rect 38790 11180 38870 16638
rect 40350 16310 40370 16700
rect 40410 16310 40430 16700
rect 39570 15477 39650 15500
rect 39570 15080 39590 15477
rect 39628 15080 39650 15477
rect 38790 11120 38800 11180
rect 38860 11120 38870 11180
rect 38790 9360 38870 11120
rect 39460 13810 39540 13820
rect 39460 13750 39470 13810
rect 39530 13750 39540 13810
rect 39460 10690 39540 13750
rect 39570 12120 39650 15080
rect 40350 14720 40430 16310
rect 40350 14660 40360 14720
rect 40420 14660 40430 14720
rect 40350 14650 40430 14660
rect 39570 12060 39580 12120
rect 39640 12060 39650 12120
rect 39570 10800 39650 12060
rect 39570 10740 39580 10800
rect 39640 10740 39650 10800
rect 39570 10730 39650 10740
rect 39680 14090 39760 14100
rect 39680 14030 39690 14090
rect 39750 14030 39760 14090
rect 39680 12350 39760 14030
rect 39680 12290 39690 12350
rect 39750 12290 39760 12350
rect 39460 10630 39470 10690
rect 39530 10630 39540 10690
rect 39460 10620 39540 10630
rect 38790 9300 38800 9360
rect 38860 9300 38870 9360
rect 38790 9290 38870 9300
rect 39680 8910 39760 12290
rect 40620 13980 40700 13990
rect 40620 13920 40630 13980
rect 40690 13920 40700 13980
rect 40620 11650 40700 13920
rect 41030 13980 41110 19200
rect 48190 19190 48270 19200
rect 48190 19130 48200 19190
rect 48260 19130 48270 19190
rect 43240 19080 43320 19090
rect 43240 19020 43250 19080
rect 43310 19020 43320 19080
rect 43240 19000 43320 19020
rect 43240 18940 43250 19000
rect 43310 18940 43320 19000
rect 43240 18920 43320 18940
rect 43240 18860 43250 18920
rect 43310 18860 43320 18920
rect 43240 18850 43320 18860
rect 45670 19080 45750 19090
rect 45670 19020 45680 19080
rect 45740 19020 45750 19080
rect 45670 19000 45750 19020
rect 45670 18940 45680 19000
rect 45740 18940 45750 19000
rect 45670 18920 45750 18940
rect 45670 18860 45680 18920
rect 45740 18860 45750 18920
rect 45670 18610 45750 18860
rect 45670 18570 45690 18610
rect 45730 18570 45750 18610
rect 41570 18414 44990 18490
rect 41570 18380 41660 18414
rect 41694 18380 41760 18414
rect 41794 18380 41860 18414
rect 41894 18380 41960 18414
rect 41994 18380 42060 18414
rect 42094 18380 42160 18414
rect 42194 18380 43020 18414
rect 43054 18380 43120 18414
rect 43154 18380 43220 18414
rect 43254 18380 43320 18414
rect 43354 18380 43420 18414
rect 43454 18380 43520 18414
rect 43554 18380 44380 18414
rect 44414 18380 44480 18414
rect 44514 18380 44580 18414
rect 44614 18380 44680 18414
rect 44714 18380 44780 18414
rect 44814 18380 44880 18414
rect 44914 18380 44990 18414
rect 41570 18314 44990 18380
rect 41570 18280 41660 18314
rect 41694 18280 41760 18314
rect 41794 18280 41860 18314
rect 41894 18280 41960 18314
rect 41994 18280 42060 18314
rect 42094 18280 42160 18314
rect 42194 18280 43020 18314
rect 43054 18280 43120 18314
rect 43154 18280 43220 18314
rect 43254 18280 43320 18314
rect 43354 18280 43420 18314
rect 43454 18280 43520 18314
rect 43554 18280 44380 18314
rect 44414 18280 44480 18314
rect 44514 18280 44580 18314
rect 44614 18280 44680 18314
rect 44714 18280 44780 18314
rect 44814 18280 44880 18314
rect 44914 18280 44990 18314
rect 41570 18214 44990 18280
rect 41570 18180 41660 18214
rect 41694 18180 41760 18214
rect 41794 18180 41860 18214
rect 41894 18180 41960 18214
rect 41994 18180 42060 18214
rect 42094 18180 42160 18214
rect 42194 18180 43020 18214
rect 43054 18180 43120 18214
rect 43154 18180 43220 18214
rect 43254 18180 43320 18214
rect 43354 18180 43420 18214
rect 43454 18180 43520 18214
rect 43554 18180 44380 18214
rect 44414 18180 44480 18214
rect 44514 18180 44580 18214
rect 44614 18180 44680 18214
rect 44714 18180 44780 18214
rect 44814 18180 44880 18214
rect 44914 18180 44990 18214
rect 41570 18114 44990 18180
rect 41570 18080 41660 18114
rect 41694 18080 41760 18114
rect 41794 18080 41860 18114
rect 41894 18080 41960 18114
rect 41994 18080 42060 18114
rect 42094 18080 42160 18114
rect 42194 18080 43020 18114
rect 43054 18080 43120 18114
rect 43154 18080 43220 18114
rect 43254 18080 43320 18114
rect 43354 18080 43420 18114
rect 43454 18080 43520 18114
rect 43554 18080 44380 18114
rect 44414 18080 44480 18114
rect 44514 18080 44580 18114
rect 44614 18080 44680 18114
rect 44714 18080 44780 18114
rect 44814 18080 44880 18114
rect 44914 18080 44990 18114
rect 41570 18014 44990 18080
rect 45670 18440 45750 18570
rect 45670 18050 45690 18440
rect 45730 18050 45750 18440
rect 45670 18030 45750 18050
rect 46780 19080 46860 19090
rect 46780 19020 46790 19080
rect 46850 19020 46860 19080
rect 46780 19000 46860 19020
rect 46780 18940 46790 19000
rect 46850 18940 46860 19000
rect 46780 18920 46860 18940
rect 46780 18860 46790 18920
rect 46850 18860 46860 18920
rect 46780 18610 46860 18860
rect 46780 18570 46800 18610
rect 46840 18570 46860 18610
rect 46780 18438 46860 18570
rect 47570 19080 47650 19090
rect 47570 19020 47580 19080
rect 47640 19020 47650 19080
rect 47570 19000 47650 19020
rect 47570 18940 47580 19000
rect 47640 18940 47650 19000
rect 47570 18920 47650 18940
rect 47570 18860 47580 18920
rect 47640 18860 47650 18920
rect 47570 18590 47650 18860
rect 48190 18850 48270 19130
rect 48190 18790 48200 18850
rect 48260 18790 48270 18850
rect 48190 18780 48270 18790
rect 47570 18550 47590 18590
rect 47630 18550 47650 18590
rect 47570 18530 47650 18550
rect 47950 18450 48030 18460
rect 46780 18041 46800 18438
rect 46838 18041 46860 18438
rect 46780 18030 46860 18041
rect 47550 18432 47668 18444
rect 47550 18035 47556 18432
rect 47662 18035 47668 18432
rect 46794 18029 46844 18030
rect 47550 18023 47668 18035
rect 47950 18390 47960 18450
rect 48020 18390 48030 18450
rect 47950 18370 48030 18390
rect 47950 18310 47960 18370
rect 48020 18310 48030 18370
rect 47950 18280 48030 18310
rect 47950 18220 47960 18280
rect 48020 18220 48030 18280
rect 47950 18190 48030 18220
rect 47950 18130 47960 18190
rect 48020 18130 48030 18190
rect 47950 18110 48030 18130
rect 47950 18050 47960 18110
rect 48020 18050 48030 18110
rect 48640 18150 48740 18170
rect 48640 18090 48660 18150
rect 48720 18090 48740 18150
rect 48640 18070 48740 18090
rect 41570 17980 41660 18014
rect 41694 17980 41760 18014
rect 41794 17980 41860 18014
rect 41894 17980 41960 18014
rect 41994 17980 42060 18014
rect 42094 17980 42160 18014
rect 42194 17980 43020 18014
rect 43054 17980 43120 18014
rect 43154 17980 43220 18014
rect 43254 17980 43320 18014
rect 43354 17980 43420 18014
rect 43454 17980 43520 18014
rect 43554 17980 44380 18014
rect 44414 17980 44480 18014
rect 44514 17980 44580 18014
rect 44614 17980 44680 18014
rect 44714 17980 44780 18014
rect 44814 17980 44880 18014
rect 44914 17980 44990 18014
rect 41570 17914 44990 17980
rect 41570 17880 41660 17914
rect 41694 17880 41760 17914
rect 41794 17880 41860 17914
rect 41894 17880 41960 17914
rect 41994 17880 42060 17914
rect 42094 17880 42160 17914
rect 42194 17880 43020 17914
rect 43054 17880 43120 17914
rect 43154 17880 43220 17914
rect 43254 17880 43320 17914
rect 43354 17880 43420 17914
rect 43454 17880 43520 17914
rect 43554 17880 44380 17914
rect 44414 17880 44480 17914
rect 44514 17880 44580 17914
rect 44614 17880 44680 17914
rect 44714 17880 44780 17914
rect 44814 17880 44880 17914
rect 44914 17880 44990 17914
rect 41570 17790 44990 17880
rect 41570 17054 42270 17790
rect 41570 17020 41660 17054
rect 41694 17020 41760 17054
rect 41794 17020 41860 17054
rect 41894 17020 41960 17054
rect 41994 17020 42060 17054
rect 42094 17020 42160 17054
rect 42194 17020 42270 17054
rect 41570 16954 42270 17020
rect 41570 16920 41660 16954
rect 41694 16920 41760 16954
rect 41794 16920 41860 16954
rect 41894 16920 41960 16954
rect 41994 16920 42060 16954
rect 42094 16920 42160 16954
rect 42194 16920 42270 16954
rect 41570 16854 42270 16920
rect 41570 16820 41660 16854
rect 41694 16820 41760 16854
rect 41794 16820 41860 16854
rect 41894 16820 41960 16854
rect 41994 16820 42060 16854
rect 42094 16820 42160 16854
rect 42194 16820 42270 16854
rect 41140 16810 41220 16820
rect 41140 16750 41150 16810
rect 41210 16750 41220 16810
rect 41140 14410 41220 16750
rect 41570 16810 42270 16820
rect 41570 16750 41580 16810
rect 41640 16754 42270 16810
rect 41640 16750 41660 16754
rect 41570 16720 41660 16750
rect 41694 16720 41760 16754
rect 41794 16720 41860 16754
rect 41894 16720 41960 16754
rect 41994 16720 42060 16754
rect 42094 16720 42160 16754
rect 42194 16720 42270 16754
rect 41570 16654 42270 16720
rect 41570 16620 41660 16654
rect 41694 16620 41760 16654
rect 41794 16620 41860 16654
rect 41894 16620 41960 16654
rect 41994 16620 42060 16654
rect 42094 16620 42160 16654
rect 42194 16620 42270 16654
rect 41570 16554 42270 16620
rect 41570 16520 41660 16554
rect 41694 16520 41760 16554
rect 41794 16520 41860 16554
rect 41894 16520 41960 16554
rect 41994 16520 42060 16554
rect 42094 16520 42160 16554
rect 42194 16520 42270 16554
rect 41570 15770 42270 16520
rect 42930 17054 43630 17130
rect 42930 17020 43020 17054
rect 43054 17020 43120 17054
rect 43154 17020 43220 17054
rect 43254 17020 43320 17054
rect 43354 17020 43420 17054
rect 43454 17020 43520 17054
rect 43554 17020 43630 17054
rect 42930 16954 43630 17020
rect 42930 16920 43020 16954
rect 43054 16920 43120 16954
rect 43154 16920 43220 16954
rect 43254 16920 43320 16954
rect 43354 16920 43420 16954
rect 43454 16920 43520 16954
rect 43554 16920 43630 16954
rect 42930 16854 43630 16920
rect 42930 16820 43020 16854
rect 43054 16820 43120 16854
rect 43154 16820 43220 16854
rect 43254 16820 43320 16854
rect 43354 16820 43420 16854
rect 43454 16820 43520 16854
rect 43554 16820 43630 16854
rect 42930 16810 43630 16820
rect 42930 16754 43250 16810
rect 43310 16754 43630 16810
rect 42930 16720 43020 16754
rect 43054 16720 43120 16754
rect 43154 16720 43220 16754
rect 43310 16750 43320 16754
rect 43254 16720 43320 16750
rect 43354 16720 43420 16754
rect 43454 16720 43520 16754
rect 43554 16720 43630 16754
rect 42930 16654 43630 16720
rect 42930 16620 43020 16654
rect 43054 16620 43120 16654
rect 43154 16620 43220 16654
rect 43254 16620 43320 16654
rect 43354 16620 43420 16654
rect 43454 16620 43520 16654
rect 43554 16620 43630 16654
rect 42930 16554 43630 16620
rect 42930 16520 43020 16554
rect 43054 16520 43120 16554
rect 43154 16520 43220 16554
rect 43254 16520 43320 16554
rect 43354 16520 43420 16554
rect 43454 16520 43520 16554
rect 43554 16520 43630 16554
rect 42930 16430 43630 16520
rect 44290 17054 44990 17790
rect 44290 17020 44380 17054
rect 44414 17020 44480 17054
rect 44514 17020 44580 17054
rect 44614 17020 44680 17054
rect 44714 17020 44780 17054
rect 44814 17020 44880 17054
rect 44914 17020 44990 17054
rect 44290 16954 44990 17020
rect 44290 16920 44380 16954
rect 44414 16920 44480 16954
rect 44514 16920 44580 16954
rect 44614 16920 44680 16954
rect 44714 16920 44780 16954
rect 44814 16920 44880 16954
rect 44914 16920 44990 16954
rect 44290 16854 44990 16920
rect 44290 16820 44380 16854
rect 44414 16820 44480 16854
rect 44514 16820 44580 16854
rect 44614 16820 44680 16854
rect 44714 16820 44780 16854
rect 44814 16820 44880 16854
rect 44914 16820 44990 16854
rect 47550 17047 47668 17059
rect 44290 16754 44990 16820
rect 44290 16720 44380 16754
rect 44414 16720 44480 16754
rect 44514 16720 44580 16754
rect 44614 16720 44680 16754
rect 44714 16720 44780 16754
rect 44814 16720 44880 16754
rect 44914 16720 44990 16754
rect 44290 16654 44990 16720
rect 44290 16620 44380 16654
rect 44414 16620 44480 16654
rect 44514 16620 44580 16654
rect 44614 16620 44680 16654
rect 44714 16620 44780 16654
rect 44814 16620 44880 16654
rect 44914 16620 44990 16654
rect 44290 16554 44990 16620
rect 44290 16520 44380 16554
rect 44414 16520 44480 16554
rect 44514 16520 44580 16554
rect 44614 16520 44680 16554
rect 44714 16520 44780 16554
rect 44814 16520 44880 16554
rect 44914 16520 44990 16554
rect 44290 15770 44990 16520
rect 41570 15694 44990 15770
rect 41570 15660 41660 15694
rect 41694 15660 41760 15694
rect 41794 15660 41860 15694
rect 41894 15660 41960 15694
rect 41994 15660 42060 15694
rect 42094 15660 42160 15694
rect 42194 15660 43020 15694
rect 43054 15660 43120 15694
rect 43154 15660 43220 15694
rect 43254 15660 43320 15694
rect 43354 15660 43420 15694
rect 43454 15660 43520 15694
rect 43554 15660 44380 15694
rect 44414 15660 44480 15694
rect 44514 15660 44580 15694
rect 44614 15660 44680 15694
rect 44714 15660 44780 15694
rect 44814 15660 44880 15694
rect 44914 15660 44990 15694
rect 41570 15594 44990 15660
rect 41570 15560 41660 15594
rect 41694 15560 41760 15594
rect 41794 15560 41860 15594
rect 41894 15560 41960 15594
rect 41994 15560 42060 15594
rect 42094 15560 42160 15594
rect 42194 15560 43020 15594
rect 43054 15560 43120 15594
rect 43154 15560 43220 15594
rect 43254 15560 43320 15594
rect 43354 15560 43420 15594
rect 43454 15560 43520 15594
rect 43554 15560 44380 15594
rect 44414 15560 44480 15594
rect 44514 15560 44580 15594
rect 44614 15560 44680 15594
rect 44714 15560 44780 15594
rect 44814 15560 44880 15594
rect 44914 15560 44990 15594
rect 41570 15494 44990 15560
rect 41570 15460 41660 15494
rect 41694 15460 41760 15494
rect 41794 15460 41860 15494
rect 41894 15460 41960 15494
rect 41994 15460 42060 15494
rect 42094 15460 42160 15494
rect 42194 15460 43020 15494
rect 43054 15460 43120 15494
rect 43154 15460 43220 15494
rect 43254 15460 43320 15494
rect 43354 15460 43420 15494
rect 43454 15460 43520 15494
rect 43554 15460 44380 15494
rect 44414 15460 44480 15494
rect 44514 15460 44580 15494
rect 44614 15460 44680 15494
rect 44714 15460 44780 15494
rect 44814 15460 44880 15494
rect 44914 15460 44990 15494
rect 41570 15394 44990 15460
rect 41570 15360 41660 15394
rect 41694 15360 41760 15394
rect 41794 15360 41860 15394
rect 41894 15360 41960 15394
rect 41994 15360 42060 15394
rect 42094 15360 42160 15394
rect 42194 15360 43020 15394
rect 43054 15360 43120 15394
rect 43154 15360 43220 15394
rect 43254 15360 43320 15394
rect 43354 15360 43420 15394
rect 43454 15360 43520 15394
rect 43554 15360 44380 15394
rect 44414 15360 44480 15394
rect 44514 15360 44580 15394
rect 44614 15360 44680 15394
rect 44714 15360 44780 15394
rect 44814 15360 44880 15394
rect 44914 15360 44990 15394
rect 41570 15294 44990 15360
rect 41570 15260 41660 15294
rect 41694 15260 41760 15294
rect 41794 15260 41860 15294
rect 41894 15260 41960 15294
rect 41994 15260 42060 15294
rect 42094 15260 42160 15294
rect 42194 15260 43020 15294
rect 43054 15260 43120 15294
rect 43154 15260 43220 15294
rect 43254 15260 43320 15294
rect 43354 15260 43420 15294
rect 43454 15260 43520 15294
rect 43554 15260 44380 15294
rect 44414 15260 44480 15294
rect 44514 15260 44580 15294
rect 44614 15260 44680 15294
rect 44714 15260 44780 15294
rect 44814 15260 44880 15294
rect 44914 15260 44990 15294
rect 41570 15194 44990 15260
rect 41570 15160 41660 15194
rect 41694 15160 41760 15194
rect 41794 15160 41860 15194
rect 41894 15160 41960 15194
rect 41994 15160 42060 15194
rect 42094 15160 42160 15194
rect 42194 15160 43020 15194
rect 43054 15160 43120 15194
rect 43154 15160 43220 15194
rect 43254 15160 43320 15194
rect 43354 15160 43420 15194
rect 43454 15160 43520 15194
rect 43554 15160 44380 15194
rect 44414 15160 44480 15194
rect 44514 15160 44580 15194
rect 44614 15160 44680 15194
rect 44714 15160 44780 15194
rect 44814 15160 44880 15194
rect 44914 15160 44990 15194
rect 41570 15070 44990 15160
rect 45340 16810 45420 16820
rect 45340 16750 45350 16810
rect 45410 16750 45420 16810
rect 45340 14800 45420 16750
rect 45340 14740 45350 14800
rect 45410 14740 45420 14800
rect 45340 14730 45420 14740
rect 46000 16700 46080 16720
rect 46000 16310 46020 16700
rect 46060 16310 46080 16700
rect 47550 16650 47556 17047
rect 47662 16650 47668 17047
rect 47550 16638 47668 16650
rect 46000 14800 46080 16310
rect 46780 16367 46860 16390
rect 46780 15970 46800 16367
rect 46838 15970 46860 16367
rect 46350 15350 46590 15370
rect 46350 15290 46360 15350
rect 46420 15290 46440 15350
rect 46500 15290 46520 15350
rect 46580 15290 46590 15350
rect 46000 14740 46010 14800
rect 46070 14740 46080 14800
rect 46000 14730 46080 14740
rect 46240 14800 46320 14810
rect 46240 14740 46250 14800
rect 46310 14740 46320 14800
rect 46240 14730 46320 14740
rect 44580 14720 45020 14730
rect 44580 14660 44590 14720
rect 44650 14660 44680 14720
rect 44740 14660 44770 14720
rect 44830 14660 44860 14720
rect 44920 14660 44950 14720
rect 45010 14660 45020 14720
rect 41140 14350 41150 14410
rect 41210 14350 41220 14410
rect 41140 14340 41220 14350
rect 41540 14402 41980 14420
rect 41540 14350 41560 14402
rect 41960 14350 41980 14402
rect 41540 14340 41980 14350
rect 44580 14402 45020 14660
rect 44580 14398 44600 14402
rect 44580 14360 44599 14398
rect 44580 14350 44600 14360
rect 45000 14350 45020 14402
rect 44580 14340 45020 14350
rect 46150 14410 46230 14420
rect 46150 14350 46160 14410
rect 46220 14350 46230 14410
rect 46150 14340 46230 14350
rect 41030 13920 41040 13980
rect 41100 13920 41110 13980
rect 41030 13910 41110 13920
rect 45470 13850 45550 13860
rect 41080 13810 41160 13820
rect 41080 13750 41090 13810
rect 41150 13750 41160 13810
rect 41080 13740 41160 13750
rect 45470 13790 45480 13850
rect 45540 13790 45550 13850
rect 45470 13770 45550 13790
rect 45470 13710 45480 13770
rect 45540 13710 45550 13770
rect 45470 13700 45550 13710
rect 41160 13640 41240 13650
rect 41160 13580 41170 13640
rect 41230 13580 41240 13640
rect 41160 13570 41240 13580
rect 41320 13640 41400 13650
rect 41320 13580 41330 13640
rect 41390 13580 41400 13640
rect 41320 13570 41400 13580
rect 41480 13640 41560 13650
rect 41480 13580 41490 13640
rect 41550 13580 41560 13640
rect 41480 13570 41560 13580
rect 41640 13640 41720 13650
rect 41640 13580 41650 13640
rect 41710 13580 41720 13640
rect 41640 13570 41720 13580
rect 41800 13640 41880 13650
rect 41800 13580 41810 13640
rect 41870 13580 41880 13640
rect 41800 13570 41880 13580
rect 41960 13640 42040 13650
rect 41960 13580 41970 13640
rect 42030 13580 42040 13640
rect 41960 13570 42040 13580
rect 42120 13640 42200 13650
rect 42120 13580 42130 13640
rect 42190 13580 42200 13640
rect 42120 13570 42200 13580
rect 42280 13640 42360 13650
rect 42280 13580 42290 13640
rect 42350 13580 42360 13640
rect 42280 13570 42360 13580
rect 42440 13640 42520 13650
rect 42440 13580 42450 13640
rect 42510 13580 42520 13640
rect 42440 13570 42520 13580
rect 42600 13640 42680 13650
rect 42600 13580 42610 13640
rect 42670 13580 42680 13640
rect 42600 13570 42680 13580
rect 42760 13640 42840 13650
rect 42760 13580 42770 13640
rect 42830 13580 42840 13640
rect 42760 13570 42840 13580
rect 42920 13640 43000 13650
rect 42920 13580 42930 13640
rect 42990 13580 43000 13640
rect 42920 13570 43000 13580
rect 43080 13640 43160 13650
rect 43080 13580 43090 13640
rect 43150 13580 43160 13640
rect 43080 13570 43160 13580
rect 43240 13640 43320 13650
rect 43240 13580 43250 13640
rect 43310 13580 43320 13640
rect 43240 13570 43320 13580
rect 43400 13640 43480 13650
rect 43400 13580 43410 13640
rect 43470 13580 43480 13640
rect 43400 13570 43480 13580
rect 43560 13640 43640 13650
rect 43560 13580 43570 13640
rect 43630 13580 43640 13640
rect 43560 13570 43640 13580
rect 43720 13640 43800 13650
rect 43720 13580 43730 13640
rect 43790 13580 43800 13640
rect 43720 13570 43800 13580
rect 43880 13640 43960 13650
rect 43880 13580 43890 13640
rect 43950 13580 43960 13640
rect 43880 13570 43960 13580
rect 44040 13640 44120 13650
rect 44040 13580 44050 13640
rect 44110 13580 44120 13640
rect 44040 13570 44120 13580
rect 44200 13640 44280 13650
rect 44200 13580 44210 13640
rect 44270 13580 44280 13640
rect 44200 13570 44280 13580
rect 44360 13640 44440 13650
rect 44360 13580 44370 13640
rect 44430 13580 44440 13640
rect 44360 13570 44440 13580
rect 44520 13640 44600 13650
rect 44520 13580 44530 13640
rect 44590 13580 44600 13640
rect 44520 13570 44600 13580
rect 44680 13640 44760 13650
rect 44680 13580 44690 13640
rect 44750 13580 44760 13640
rect 44680 13570 44760 13580
rect 44840 13640 44920 13650
rect 44840 13580 44850 13640
rect 44910 13580 44920 13640
rect 44840 13570 44920 13580
rect 45000 13640 45080 13650
rect 45000 13580 45010 13640
rect 45070 13580 45080 13640
rect 45000 13570 45080 13580
rect 45160 13640 45240 13650
rect 45160 13580 45170 13640
rect 45230 13580 45240 13640
rect 45160 13570 45240 13580
rect 41900 13530 41980 13540
rect 41900 13470 41910 13530
rect 41970 13470 41980 13530
rect 41900 13450 41980 13470
rect 41900 13390 41910 13450
rect 41970 13390 41980 13450
rect 41900 13370 41980 13390
rect 41900 13310 41910 13370
rect 41970 13310 41980 13370
rect 41900 13300 41980 13310
rect 43160 13530 43400 13540
rect 43160 13470 43170 13530
rect 43230 13470 43250 13530
rect 43310 13470 43330 13530
rect 43390 13470 43400 13530
rect 43160 13450 43400 13470
rect 43160 13390 43170 13450
rect 43230 13390 43250 13450
rect 43310 13390 43330 13450
rect 43390 13390 43400 13450
rect 43160 13370 43400 13390
rect 43160 13310 43170 13370
rect 43230 13310 43250 13370
rect 43310 13310 43330 13370
rect 43390 13310 43400 13370
rect 40740 12760 40820 12780
rect 40740 12720 40760 12760
rect 40800 12720 40820 12760
rect 43070 12750 43130 12770
rect 40740 12460 40820 12720
rect 40920 12730 41000 12740
rect 40920 12670 40930 12730
rect 40990 12670 41000 12730
rect 40920 12650 41000 12670
rect 40920 12590 40930 12650
rect 40990 12590 41000 12650
rect 40920 12570 41000 12590
rect 40920 12510 40930 12570
rect 40990 12510 41000 12570
rect 40920 12500 41000 12510
rect 41160 12730 41240 12740
rect 41160 12670 41170 12730
rect 41230 12670 41240 12730
rect 41160 12650 41240 12670
rect 41160 12590 41170 12650
rect 41230 12590 41240 12650
rect 41160 12570 41240 12590
rect 41160 12510 41170 12570
rect 41230 12510 41240 12570
rect 41160 12500 41240 12510
rect 41400 12730 41480 12740
rect 41400 12670 41410 12730
rect 41470 12670 41480 12730
rect 41400 12650 41480 12670
rect 41400 12590 41410 12650
rect 41470 12590 41480 12650
rect 41400 12570 41480 12590
rect 41400 12510 41410 12570
rect 41470 12510 41480 12570
rect 41400 12500 41480 12510
rect 41640 12730 41720 12740
rect 41640 12670 41650 12730
rect 41710 12670 41720 12730
rect 41640 12650 41720 12670
rect 41640 12590 41650 12650
rect 41710 12590 41720 12650
rect 41640 12570 41720 12590
rect 41640 12510 41650 12570
rect 41710 12510 41720 12570
rect 41640 12500 41720 12510
rect 42280 12730 42360 12740
rect 42280 12670 42290 12730
rect 42350 12670 42360 12730
rect 42280 12650 42360 12670
rect 42280 12590 42290 12650
rect 42350 12590 42360 12650
rect 42280 12570 42360 12590
rect 42280 12510 42290 12570
rect 42350 12510 42360 12570
rect 42280 12500 42360 12510
rect 42520 12730 42600 12740
rect 42520 12670 42530 12730
rect 42590 12670 42600 12730
rect 42520 12650 42600 12670
rect 42520 12590 42530 12650
rect 42590 12590 42600 12650
rect 42520 12570 42600 12590
rect 42520 12510 42530 12570
rect 42590 12510 42600 12570
rect 42520 12500 42600 12510
rect 42760 12730 42840 12740
rect 42760 12670 42770 12730
rect 42830 12670 42840 12730
rect 42760 12650 42840 12670
rect 42760 12590 42770 12650
rect 42830 12590 42840 12650
rect 42760 12570 42840 12590
rect 42760 12510 42770 12570
rect 42830 12510 42840 12570
rect 42760 12500 42840 12510
rect 43070 12710 43080 12750
rect 43120 12710 43130 12750
rect 40740 12400 40750 12460
rect 40810 12400 40820 12460
rect 40740 12390 40820 12400
rect 41490 12460 41570 12470
rect 41490 12400 41500 12460
rect 41560 12400 41570 12460
rect 41490 12390 41570 12400
rect 41710 12460 41790 12470
rect 41710 12400 41720 12460
rect 41780 12400 41790 12460
rect 41710 12390 41790 12400
rect 41970 12460 42050 12470
rect 41970 12400 41980 12460
rect 42040 12400 42050 12460
rect 41970 12390 42050 12400
rect 42190 12460 42270 12470
rect 42190 12400 42200 12460
rect 42260 12400 42270 12460
rect 42190 12390 42270 12400
rect 42450 12460 42530 12470
rect 42450 12400 42460 12460
rect 42520 12400 42530 12460
rect 42450 12390 42530 12400
rect 41431 12350 41489 12360
rect 41431 12298 41433 12350
rect 41485 12298 41489 12350
rect 41431 12290 41489 12298
rect 41520 12250 41550 12390
rect 41730 12250 41760 12390
rect 41791 12350 41849 12360
rect 41791 12298 41793 12350
rect 41845 12298 41849 12350
rect 41791 12290 41849 12298
rect 41911 12350 41969 12360
rect 41911 12298 41913 12350
rect 41965 12298 41969 12350
rect 41911 12290 41969 12298
rect 42000 12250 42030 12390
rect 42210 12250 42240 12390
rect 42271 12350 42329 12360
rect 42271 12298 42273 12350
rect 42325 12298 42329 12350
rect 42271 12290 42329 12298
rect 42391 12350 42449 12360
rect 42391 12298 42393 12350
rect 42445 12298 42449 12350
rect 42391 12290 42449 12298
rect 42480 12250 42510 12390
rect 42800 12330 42880 12340
rect 42800 12270 42810 12330
rect 42870 12270 42880 12330
rect 42800 12250 42880 12270
rect 41370 12230 41430 12250
rect 41370 12190 41380 12230
rect 41420 12190 41430 12230
rect 41370 11920 41430 12190
rect 41490 12230 41550 12250
rect 41490 12190 41500 12230
rect 41540 12190 41550 12230
rect 41490 12170 41550 12190
rect 41610 12230 41670 12250
rect 41610 12190 41620 12230
rect 41660 12190 41670 12230
rect 41610 12170 41670 12190
rect 41730 12230 41790 12250
rect 41730 12190 41740 12230
rect 41780 12190 41790 12230
rect 41730 12170 41790 12190
rect 41850 12230 41910 12250
rect 41850 12190 41860 12230
rect 41900 12190 41910 12230
rect 41850 12170 41910 12190
rect 41970 12230 42030 12250
rect 41970 12190 41980 12230
rect 42020 12190 42030 12230
rect 41970 12170 42030 12190
rect 42090 12230 42150 12250
rect 42090 12190 42100 12230
rect 42140 12190 42150 12230
rect 42090 12170 42150 12190
rect 42210 12230 42270 12250
rect 42210 12190 42220 12230
rect 42260 12190 42270 12230
rect 42210 12170 42270 12190
rect 42330 12230 42390 12250
rect 42330 12190 42340 12230
rect 42380 12190 42390 12230
rect 42330 12170 42390 12190
rect 42450 12230 42510 12250
rect 42450 12190 42460 12230
rect 42500 12190 42510 12230
rect 42450 12170 42510 12190
rect 42570 12230 42630 12250
rect 42570 12190 42580 12230
rect 42620 12190 42630 12230
rect 42570 12170 42630 12190
rect 42800 12190 42810 12250
rect 42870 12190 42880 12250
rect 42800 12170 42880 12190
rect 41532 12122 41590 12130
rect 41532 12070 41536 12122
rect 41588 12070 41590 12122
rect 41532 12060 41590 12070
rect 41620 12030 41660 12170
rect 41690 12122 41748 12130
rect 41690 12070 41694 12122
rect 41746 12070 41748 12122
rect 41690 12060 41748 12070
rect 41600 12020 41680 12030
rect 41600 11960 41610 12020
rect 41670 11960 41680 12020
rect 41360 11910 41440 11920
rect 41360 11850 41370 11910
rect 41430 11850 41440 11910
rect 40620 11640 40780 11650
rect 40620 11580 40630 11640
rect 40690 11580 40710 11640
rect 40770 11580 40780 11640
rect 40620 11570 40780 11580
rect 41120 11640 41200 11650
rect 41120 11580 41130 11640
rect 41190 11580 41200 11640
rect 41120 11570 41200 11580
rect 41360 11640 41440 11850
rect 41360 11580 41370 11640
rect 41430 11580 41440 11640
rect 41360 11570 41440 11580
rect 40710 11520 40770 11570
rect 40710 11480 40720 11520
rect 40760 11480 40770 11520
rect 40710 11460 40770 11480
rect 40880 11520 40960 11530
rect 40880 11460 40890 11520
rect 40950 11460 40960 11520
rect 40880 11450 40960 11460
rect 40530 11390 40590 11410
rect 40530 11350 40540 11390
rect 40580 11350 40590 11390
rect 40530 11290 40590 11350
rect 40530 11250 40540 11290
rect 40580 11250 40590 11290
rect 40530 11170 40590 11250
rect 40650 11390 40710 11410
rect 40650 11350 40660 11390
rect 40700 11350 40710 11390
rect 40650 11290 40710 11350
rect 40650 11250 40660 11290
rect 40700 11250 40710 11290
rect 40650 11190 40710 11250
rect 40770 11390 40830 11410
rect 40770 11350 40780 11390
rect 40820 11350 40830 11390
rect 40770 11290 40830 11350
rect 40770 11250 40780 11290
rect 40820 11250 40830 11290
rect 40530 11130 40540 11170
rect 40580 11130 40590 11170
rect 40530 11080 40590 11130
rect 40640 11180 40720 11190
rect 40640 11120 40650 11180
rect 40710 11120 40720 11180
rect 40640 11110 40720 11120
rect 40770 11080 40830 11250
rect 40890 11390 40950 11450
rect 40890 11350 40900 11390
rect 40940 11350 40950 11390
rect 40890 11290 40950 11350
rect 40890 11250 40900 11290
rect 40940 11250 40950 11290
rect 40890 11230 40950 11250
rect 41010 11390 41070 11410
rect 41010 11350 41020 11390
rect 41060 11350 41070 11390
rect 41010 11290 41070 11350
rect 41010 11250 41020 11290
rect 41060 11250 41070 11290
rect 41010 11080 41070 11250
rect 41130 11390 41190 11570
rect 41370 11510 41430 11570
rect 41370 11470 41380 11510
rect 41420 11470 41430 11510
rect 41370 11450 41430 11470
rect 41600 11520 41680 11960
rect 41860 11920 41900 12170
rect 42014 12122 42072 12130
rect 42014 12070 42018 12122
rect 42070 12070 42072 12122
rect 42014 12060 42072 12070
rect 42100 12030 42140 12170
rect 42168 12122 42226 12130
rect 42168 12070 42172 12122
rect 42224 12070 42226 12122
rect 42168 12060 42226 12070
rect 42080 12020 42160 12030
rect 42080 11960 42090 12020
rect 42150 11960 42160 12020
rect 42080 11950 42160 11960
rect 42340 11920 42380 12170
rect 42492 12122 42550 12130
rect 42492 12070 42496 12122
rect 42548 12070 42550 12122
rect 42492 12060 42550 12070
rect 42580 12030 42620 12170
rect 42800 12110 42810 12170
rect 42870 12110 42880 12170
rect 42800 12100 42880 12110
rect 42560 12020 42640 12030
rect 42560 11960 42570 12020
rect 42630 11960 42640 12020
rect 42560 11950 42640 11960
rect 41840 11910 41920 11920
rect 41840 11850 41850 11910
rect 41910 11850 41920 11910
rect 41840 11840 41920 11850
rect 42320 11910 42400 11920
rect 42320 11850 42330 11910
rect 42390 11850 42400 11910
rect 42320 11840 42400 11850
rect 41840 11640 41920 11650
rect 41840 11580 41850 11640
rect 41910 11580 41920 11640
rect 41840 11570 41920 11580
rect 42080 11640 42160 11650
rect 42080 11580 42090 11640
rect 42150 11580 42160 11640
rect 42080 11570 42160 11580
rect 42560 11640 42640 11650
rect 42560 11580 42570 11640
rect 42630 11580 42640 11640
rect 42560 11570 42640 11580
rect 42740 11640 42820 11650
rect 42740 11580 42750 11640
rect 42810 11580 42820 11640
rect 42740 11570 42820 11580
rect 41600 11460 41610 11520
rect 41670 11460 41680 11520
rect 41600 11450 41680 11460
rect 41130 11350 41140 11390
rect 41180 11350 41190 11390
rect 41130 11290 41190 11350
rect 41130 11250 41140 11290
rect 41180 11250 41190 11290
rect 41130 11230 41190 11250
rect 41250 11390 41310 11410
rect 41250 11350 41260 11390
rect 41300 11350 41310 11390
rect 41250 11290 41310 11350
rect 41250 11250 41260 11290
rect 41300 11250 41310 11290
rect 41250 11080 41310 11250
rect 41370 11390 41430 11410
rect 41370 11350 41380 11390
rect 41420 11350 41430 11390
rect 41370 11290 41430 11350
rect 41370 11250 41380 11290
rect 41420 11250 41430 11290
rect 41370 11190 41430 11250
rect 41490 11390 41550 11410
rect 41490 11350 41500 11390
rect 41540 11350 41550 11390
rect 41490 11290 41550 11350
rect 41490 11250 41500 11290
rect 41540 11250 41550 11290
rect 41360 11180 41440 11190
rect 41360 11120 41370 11180
rect 41430 11120 41440 11180
rect 41360 11110 41440 11120
rect 41490 11080 41550 11250
rect 41610 11390 41670 11450
rect 41610 11350 41620 11390
rect 41660 11350 41670 11390
rect 41610 11290 41670 11350
rect 41610 11250 41620 11290
rect 41660 11250 41670 11290
rect 41610 11230 41670 11250
rect 41730 11390 41790 11410
rect 41730 11350 41740 11390
rect 41780 11350 41790 11390
rect 41730 11290 41790 11350
rect 41730 11250 41740 11290
rect 41780 11250 41790 11290
rect 41730 11080 41790 11250
rect 41850 11390 41910 11570
rect 42090 11510 42150 11570
rect 42090 11470 42100 11510
rect 42140 11470 42150 11510
rect 42090 11450 42150 11470
rect 42320 11520 42400 11530
rect 42320 11460 42330 11520
rect 42390 11460 42400 11520
rect 42320 11450 42400 11460
rect 41850 11350 41860 11390
rect 41900 11350 41910 11390
rect 41850 11290 41910 11350
rect 41850 11250 41860 11290
rect 41900 11250 41910 11290
rect 41850 11230 41910 11250
rect 41970 11390 42030 11410
rect 41970 11350 41980 11390
rect 42020 11350 42030 11390
rect 41970 11290 42030 11350
rect 41970 11250 41980 11290
rect 42020 11250 42030 11290
rect 41970 11080 42030 11250
rect 42090 11390 42150 11410
rect 42090 11350 42100 11390
rect 42140 11350 42150 11390
rect 42090 11290 42150 11350
rect 42090 11250 42100 11290
rect 42140 11250 42150 11290
rect 42090 11190 42150 11250
rect 42210 11390 42270 11410
rect 42210 11350 42220 11390
rect 42260 11350 42270 11390
rect 42210 11290 42270 11350
rect 42210 11250 42220 11290
rect 42260 11250 42270 11290
rect 42080 11180 42160 11190
rect 42080 11120 42090 11180
rect 42150 11120 42160 11180
rect 42080 11110 42160 11120
rect 42210 11080 42270 11250
rect 42330 11390 42390 11450
rect 42330 11350 42340 11390
rect 42380 11350 42390 11390
rect 42330 11290 42390 11350
rect 42330 11250 42340 11290
rect 42380 11250 42390 11290
rect 42330 11230 42390 11250
rect 42450 11390 42510 11410
rect 42450 11350 42460 11390
rect 42500 11350 42510 11390
rect 42450 11290 42510 11350
rect 42450 11250 42460 11290
rect 42500 11250 42510 11290
rect 42450 11080 42510 11250
rect 42570 11390 42630 11570
rect 42750 11510 42810 11570
rect 42750 11470 42760 11510
rect 42800 11470 42810 11510
rect 42750 11450 42810 11470
rect 42570 11350 42580 11390
rect 42620 11350 42630 11390
rect 42570 11290 42630 11350
rect 42570 11250 42580 11290
rect 42620 11250 42630 11290
rect 42570 11230 42630 11250
rect 42690 11390 42750 11410
rect 42690 11350 42700 11390
rect 42740 11350 42750 11390
rect 42690 11290 42750 11350
rect 42690 11250 42700 11290
rect 42740 11250 42750 11290
rect 42690 11080 42750 11250
rect 42810 11390 42870 11410
rect 42810 11350 42820 11390
rect 42860 11350 42870 11390
rect 42810 11290 42870 11350
rect 42810 11250 42820 11290
rect 42860 11250 42870 11290
rect 42810 11190 42870 11250
rect 42930 11390 42990 11410
rect 42930 11350 42940 11390
rect 42980 11350 42990 11390
rect 42930 11290 42990 11350
rect 42930 11250 42940 11290
rect 42980 11250 42990 11290
rect 42800 11180 42880 11190
rect 42800 11120 42810 11180
rect 42870 11120 42880 11180
rect 42800 11110 42880 11120
rect 42930 11170 42990 11250
rect 43070 11190 43130 12710
rect 43160 12330 43400 13310
rect 44580 13530 44660 13540
rect 44580 13470 44590 13530
rect 44650 13470 44660 13530
rect 44580 13450 44660 13470
rect 44580 13390 44590 13450
rect 44650 13390 44660 13450
rect 44580 13370 44660 13390
rect 44580 13310 44590 13370
rect 44650 13310 44660 13370
rect 44580 13300 44660 13310
rect 45750 13240 45810 13260
rect 45750 13200 45760 13240
rect 45800 13200 45810 13240
rect 45750 13140 45810 13200
rect 45750 13100 45760 13140
rect 45800 13100 45810 13140
rect 45750 13040 45810 13100
rect 45750 13000 45760 13040
rect 45800 13000 45810 13040
rect 45750 12940 45810 13000
rect 45750 12900 45760 12940
rect 45800 12900 45810 12940
rect 45750 12840 45810 12900
rect 45750 12800 45760 12840
rect 45800 12800 45810 12840
rect 43160 12270 43170 12330
rect 43230 12270 43250 12330
rect 43310 12270 43330 12330
rect 43390 12270 43400 12330
rect 43160 12250 43400 12270
rect 43160 12190 43170 12250
rect 43230 12190 43250 12250
rect 43310 12190 43330 12250
rect 43390 12190 43400 12250
rect 43160 12170 43400 12190
rect 43160 12110 43170 12170
rect 43230 12110 43250 12170
rect 43310 12110 43330 12170
rect 43390 12110 43400 12170
rect 43160 12100 43400 12110
rect 43430 12750 43490 12770
rect 43430 12710 43440 12750
rect 43480 12710 43490 12750
rect 43430 11190 43490 12710
rect 43720 12730 43800 12740
rect 43720 12670 43730 12730
rect 43790 12670 43800 12730
rect 43720 12650 43800 12670
rect 43720 12590 43730 12650
rect 43790 12590 43800 12650
rect 43720 12570 43800 12590
rect 43720 12510 43730 12570
rect 43790 12510 43800 12570
rect 43720 12500 43800 12510
rect 43960 12730 44040 12740
rect 43960 12670 43970 12730
rect 44030 12670 44040 12730
rect 43960 12650 44040 12670
rect 43960 12590 43970 12650
rect 44030 12590 44040 12650
rect 43960 12570 44040 12590
rect 43960 12510 43970 12570
rect 44030 12510 44040 12570
rect 43960 12500 44040 12510
rect 44200 12730 44280 12740
rect 44200 12670 44210 12730
rect 44270 12670 44280 12730
rect 44200 12650 44280 12670
rect 44200 12590 44210 12650
rect 44270 12590 44280 12650
rect 44200 12570 44280 12590
rect 44200 12510 44210 12570
rect 44270 12510 44280 12570
rect 44200 12500 44280 12510
rect 44840 12730 44920 12740
rect 44840 12670 44850 12730
rect 44910 12670 44920 12730
rect 44840 12650 44920 12670
rect 44840 12590 44850 12650
rect 44910 12590 44920 12650
rect 44840 12570 44920 12590
rect 44840 12510 44850 12570
rect 44910 12510 44920 12570
rect 44840 12500 44920 12510
rect 45080 12730 45160 12740
rect 45080 12670 45090 12730
rect 45150 12670 45160 12730
rect 45080 12650 45160 12670
rect 45080 12590 45090 12650
rect 45150 12590 45160 12650
rect 45080 12570 45160 12590
rect 45080 12510 45090 12570
rect 45150 12510 45160 12570
rect 45080 12500 45160 12510
rect 45320 12730 45400 12740
rect 45320 12670 45330 12730
rect 45390 12670 45400 12730
rect 45320 12650 45400 12670
rect 45320 12590 45330 12650
rect 45390 12590 45400 12650
rect 45320 12570 45400 12590
rect 45320 12510 45330 12570
rect 45390 12510 45400 12570
rect 45320 12500 45400 12510
rect 45560 12730 45640 12740
rect 45560 12670 45570 12730
rect 45630 12670 45640 12730
rect 45560 12650 45640 12670
rect 45560 12590 45570 12650
rect 45630 12590 45640 12650
rect 45560 12570 45640 12590
rect 45560 12510 45570 12570
rect 45630 12510 45640 12570
rect 45560 12500 45640 12510
rect 45750 12470 45810 12800
rect 44030 12460 44110 12470
rect 44030 12400 44040 12460
rect 44100 12400 44110 12460
rect 44030 12390 44110 12400
rect 44290 12460 44370 12470
rect 44290 12400 44300 12460
rect 44360 12400 44370 12460
rect 44290 12390 44370 12400
rect 44510 12460 44590 12470
rect 44510 12400 44520 12460
rect 44580 12400 44590 12460
rect 44510 12390 44590 12400
rect 44770 12460 44850 12470
rect 44770 12400 44780 12460
rect 44840 12400 44850 12460
rect 44770 12390 44850 12400
rect 44990 12460 45070 12470
rect 44990 12400 45000 12460
rect 45060 12400 45070 12460
rect 44990 12390 45070 12400
rect 45740 12460 45820 12470
rect 45740 12400 45750 12460
rect 45810 12400 45820 12460
rect 45740 12390 45820 12400
rect 43680 12330 43760 12340
rect 43680 12270 43690 12330
rect 43750 12270 43760 12330
rect 43680 12250 43760 12270
rect 44050 12250 44080 12390
rect 44111 12350 44169 12360
rect 44111 12298 44115 12350
rect 44167 12298 44169 12350
rect 44111 12290 44169 12298
rect 44231 12350 44289 12360
rect 44231 12298 44235 12350
rect 44287 12298 44289 12350
rect 44231 12290 44289 12298
rect 44320 12250 44350 12390
rect 44530 12250 44560 12390
rect 44591 12350 44649 12360
rect 44591 12298 44595 12350
rect 44647 12298 44649 12350
rect 44591 12290 44649 12298
rect 44711 12350 44769 12360
rect 44711 12298 44715 12350
rect 44767 12298 44769 12350
rect 44711 12290 44769 12298
rect 44800 12250 44830 12390
rect 45010 12250 45040 12390
rect 46170 12360 46210 14340
rect 45071 12350 45129 12360
rect 45071 12298 45075 12350
rect 45127 12298 45129 12350
rect 45071 12290 45129 12298
rect 46150 12350 46230 12360
rect 46150 12290 46160 12350
rect 46220 12290 46230 12350
rect 46150 12280 46230 12290
rect 43680 12190 43690 12250
rect 43750 12190 43760 12250
rect 43680 12170 43760 12190
rect 43930 12230 43990 12250
rect 43930 12190 43940 12230
rect 43980 12190 43990 12230
rect 43930 12170 43990 12190
rect 44050 12230 44110 12250
rect 44050 12190 44060 12230
rect 44100 12190 44110 12230
rect 44050 12170 44110 12190
rect 44170 12230 44230 12250
rect 44170 12190 44180 12230
rect 44220 12190 44230 12230
rect 44170 12170 44230 12190
rect 44290 12230 44350 12250
rect 44290 12190 44300 12230
rect 44340 12190 44350 12230
rect 44290 12170 44350 12190
rect 44410 12230 44470 12250
rect 44410 12190 44420 12230
rect 44460 12190 44470 12230
rect 44410 12170 44470 12190
rect 44530 12230 44590 12250
rect 44530 12190 44540 12230
rect 44580 12190 44590 12230
rect 44530 12170 44590 12190
rect 44650 12230 44710 12250
rect 44650 12190 44660 12230
rect 44700 12190 44710 12230
rect 44650 12170 44710 12190
rect 44770 12230 44830 12250
rect 44770 12190 44780 12230
rect 44820 12190 44830 12230
rect 44770 12170 44830 12190
rect 44890 12230 44950 12250
rect 44890 12190 44900 12230
rect 44940 12190 44950 12230
rect 44890 12170 44950 12190
rect 45010 12230 45070 12250
rect 45010 12190 45020 12230
rect 45060 12190 45070 12230
rect 45010 12170 45070 12190
rect 45130 12230 45190 12250
rect 45130 12190 45140 12230
rect 45180 12190 45190 12230
rect 43680 12110 43690 12170
rect 43750 12110 43760 12170
rect 43680 12100 43760 12110
rect 43940 12030 43980 12170
rect 44010 12122 44068 12130
rect 44010 12070 44012 12122
rect 44064 12070 44068 12122
rect 44010 12060 44068 12070
rect 43920 12020 44000 12030
rect 43920 11960 43930 12020
rect 43990 11960 44000 12020
rect 43920 11950 44000 11960
rect 44180 11920 44220 12170
rect 44334 12122 44392 12130
rect 44334 12070 44336 12122
rect 44388 12070 44392 12122
rect 44334 12060 44392 12070
rect 44420 12030 44460 12170
rect 44488 12122 44546 12130
rect 44488 12070 44490 12122
rect 44542 12070 44546 12122
rect 44488 12060 44546 12070
rect 44400 12020 44480 12030
rect 44400 11960 44410 12020
rect 44470 11960 44480 12020
rect 44400 11950 44480 11960
rect 44660 11920 44700 12170
rect 44812 12122 44870 12130
rect 44812 12070 44814 12122
rect 44866 12070 44870 12122
rect 44812 12060 44870 12070
rect 44900 12030 44940 12170
rect 44970 12122 45028 12130
rect 44970 12070 44972 12122
rect 45024 12070 45028 12122
rect 44970 12060 45028 12070
rect 44880 12020 44960 12030
rect 44880 11960 44890 12020
rect 44950 11960 44960 12020
rect 44160 11910 44240 11920
rect 44160 11850 44170 11910
rect 44230 11850 44240 11910
rect 44160 11840 44240 11850
rect 44640 11910 44720 11920
rect 44640 11850 44650 11910
rect 44710 11850 44720 11910
rect 44640 11840 44720 11850
rect 43740 11800 43820 11810
rect 43740 11740 43750 11800
rect 43810 11740 43820 11800
rect 43740 11720 43820 11740
rect 43740 11660 43750 11720
rect 43810 11660 43820 11720
rect 43740 11640 43820 11660
rect 43740 11580 43750 11640
rect 43810 11580 43820 11640
rect 43740 11570 43820 11580
rect 43920 11800 44000 11810
rect 43920 11740 43930 11800
rect 43990 11740 44000 11800
rect 43920 11720 44000 11740
rect 43920 11660 43930 11720
rect 43990 11660 44000 11720
rect 43920 11640 44000 11660
rect 43920 11580 43930 11640
rect 43990 11580 44000 11640
rect 43920 11570 44000 11580
rect 44160 11800 44240 11810
rect 44160 11740 44170 11800
rect 44230 11740 44240 11800
rect 44160 11720 44240 11740
rect 44160 11660 44170 11720
rect 44230 11660 44240 11720
rect 44160 11640 44240 11660
rect 44160 11580 44170 11640
rect 44230 11580 44240 11640
rect 44160 11570 44240 11580
rect 44400 11800 44480 11810
rect 44400 11740 44410 11800
rect 44470 11740 44480 11800
rect 44400 11720 44480 11740
rect 44400 11660 44410 11720
rect 44470 11660 44480 11720
rect 44400 11640 44480 11660
rect 44400 11580 44410 11640
rect 44470 11580 44480 11640
rect 44400 11570 44480 11580
rect 44640 11800 44720 11810
rect 44640 11740 44650 11800
rect 44710 11740 44720 11800
rect 44640 11720 44720 11740
rect 44640 11660 44650 11720
rect 44710 11660 44720 11720
rect 44640 11640 44720 11660
rect 44640 11580 44650 11640
rect 44710 11580 44720 11640
rect 44640 11570 44720 11580
rect 43750 11510 43810 11570
rect 43750 11470 43760 11510
rect 43800 11470 43810 11510
rect 43750 11450 43810 11470
rect 43570 11390 43630 11410
rect 43570 11350 43580 11390
rect 43620 11350 43630 11390
rect 43570 11290 43630 11350
rect 43570 11250 43580 11290
rect 43620 11250 43630 11290
rect 42930 11130 42940 11170
rect 42980 11130 42990 11170
rect 42930 11080 42990 11130
rect 43060 11180 43140 11190
rect 43060 11120 43070 11180
rect 43130 11120 43140 11180
rect 43060 11110 43140 11120
rect 43420 11180 43500 11190
rect 43420 11120 43430 11180
rect 43490 11120 43500 11180
rect 40520 11070 40600 11080
rect 40520 11010 40530 11070
rect 40590 11010 40600 11070
rect 40520 10990 40600 11010
rect 40520 10930 40530 10990
rect 40590 10930 40600 10990
rect 40520 10910 40600 10930
rect 40520 10850 40530 10910
rect 40590 10850 40600 10910
rect 40520 10840 40600 10850
rect 40760 11070 40840 11080
rect 40760 11010 40770 11070
rect 40830 11010 40840 11070
rect 40760 10990 40840 11010
rect 40760 10930 40770 10990
rect 40830 10930 40840 10990
rect 40760 10910 40840 10930
rect 40760 10850 40770 10910
rect 40830 10850 40840 10910
rect 40760 10840 40840 10850
rect 41000 11070 41080 11080
rect 41000 11010 41010 11070
rect 41070 11010 41080 11070
rect 41000 10990 41080 11010
rect 41000 10930 41010 10990
rect 41070 10930 41080 10990
rect 41000 10910 41080 10930
rect 41000 10850 41010 10910
rect 41070 10850 41080 10910
rect 41000 10840 41080 10850
rect 41240 11070 41320 11080
rect 41240 11010 41250 11070
rect 41310 11010 41320 11070
rect 41240 10990 41320 11010
rect 41240 10930 41250 10990
rect 41310 10930 41320 10990
rect 41240 10910 41320 10930
rect 41240 10850 41250 10910
rect 41310 10850 41320 10910
rect 41240 10840 41320 10850
rect 41480 11070 41560 11080
rect 41480 11010 41490 11070
rect 41550 11010 41560 11070
rect 41480 10990 41560 11010
rect 41480 10930 41490 10990
rect 41550 10930 41560 10990
rect 41480 10910 41560 10930
rect 41480 10850 41490 10910
rect 41550 10850 41560 10910
rect 41480 10840 41560 10850
rect 41720 11070 41800 11080
rect 41720 11010 41730 11070
rect 41790 11010 41800 11070
rect 41720 10990 41800 11010
rect 41720 10930 41730 10990
rect 41790 10930 41800 10990
rect 41720 10910 41800 10930
rect 41720 10850 41730 10910
rect 41790 10850 41800 10910
rect 41720 10840 41800 10850
rect 41960 11070 42040 11080
rect 41960 11010 41970 11070
rect 42030 11010 42040 11070
rect 41960 10990 42040 11010
rect 41960 10930 41970 10990
rect 42030 10930 42040 10990
rect 41960 10910 42040 10930
rect 41960 10850 41970 10910
rect 42030 10850 42040 10910
rect 41960 10840 42040 10850
rect 42200 11070 42280 11080
rect 42200 11010 42210 11070
rect 42270 11010 42280 11070
rect 42200 10990 42280 11010
rect 42200 10930 42210 10990
rect 42270 10930 42280 10990
rect 42200 10910 42280 10930
rect 42200 10850 42210 10910
rect 42270 10850 42280 10910
rect 42200 10840 42280 10850
rect 42440 11070 42520 11080
rect 42440 11010 42450 11070
rect 42510 11010 42520 11070
rect 42440 10990 42520 11010
rect 42440 10930 42450 10990
rect 42510 10930 42520 10990
rect 42440 10910 42520 10930
rect 42440 10850 42450 10910
rect 42510 10850 42520 10910
rect 42440 10840 42520 10850
rect 42680 11070 42760 11080
rect 42680 11010 42690 11070
rect 42750 11010 42760 11070
rect 42680 10990 42760 11010
rect 42680 10930 42690 10990
rect 42750 10930 42760 10990
rect 42680 10910 42760 10930
rect 42680 10850 42690 10910
rect 42750 10850 42760 10910
rect 42680 10840 42760 10850
rect 42920 11070 43000 11080
rect 42920 11010 42930 11070
rect 42990 11010 43000 11070
rect 42920 10990 43000 11010
rect 42920 10930 42930 10990
rect 42990 10930 43000 10990
rect 42920 10910 43000 10930
rect 42920 10850 42930 10910
rect 42990 10850 43000 10910
rect 42920 10840 43000 10850
rect 41800 10800 41880 10810
rect 41800 10740 41810 10800
rect 41870 10740 41880 10800
rect 41800 10730 41880 10740
rect 43240 10800 43320 10810
rect 43240 10740 43250 10800
rect 43310 10740 43320 10800
rect 43240 10730 43320 10740
rect 41630 10230 41690 10250
rect 41630 10190 41640 10230
rect 41680 10190 41690 10230
rect 41630 10130 41690 10190
rect 41630 10090 41640 10130
rect 41680 10090 41690 10130
rect 41630 10030 41690 10090
rect 41630 9990 41640 10030
rect 41680 9990 41690 10030
rect 41630 9930 41690 9990
rect 41630 9890 41640 9930
rect 41680 9890 41690 9930
rect 41630 9830 41690 9890
rect 41630 9790 41640 9830
rect 41680 9790 41690 9830
rect 41630 9730 41690 9790
rect 41630 9690 41640 9730
rect 41680 9690 41690 9730
rect 41630 9670 41690 9690
rect 41810 10230 41870 10730
rect 42160 10690 42240 10700
rect 42160 10630 42170 10690
rect 42230 10630 42240 10690
rect 42160 10620 42240 10630
rect 41900 10360 41970 10370
rect 41960 10300 41970 10360
rect 41900 10290 41970 10300
rect 42070 10360 42150 10370
rect 42070 10300 42080 10360
rect 42140 10300 42150 10360
rect 42070 10290 42150 10300
rect 42180 10250 42220 10620
rect 42520 10580 42600 10590
rect 42520 10520 42530 10580
rect 42590 10520 42600 10580
rect 42520 10510 42600 10520
rect 42250 10360 42330 10370
rect 42250 10300 42260 10360
rect 42320 10300 42330 10360
rect 42250 10290 42330 10300
rect 42430 10360 42510 10370
rect 42430 10300 42440 10360
rect 42500 10300 42510 10360
rect 42430 10290 42510 10300
rect 42540 10250 42580 10510
rect 42880 10470 42960 10480
rect 42880 10410 42890 10470
rect 42950 10410 42960 10470
rect 42880 10400 42960 10410
rect 42610 10360 42690 10370
rect 42610 10300 42620 10360
rect 42680 10300 42690 10360
rect 42610 10290 42690 10300
rect 42790 10360 42870 10370
rect 42790 10300 42800 10360
rect 42860 10300 42870 10360
rect 42790 10290 42870 10300
rect 42900 10250 42940 10400
rect 42970 10360 43050 10370
rect 42970 10300 42980 10360
rect 43040 10300 43050 10360
rect 42970 10290 43050 10300
rect 43150 10360 43220 10370
rect 43150 10300 43160 10360
rect 43150 10290 43220 10300
rect 41810 10190 41820 10230
rect 41860 10190 41870 10230
rect 41810 10130 41870 10190
rect 41810 10090 41820 10130
rect 41860 10090 41870 10130
rect 41810 10030 41870 10090
rect 41810 9990 41820 10030
rect 41860 9990 41870 10030
rect 41810 9930 41870 9990
rect 41810 9890 41820 9930
rect 41860 9890 41870 9930
rect 41810 9830 41870 9890
rect 41810 9790 41820 9830
rect 41860 9790 41870 9830
rect 41810 9730 41870 9790
rect 41810 9690 41820 9730
rect 41860 9690 41870 9730
rect 41810 9670 41870 9690
rect 41990 10230 42050 10250
rect 41990 10190 42000 10230
rect 42040 10190 42050 10230
rect 41990 10130 42050 10190
rect 41990 10090 42000 10130
rect 42040 10090 42050 10130
rect 41990 10030 42050 10090
rect 41990 9990 42000 10030
rect 42040 9990 42050 10030
rect 41990 9930 42050 9990
rect 41990 9890 42000 9930
rect 42040 9890 42050 9930
rect 41990 9830 42050 9890
rect 41990 9790 42000 9830
rect 42040 9790 42050 9830
rect 41990 9730 42050 9790
rect 41990 9690 42000 9730
rect 42040 9690 42050 9730
rect 41990 9670 42050 9690
rect 42170 10230 42230 10250
rect 42170 10190 42180 10230
rect 42220 10190 42230 10230
rect 42170 10130 42230 10190
rect 42170 10090 42180 10130
rect 42220 10090 42230 10130
rect 42170 10030 42230 10090
rect 42170 9990 42180 10030
rect 42220 9990 42230 10030
rect 42170 9930 42230 9990
rect 42170 9890 42180 9930
rect 42220 9890 42230 9930
rect 42170 9830 42230 9890
rect 42170 9790 42180 9830
rect 42220 9790 42230 9830
rect 42170 9730 42230 9790
rect 42170 9690 42180 9730
rect 42220 9690 42230 9730
rect 42170 9670 42230 9690
rect 42350 10230 42410 10250
rect 42350 10190 42360 10230
rect 42400 10190 42410 10230
rect 42350 10130 42410 10190
rect 42350 10090 42360 10130
rect 42400 10090 42410 10130
rect 42350 10030 42410 10090
rect 42350 9990 42360 10030
rect 42400 9990 42410 10030
rect 42350 9930 42410 9990
rect 42350 9890 42360 9930
rect 42400 9890 42410 9930
rect 42350 9830 42410 9890
rect 42350 9790 42360 9830
rect 42400 9790 42410 9830
rect 42350 9730 42410 9790
rect 42350 9690 42360 9730
rect 42400 9690 42410 9730
rect 42350 9670 42410 9690
rect 42530 10230 42590 10250
rect 42530 10190 42540 10230
rect 42580 10190 42590 10230
rect 42530 10130 42590 10190
rect 42530 10090 42540 10130
rect 42580 10090 42590 10130
rect 42530 10030 42590 10090
rect 42530 9990 42540 10030
rect 42580 9990 42590 10030
rect 42530 9930 42590 9990
rect 42530 9890 42540 9930
rect 42580 9890 42590 9930
rect 42530 9830 42590 9890
rect 42530 9790 42540 9830
rect 42580 9790 42590 9830
rect 42530 9730 42590 9790
rect 42530 9690 42540 9730
rect 42580 9690 42590 9730
rect 42530 9670 42590 9690
rect 42710 10230 42770 10250
rect 42710 10190 42720 10230
rect 42760 10190 42770 10230
rect 42710 10130 42770 10190
rect 42710 10090 42720 10130
rect 42760 10090 42770 10130
rect 42710 10030 42770 10090
rect 42710 9990 42720 10030
rect 42760 9990 42770 10030
rect 42710 9930 42770 9990
rect 42710 9890 42720 9930
rect 42760 9890 42770 9930
rect 42710 9830 42770 9890
rect 42710 9790 42720 9830
rect 42760 9790 42770 9830
rect 42710 9730 42770 9790
rect 42710 9690 42720 9730
rect 42760 9690 42770 9730
rect 42710 9670 42770 9690
rect 42890 10230 42950 10250
rect 42890 10190 42900 10230
rect 42940 10190 42950 10230
rect 42890 10130 42950 10190
rect 42890 10090 42900 10130
rect 42940 10090 42950 10130
rect 42890 10030 42950 10090
rect 42890 9990 42900 10030
rect 42940 9990 42950 10030
rect 42890 9930 42950 9990
rect 42890 9890 42900 9930
rect 42940 9890 42950 9930
rect 42890 9830 42950 9890
rect 42890 9790 42900 9830
rect 42940 9790 42950 9830
rect 42890 9730 42950 9790
rect 42890 9690 42900 9730
rect 42940 9690 42950 9730
rect 42890 9670 42950 9690
rect 43070 10230 43130 10250
rect 43070 10190 43080 10230
rect 43120 10190 43130 10230
rect 43070 10130 43130 10190
rect 43070 10090 43080 10130
rect 43120 10090 43130 10130
rect 43070 10030 43130 10090
rect 43070 9990 43080 10030
rect 43120 9990 43130 10030
rect 43070 9930 43130 9990
rect 43070 9890 43080 9930
rect 43120 9890 43130 9930
rect 43070 9830 43130 9890
rect 43070 9790 43080 9830
rect 43120 9790 43130 9830
rect 43070 9730 43130 9790
rect 43070 9690 43080 9730
rect 43120 9690 43130 9730
rect 43070 9670 43130 9690
rect 43250 10230 43310 10730
rect 43420 10370 43500 11120
rect 43570 11170 43630 11250
rect 43690 11390 43750 11410
rect 43690 11350 43700 11390
rect 43740 11350 43750 11390
rect 43690 11290 43750 11350
rect 43690 11250 43700 11290
rect 43740 11250 43750 11290
rect 43690 11190 43750 11250
rect 43810 11390 43870 11410
rect 43810 11350 43820 11390
rect 43860 11350 43870 11390
rect 43810 11290 43870 11350
rect 43810 11250 43820 11290
rect 43860 11250 43870 11290
rect 43570 11130 43580 11170
rect 43620 11130 43630 11170
rect 43570 11080 43630 11130
rect 43680 11180 43760 11190
rect 43680 11120 43690 11180
rect 43750 11120 43760 11180
rect 43680 11110 43760 11120
rect 43810 11080 43870 11250
rect 43930 11390 43990 11570
rect 44160 11520 44240 11530
rect 44160 11460 44170 11520
rect 44230 11460 44240 11520
rect 44160 11450 44240 11460
rect 44410 11510 44470 11570
rect 44410 11470 44420 11510
rect 44460 11470 44470 11510
rect 44410 11450 44470 11470
rect 43930 11350 43940 11390
rect 43980 11350 43990 11390
rect 43930 11290 43990 11350
rect 43930 11250 43940 11290
rect 43980 11250 43990 11290
rect 43930 11230 43990 11250
rect 44050 11390 44110 11410
rect 44050 11350 44060 11390
rect 44100 11350 44110 11390
rect 44050 11290 44110 11350
rect 44050 11250 44060 11290
rect 44100 11250 44110 11290
rect 44050 11080 44110 11250
rect 44170 11390 44230 11450
rect 44170 11350 44180 11390
rect 44220 11350 44230 11390
rect 44170 11290 44230 11350
rect 44170 11250 44180 11290
rect 44220 11250 44230 11290
rect 44170 11230 44230 11250
rect 44290 11390 44350 11410
rect 44290 11350 44300 11390
rect 44340 11350 44350 11390
rect 44290 11290 44350 11350
rect 44290 11250 44300 11290
rect 44340 11250 44350 11290
rect 44290 11080 44350 11250
rect 44410 11390 44470 11410
rect 44410 11350 44420 11390
rect 44460 11350 44470 11390
rect 44410 11290 44470 11350
rect 44410 11250 44420 11290
rect 44460 11250 44470 11290
rect 44410 11190 44470 11250
rect 44530 11390 44590 11410
rect 44530 11350 44540 11390
rect 44580 11350 44590 11390
rect 44530 11290 44590 11350
rect 44530 11250 44540 11290
rect 44580 11250 44590 11290
rect 44400 11180 44480 11190
rect 44400 11120 44410 11180
rect 44470 11120 44480 11180
rect 44400 11110 44480 11120
rect 44530 11080 44590 11250
rect 44650 11390 44710 11570
rect 44880 11520 44960 11960
rect 45130 11920 45190 12190
rect 45120 11910 45200 11920
rect 45120 11850 45130 11910
rect 45190 11850 45200 11910
rect 45120 11800 45200 11850
rect 45120 11740 45130 11800
rect 45190 11740 45200 11800
rect 45120 11720 45200 11740
rect 45120 11660 45130 11720
rect 45190 11660 45200 11720
rect 45120 11640 45200 11660
rect 45120 11580 45130 11640
rect 45190 11580 45200 11640
rect 45120 11570 45200 11580
rect 45360 11800 45440 11810
rect 45360 11740 45370 11800
rect 45430 11740 45440 11800
rect 45360 11720 45440 11740
rect 45360 11660 45370 11720
rect 45430 11660 45440 11720
rect 45360 11640 45440 11660
rect 45360 11580 45370 11640
rect 45430 11580 45440 11640
rect 45360 11570 45440 11580
rect 45780 11800 45860 11810
rect 45780 11740 45790 11800
rect 45850 11740 45860 11800
rect 45780 11720 45860 11740
rect 45780 11660 45790 11720
rect 45850 11660 45860 11720
rect 45780 11640 45860 11660
rect 45780 11580 45790 11640
rect 45850 11580 45860 11640
rect 45780 11570 45860 11580
rect 44880 11460 44890 11520
rect 44950 11460 44960 11520
rect 44880 11450 44960 11460
rect 45130 11510 45190 11570
rect 45130 11470 45140 11510
rect 45180 11470 45190 11510
rect 45130 11450 45190 11470
rect 44650 11350 44660 11390
rect 44700 11350 44710 11390
rect 44650 11290 44710 11350
rect 44650 11250 44660 11290
rect 44700 11250 44710 11290
rect 44650 11230 44710 11250
rect 44770 11390 44830 11410
rect 44770 11350 44780 11390
rect 44820 11350 44830 11390
rect 44770 11290 44830 11350
rect 44770 11250 44780 11290
rect 44820 11250 44830 11290
rect 44770 11080 44830 11250
rect 44890 11390 44950 11450
rect 44890 11350 44900 11390
rect 44940 11350 44950 11390
rect 44890 11290 44950 11350
rect 44890 11250 44900 11290
rect 44940 11250 44950 11290
rect 44890 11230 44950 11250
rect 45010 11390 45070 11410
rect 45010 11350 45020 11390
rect 45060 11350 45070 11390
rect 45010 11290 45070 11350
rect 45010 11250 45020 11290
rect 45060 11250 45070 11290
rect 45010 11080 45070 11250
rect 45130 11390 45190 11410
rect 45130 11350 45140 11390
rect 45180 11350 45190 11390
rect 45130 11290 45190 11350
rect 45130 11250 45140 11290
rect 45180 11250 45190 11290
rect 45130 11190 45190 11250
rect 45250 11390 45310 11410
rect 45250 11350 45260 11390
rect 45300 11350 45310 11390
rect 45250 11290 45310 11350
rect 45250 11250 45260 11290
rect 45300 11250 45310 11290
rect 45120 11180 45200 11190
rect 45120 11120 45130 11180
rect 45190 11120 45200 11180
rect 45120 11110 45200 11120
rect 45250 11080 45310 11250
rect 45370 11390 45430 11570
rect 45600 11520 45680 11530
rect 45600 11460 45610 11520
rect 45670 11460 45680 11520
rect 45790 11520 45850 11570
rect 45790 11480 45800 11520
rect 45840 11480 45850 11520
rect 45790 11460 45850 11480
rect 45600 11450 45680 11460
rect 45370 11350 45380 11390
rect 45420 11350 45430 11390
rect 45370 11290 45430 11350
rect 45370 11250 45380 11290
rect 45420 11250 45430 11290
rect 45370 11230 45430 11250
rect 45490 11390 45550 11410
rect 45490 11350 45500 11390
rect 45540 11350 45550 11390
rect 45490 11290 45550 11350
rect 45490 11250 45500 11290
rect 45540 11250 45550 11290
rect 45490 11080 45550 11250
rect 45610 11390 45670 11450
rect 45610 11350 45620 11390
rect 45660 11350 45670 11390
rect 45610 11290 45670 11350
rect 45610 11250 45620 11290
rect 45660 11250 45670 11290
rect 45610 11230 45670 11250
rect 45730 11390 45790 11410
rect 45730 11350 45740 11390
rect 45780 11350 45790 11390
rect 45730 11290 45790 11350
rect 45730 11250 45740 11290
rect 45780 11250 45790 11290
rect 45730 11080 45790 11250
rect 45850 11390 45910 11410
rect 45850 11350 45860 11390
rect 45900 11350 45910 11390
rect 45850 11290 45910 11350
rect 45850 11250 45860 11290
rect 45900 11250 45910 11290
rect 45850 11190 45910 11250
rect 45970 11390 46030 11410
rect 45970 11350 45980 11390
rect 46020 11350 46030 11390
rect 45970 11290 46030 11350
rect 45970 11250 45980 11290
rect 46020 11250 46030 11290
rect 45840 11180 45920 11190
rect 45840 11120 45850 11180
rect 45910 11120 45920 11180
rect 43560 11070 43640 11080
rect 43560 11010 43570 11070
rect 43630 11010 43640 11070
rect 43560 10990 43640 11010
rect 43560 10930 43570 10990
rect 43630 10930 43640 10990
rect 43560 10910 43640 10930
rect 43560 10850 43570 10910
rect 43630 10850 43640 10910
rect 43560 10840 43640 10850
rect 43800 11070 43880 11080
rect 43800 11010 43810 11070
rect 43870 11010 43880 11070
rect 43800 10990 43880 11010
rect 43800 10930 43810 10990
rect 43870 10930 43880 10990
rect 43800 10910 43880 10930
rect 43800 10850 43810 10910
rect 43870 10850 43880 10910
rect 43800 10840 43880 10850
rect 44040 11070 44120 11080
rect 44040 11010 44050 11070
rect 44110 11010 44120 11070
rect 44040 10990 44120 11010
rect 44040 10930 44050 10990
rect 44110 10930 44120 10990
rect 44040 10910 44120 10930
rect 44040 10850 44050 10910
rect 44110 10850 44120 10910
rect 44040 10840 44120 10850
rect 44280 11070 44360 11080
rect 44280 11010 44290 11070
rect 44350 11010 44360 11070
rect 44280 10990 44360 11010
rect 44280 10930 44290 10990
rect 44350 10930 44360 10990
rect 44280 10910 44360 10930
rect 44280 10850 44290 10910
rect 44350 10850 44360 10910
rect 44280 10840 44360 10850
rect 44520 11070 44600 11080
rect 44520 11010 44530 11070
rect 44590 11010 44600 11070
rect 44520 10990 44600 11010
rect 44520 10930 44530 10990
rect 44590 10930 44600 10990
rect 44520 10910 44600 10930
rect 44520 10850 44530 10910
rect 44590 10850 44600 10910
rect 44520 10840 44600 10850
rect 44760 11070 44840 11080
rect 44760 11010 44770 11070
rect 44830 11010 44840 11070
rect 44760 10990 44840 11010
rect 44760 10930 44770 10990
rect 44830 10930 44840 10990
rect 44760 10910 44840 10930
rect 44760 10850 44770 10910
rect 44830 10850 44840 10910
rect 44760 10840 44840 10850
rect 45000 11070 45080 11080
rect 45000 11010 45010 11070
rect 45070 11010 45080 11070
rect 45000 10990 45080 11010
rect 45000 10930 45010 10990
rect 45070 10930 45080 10990
rect 45000 10910 45080 10930
rect 45000 10850 45010 10910
rect 45070 10850 45080 10910
rect 45000 10840 45080 10850
rect 45240 11070 45320 11080
rect 45240 11010 45250 11070
rect 45310 11010 45320 11070
rect 45240 10990 45320 11010
rect 45240 10930 45250 10990
rect 45310 10930 45320 10990
rect 45240 10910 45320 10930
rect 45240 10850 45250 10910
rect 45310 10850 45320 10910
rect 45240 10840 45320 10850
rect 45480 11070 45560 11080
rect 45480 11010 45490 11070
rect 45550 11010 45560 11070
rect 45480 10990 45560 11010
rect 45480 10930 45490 10990
rect 45550 10930 45560 10990
rect 45480 10910 45560 10930
rect 45480 10850 45490 10910
rect 45550 10850 45560 10910
rect 45480 10840 45560 10850
rect 45720 11070 45800 11080
rect 45720 11010 45730 11070
rect 45790 11010 45800 11070
rect 45720 10990 45800 11010
rect 45720 10930 45730 10990
rect 45790 10930 45800 10990
rect 45720 10910 45800 10930
rect 45720 10850 45730 10910
rect 45790 10850 45800 10910
rect 45720 10840 45800 10850
rect 44680 10800 44760 10810
rect 44680 10740 44690 10800
rect 44750 10740 44760 10800
rect 44680 10730 44760 10740
rect 44320 10690 44400 10700
rect 44320 10630 44330 10690
rect 44390 10630 44400 10690
rect 44320 10620 44400 10630
rect 43960 10580 44040 10590
rect 43960 10520 43970 10580
rect 44030 10520 44040 10580
rect 43960 10510 44040 10520
rect 43600 10470 43680 10480
rect 43600 10410 43610 10470
rect 43670 10410 43680 10470
rect 43600 10400 43680 10410
rect 43340 10360 43590 10370
rect 43400 10300 43430 10360
rect 43490 10300 43520 10360
rect 43580 10300 43590 10360
rect 43340 10290 43590 10300
rect 43620 10250 43660 10400
rect 43690 10360 43770 10370
rect 43690 10300 43700 10360
rect 43760 10300 43770 10360
rect 43690 10290 43770 10300
rect 43870 10360 43950 10370
rect 43870 10300 43880 10360
rect 43940 10300 43950 10360
rect 43870 10290 43950 10300
rect 43980 10250 44020 10510
rect 44050 10360 44130 10370
rect 44050 10300 44060 10360
rect 44120 10300 44130 10360
rect 44050 10290 44130 10300
rect 44230 10360 44310 10370
rect 44230 10300 44240 10360
rect 44300 10300 44310 10360
rect 44230 10290 44310 10300
rect 44340 10250 44380 10620
rect 44410 10360 44490 10370
rect 44410 10300 44420 10360
rect 44480 10300 44490 10360
rect 44410 10290 44490 10300
rect 44590 10360 44660 10370
rect 44590 10300 44600 10360
rect 44590 10290 44660 10300
rect 43250 10190 43260 10230
rect 43300 10190 43310 10230
rect 43250 10130 43310 10190
rect 43250 10090 43260 10130
rect 43300 10090 43310 10130
rect 43250 10030 43310 10090
rect 43250 9990 43260 10030
rect 43300 9990 43310 10030
rect 43250 9930 43310 9990
rect 43250 9890 43260 9930
rect 43300 9890 43310 9930
rect 43250 9830 43310 9890
rect 43250 9790 43260 9830
rect 43300 9790 43310 9830
rect 43250 9730 43310 9790
rect 43250 9690 43260 9730
rect 43300 9690 43310 9730
rect 43250 9670 43310 9690
rect 43430 10230 43490 10250
rect 43430 10190 43440 10230
rect 43480 10190 43490 10230
rect 43430 10130 43490 10190
rect 43430 10090 43440 10130
rect 43480 10090 43490 10130
rect 43430 10030 43490 10090
rect 43430 9990 43440 10030
rect 43480 9990 43490 10030
rect 43430 9930 43490 9990
rect 43430 9890 43440 9930
rect 43480 9890 43490 9930
rect 43430 9830 43490 9890
rect 43430 9790 43440 9830
rect 43480 9790 43490 9830
rect 43430 9730 43490 9790
rect 43430 9690 43440 9730
rect 43480 9690 43490 9730
rect 43430 9670 43490 9690
rect 43610 10230 43670 10250
rect 43610 10190 43620 10230
rect 43660 10190 43670 10230
rect 43610 10130 43670 10190
rect 43610 10090 43620 10130
rect 43660 10090 43670 10130
rect 43610 10030 43670 10090
rect 43610 9990 43620 10030
rect 43660 9990 43670 10030
rect 43610 9930 43670 9990
rect 43610 9890 43620 9930
rect 43660 9890 43670 9930
rect 43610 9830 43670 9890
rect 43610 9790 43620 9830
rect 43660 9790 43670 9830
rect 43610 9730 43670 9790
rect 43610 9690 43620 9730
rect 43660 9690 43670 9730
rect 43610 9670 43670 9690
rect 43790 10230 43850 10250
rect 43790 10190 43800 10230
rect 43840 10190 43850 10230
rect 43790 10130 43850 10190
rect 43790 10090 43800 10130
rect 43840 10090 43850 10130
rect 43790 10030 43850 10090
rect 43790 9990 43800 10030
rect 43840 9990 43850 10030
rect 43790 9930 43850 9990
rect 43790 9890 43800 9930
rect 43840 9890 43850 9930
rect 43790 9830 43850 9890
rect 43790 9790 43800 9830
rect 43840 9790 43850 9830
rect 43790 9730 43850 9790
rect 43790 9690 43800 9730
rect 43840 9690 43850 9730
rect 43790 9670 43850 9690
rect 43970 10230 44030 10250
rect 43970 10190 43980 10230
rect 44020 10190 44030 10230
rect 43970 10130 44030 10190
rect 43970 10090 43980 10130
rect 44020 10090 44030 10130
rect 43970 10030 44030 10090
rect 43970 9990 43980 10030
rect 44020 9990 44030 10030
rect 43970 9930 44030 9990
rect 43970 9890 43980 9930
rect 44020 9890 44030 9930
rect 43970 9830 44030 9890
rect 43970 9790 43980 9830
rect 44020 9790 44030 9830
rect 43970 9730 44030 9790
rect 43970 9690 43980 9730
rect 44020 9690 44030 9730
rect 43970 9670 44030 9690
rect 44150 10230 44210 10250
rect 44150 10190 44160 10230
rect 44200 10190 44210 10230
rect 44150 10130 44210 10190
rect 44150 10090 44160 10130
rect 44200 10090 44210 10130
rect 44150 10030 44210 10090
rect 44150 9990 44160 10030
rect 44200 9990 44210 10030
rect 44150 9930 44210 9990
rect 44150 9890 44160 9930
rect 44200 9890 44210 9930
rect 44150 9830 44210 9890
rect 44150 9790 44160 9830
rect 44200 9790 44210 9830
rect 44150 9730 44210 9790
rect 44150 9690 44160 9730
rect 44200 9690 44210 9730
rect 44150 9670 44210 9690
rect 44330 10230 44390 10250
rect 44330 10190 44340 10230
rect 44380 10190 44390 10230
rect 44330 10130 44390 10190
rect 44330 10090 44340 10130
rect 44380 10090 44390 10130
rect 44330 10030 44390 10090
rect 44330 9990 44340 10030
rect 44380 9990 44390 10030
rect 44330 9930 44390 9990
rect 44330 9890 44340 9930
rect 44380 9890 44390 9930
rect 44330 9830 44390 9890
rect 44330 9790 44340 9830
rect 44380 9790 44390 9830
rect 44330 9730 44390 9790
rect 44330 9690 44340 9730
rect 44380 9690 44390 9730
rect 44330 9670 44390 9690
rect 44510 10230 44570 10250
rect 44510 10190 44520 10230
rect 44560 10190 44570 10230
rect 44510 10130 44570 10190
rect 44510 10090 44520 10130
rect 44560 10090 44570 10130
rect 44510 10030 44570 10090
rect 44510 9990 44520 10030
rect 44560 9990 44570 10030
rect 44510 9930 44570 9990
rect 44510 9890 44520 9930
rect 44560 9890 44570 9930
rect 44510 9830 44570 9890
rect 44510 9790 44520 9830
rect 44560 9790 44570 9830
rect 44510 9730 44570 9790
rect 44510 9690 44520 9730
rect 44560 9690 44570 9730
rect 44510 9670 44570 9690
rect 44690 10230 44750 10730
rect 45710 10690 45790 10700
rect 45710 10630 45720 10690
rect 45780 10630 45790 10690
rect 45240 10580 45320 10590
rect 45240 10520 45250 10580
rect 45310 10520 45320 10580
rect 45240 10510 45320 10520
rect 44690 10190 44700 10230
rect 44740 10190 44750 10230
rect 44690 10130 44750 10190
rect 44690 10090 44700 10130
rect 44740 10090 44750 10130
rect 44690 10030 44750 10090
rect 44690 9990 44700 10030
rect 44740 9990 44750 10030
rect 44690 9930 44750 9990
rect 44690 9890 44700 9930
rect 44740 9890 44750 9930
rect 44690 9830 44750 9890
rect 44690 9790 44700 9830
rect 44740 9790 44750 9830
rect 44690 9730 44750 9790
rect 44690 9690 44700 9730
rect 44740 9690 44750 9730
rect 44690 9670 44750 9690
rect 44870 10230 44930 10250
rect 44870 10190 44880 10230
rect 44920 10190 44930 10230
rect 44870 10130 44930 10190
rect 44870 10090 44880 10130
rect 44920 10090 44930 10130
rect 44870 10030 44930 10090
rect 44870 9990 44880 10030
rect 44920 9990 44930 10030
rect 44870 9930 44930 9990
rect 44870 9890 44880 9930
rect 44920 9890 44930 9930
rect 44870 9830 44930 9890
rect 45260 9830 45300 10510
rect 45590 10160 45670 10170
rect 45590 10100 45600 10160
rect 45660 10100 45670 10160
rect 45590 10090 45670 10100
rect 45710 10150 45790 10630
rect 45840 10170 45920 11120
rect 45970 11170 46030 11250
rect 45970 11130 45980 11170
rect 46020 11130 46030 11170
rect 45970 11080 46030 11130
rect 45960 11070 46040 11080
rect 45960 11010 45970 11070
rect 46030 11010 46040 11070
rect 45960 10990 46040 11010
rect 45960 10930 45970 10990
rect 46030 10930 46040 10990
rect 45960 10910 46040 10930
rect 45960 10850 45970 10910
rect 46030 10850 46040 10910
rect 45960 10840 46040 10850
rect 46170 10480 46210 12280
rect 46260 12130 46300 14730
rect 46240 12120 46320 12130
rect 46240 12060 46250 12120
rect 46310 12060 46320 12120
rect 46240 12050 46320 12060
rect 46260 10590 46300 12050
rect 46350 11800 46590 15290
rect 46780 14090 46860 15970
rect 46780 14030 46790 14090
rect 46850 14030 46860 14090
rect 46780 14020 46860 14030
rect 46350 11740 46360 11800
rect 46420 11740 46440 11800
rect 46500 11740 46520 11800
rect 46580 11740 46590 11800
rect 46350 11720 46590 11740
rect 46350 11660 46360 11720
rect 46420 11660 46440 11720
rect 46500 11660 46520 11720
rect 46580 11660 46590 11720
rect 46350 11640 46590 11660
rect 46350 11580 46360 11640
rect 46420 11580 46440 11640
rect 46500 11580 46520 11640
rect 46580 11580 46590 11640
rect 46350 11570 46590 11580
rect 47570 11180 47650 16638
rect 47950 16050 48030 18050
rect 47950 15990 47960 16050
rect 48020 15990 48030 16050
rect 47950 15980 48030 15990
rect 48120 17450 48200 17460
rect 48120 17390 48130 17450
rect 48190 17390 48200 17450
rect 48120 13040 48200 17390
rect 48650 13980 48730 18070
rect 48780 16750 48880 16770
rect 48780 16690 48800 16750
rect 48860 16690 48880 16750
rect 48780 16670 48880 16690
rect 48780 15350 48880 15370
rect 48780 15290 48800 15350
rect 48860 15290 48880 15350
rect 48780 15270 48880 15290
rect 48650 13920 48660 13980
rect 48720 13920 48730 13980
rect 48650 13910 48730 13920
rect 47570 11120 47580 11180
rect 47640 11120 47650 11180
rect 47570 11110 47650 11120
rect 46240 10580 46320 10590
rect 46240 10520 46250 10580
rect 46310 10520 46320 10580
rect 46240 10510 46320 10520
rect 46150 10470 46230 10480
rect 46150 10410 46160 10470
rect 46220 10410 46230 10470
rect 46150 10400 46230 10410
rect 45710 10110 45730 10150
rect 45770 10110 45790 10150
rect 45710 10090 45790 10110
rect 45830 10160 45910 10170
rect 45830 10100 45840 10160
rect 45900 10100 45910 10160
rect 45830 10090 45910 10100
rect 45500 10030 45560 10050
rect 45500 9990 45510 10030
rect 45550 9990 45560 10030
rect 45500 9930 45560 9990
rect 45500 9890 45510 9930
rect 45550 9890 45560 9930
rect 45500 9830 45560 9890
rect 45610 10030 45670 10090
rect 45610 9990 45620 10030
rect 45660 9990 45670 10030
rect 45610 9930 45670 9990
rect 45610 9890 45620 9930
rect 45660 9890 45670 9930
rect 45610 9870 45670 9890
rect 45720 10030 45780 10050
rect 45720 9990 45730 10030
rect 45770 9990 45780 10030
rect 45720 9930 45780 9990
rect 45720 9890 45730 9930
rect 45770 9890 45780 9930
rect 45720 9830 45780 9890
rect 45830 10030 45890 10090
rect 45830 9990 45840 10030
rect 45880 9990 45890 10030
rect 45830 9930 45890 9990
rect 45830 9890 45840 9930
rect 45880 9890 45890 9930
rect 45830 9870 45890 9890
rect 45940 10030 46000 10050
rect 45940 9990 45950 10030
rect 45990 9990 46000 10030
rect 45940 9930 46000 9990
rect 45940 9890 45950 9930
rect 45990 9890 46000 9930
rect 45940 9830 46000 9890
rect 44870 9790 44880 9830
rect 44920 9790 44930 9830
rect 44870 9730 44930 9790
rect 45240 9820 45320 9830
rect 45240 9760 45250 9820
rect 45310 9760 45320 9820
rect 45240 9750 45320 9760
rect 45490 9810 45570 9830
rect 45490 9770 45510 9810
rect 45550 9770 45570 9810
rect 45490 9750 45570 9770
rect 45710 9820 45790 9830
rect 45710 9760 45720 9820
rect 45780 9760 45790 9820
rect 45710 9750 45790 9760
rect 45930 9810 46010 9830
rect 45930 9770 45950 9810
rect 45990 9770 46010 9810
rect 45930 9750 46010 9770
rect 44870 9690 44880 9730
rect 44920 9690 44930 9730
rect 44870 9670 44930 9690
rect 45500 9630 45560 9750
rect 45940 9630 46000 9750
rect 41620 9620 41700 9630
rect 41620 9560 41630 9620
rect 41690 9560 41700 9620
rect 41620 9540 41700 9560
rect 41620 9480 41630 9540
rect 41690 9480 41700 9540
rect 41620 9460 41700 9480
rect 41620 9400 41630 9460
rect 41690 9400 41700 9460
rect 41620 9390 41700 9400
rect 41980 9620 42060 9630
rect 41980 9560 41990 9620
rect 42050 9560 42060 9620
rect 41980 9540 42060 9560
rect 41980 9480 41990 9540
rect 42050 9480 42060 9540
rect 41980 9460 42060 9480
rect 41980 9400 41990 9460
rect 42050 9400 42060 9460
rect 41980 9390 42060 9400
rect 42340 9620 42420 9630
rect 42340 9560 42350 9620
rect 42410 9560 42420 9620
rect 42340 9540 42420 9560
rect 42340 9480 42350 9540
rect 42410 9480 42420 9540
rect 42340 9460 42420 9480
rect 42340 9400 42350 9460
rect 42410 9400 42420 9460
rect 42340 9390 42420 9400
rect 42700 9620 42780 9630
rect 42700 9560 42710 9620
rect 42770 9560 42780 9620
rect 42700 9540 42780 9560
rect 42700 9480 42710 9540
rect 42770 9480 42780 9540
rect 42700 9460 42780 9480
rect 42700 9400 42710 9460
rect 42770 9400 42780 9460
rect 42700 9390 42780 9400
rect 43060 9620 43140 9630
rect 43060 9560 43070 9620
rect 43130 9560 43140 9620
rect 43060 9540 43140 9560
rect 43060 9480 43070 9540
rect 43130 9480 43140 9540
rect 43060 9460 43140 9480
rect 43060 9400 43070 9460
rect 43130 9400 43140 9460
rect 43060 9390 43140 9400
rect 43420 9620 43500 9630
rect 43420 9560 43430 9620
rect 43490 9560 43500 9620
rect 43420 9540 43500 9560
rect 43420 9480 43430 9540
rect 43490 9480 43500 9540
rect 43420 9460 43500 9480
rect 43420 9400 43430 9460
rect 43490 9400 43500 9460
rect 43420 9390 43500 9400
rect 43780 9620 43860 9630
rect 43780 9560 43790 9620
rect 43850 9560 43860 9620
rect 43780 9540 43860 9560
rect 43780 9480 43790 9540
rect 43850 9480 43860 9540
rect 43780 9460 43860 9480
rect 43780 9400 43790 9460
rect 43850 9400 43860 9460
rect 43780 9390 43860 9400
rect 44140 9620 44220 9630
rect 44140 9560 44150 9620
rect 44210 9560 44220 9620
rect 44140 9540 44220 9560
rect 44140 9480 44150 9540
rect 44210 9480 44220 9540
rect 44140 9460 44220 9480
rect 44140 9400 44150 9460
rect 44210 9400 44220 9460
rect 44140 9390 44220 9400
rect 44500 9620 44580 9630
rect 44500 9560 44510 9620
rect 44570 9560 44580 9620
rect 44500 9540 44580 9560
rect 44500 9480 44510 9540
rect 44570 9480 44580 9540
rect 44500 9460 44580 9480
rect 44500 9400 44510 9460
rect 44570 9400 44580 9460
rect 44500 9390 44580 9400
rect 44860 9620 44940 9630
rect 44860 9560 44870 9620
rect 44930 9560 44940 9620
rect 44860 9540 44940 9560
rect 44860 9480 44870 9540
rect 44930 9480 44940 9540
rect 44860 9460 44940 9480
rect 44860 9400 44870 9460
rect 44930 9400 44940 9460
rect 44860 9390 44940 9400
rect 45490 9620 45570 9630
rect 45490 9560 45500 9620
rect 45560 9560 45570 9620
rect 45490 9540 45570 9560
rect 45490 9480 45500 9540
rect 45560 9480 45570 9540
rect 45490 9460 45570 9480
rect 45490 9400 45500 9460
rect 45560 9400 45570 9460
rect 45490 9390 45570 9400
rect 45930 9620 46010 9630
rect 45930 9560 45940 9620
rect 46000 9560 46010 9620
rect 45930 9540 46010 9560
rect 45930 9480 45940 9540
rect 46000 9480 46010 9540
rect 45930 9460 46010 9480
rect 45930 9400 45940 9460
rect 46000 9400 46010 9460
rect 45930 9390 46010 9400
rect 41806 9350 41864 9360
rect 41806 9298 41808 9350
rect 41860 9298 41864 9350
rect 41806 9290 41864 9298
rect 41916 9350 41974 9360
rect 41916 9298 41918 9350
rect 41970 9298 41974 9350
rect 41916 9290 41974 9298
rect 42026 9350 42084 9360
rect 42026 9298 42028 9350
rect 42080 9298 42084 9350
rect 42026 9290 42084 9298
rect 42136 9350 42194 9360
rect 42136 9298 42138 9350
rect 42190 9298 42194 9350
rect 42136 9290 42194 9298
rect 42246 9350 42304 9360
rect 42246 9298 42248 9350
rect 42300 9298 42304 9350
rect 42246 9290 42304 9298
rect 42356 9350 42414 9360
rect 42356 9298 42358 9350
rect 42410 9298 42414 9350
rect 42356 9290 42414 9298
rect 42466 9350 42524 9360
rect 42466 9298 42468 9350
rect 42520 9298 42524 9350
rect 42466 9290 42524 9298
rect 42576 9350 42634 9360
rect 42576 9298 42578 9350
rect 42630 9298 42634 9350
rect 42576 9290 42634 9298
rect 42686 9350 42744 9360
rect 42686 9298 42688 9350
rect 42740 9298 42744 9350
rect 42686 9290 42744 9298
rect 42796 9350 42854 9360
rect 42796 9298 42798 9350
rect 42850 9298 42854 9350
rect 42796 9290 42854 9298
rect 43706 9350 43764 9360
rect 43706 9298 43708 9350
rect 43760 9298 43764 9350
rect 43706 9290 43764 9298
rect 43816 9350 43874 9360
rect 43816 9298 43818 9350
rect 43870 9298 43874 9350
rect 43816 9290 43874 9298
rect 43926 9350 43984 9360
rect 43926 9298 43928 9350
rect 43980 9298 43984 9350
rect 43926 9290 43984 9298
rect 44036 9350 44094 9360
rect 44036 9298 44038 9350
rect 44090 9298 44094 9350
rect 44036 9290 44094 9298
rect 44146 9350 44204 9360
rect 44146 9298 44148 9350
rect 44200 9298 44204 9350
rect 44146 9290 44204 9298
rect 44256 9350 44314 9360
rect 44256 9298 44258 9350
rect 44310 9298 44314 9350
rect 44256 9290 44314 9298
rect 44366 9350 44424 9360
rect 44366 9298 44368 9350
rect 44420 9298 44424 9350
rect 44366 9290 44424 9298
rect 44476 9350 44534 9360
rect 44476 9298 44478 9350
rect 44530 9298 44534 9350
rect 44476 9290 44534 9298
rect 44586 9350 44644 9360
rect 44586 9298 44588 9350
rect 44640 9298 44644 9350
rect 44586 9290 44644 9298
rect 44696 9350 44754 9360
rect 44696 9298 44698 9350
rect 44750 9298 44754 9350
rect 44696 9290 44754 9298
rect 41560 9230 41700 9250
rect 41560 9190 41570 9230
rect 41610 9190 41650 9230
rect 41690 9190 41700 9230
rect 41560 9130 41700 9190
rect 41560 9090 41570 9130
rect 41610 9090 41650 9130
rect 41690 9090 41700 9130
rect 41560 9070 41700 9090
rect 41640 9030 41700 9070
rect 41750 9230 41810 9250
rect 41750 9190 41760 9230
rect 41800 9190 41810 9230
rect 41750 9130 41810 9190
rect 41750 9090 41760 9130
rect 41800 9090 41810 9130
rect 41630 9020 41710 9030
rect 41630 8960 41640 9020
rect 41700 8960 41710 9020
rect 41630 8950 41710 8960
rect 41750 8920 41810 9090
rect 41860 9230 41920 9250
rect 41860 9190 41870 9230
rect 41910 9190 41920 9230
rect 41860 9130 41920 9190
rect 41860 9090 41870 9130
rect 41910 9090 41920 9130
rect 41860 9030 41920 9090
rect 41970 9230 42030 9250
rect 41970 9190 41980 9230
rect 42020 9190 42030 9230
rect 41970 9130 42030 9190
rect 41970 9090 41980 9130
rect 42020 9090 42030 9130
rect 41850 9020 41930 9030
rect 41850 8960 41860 9020
rect 41920 8960 41930 9020
rect 41850 8950 41930 8960
rect 41970 8920 42030 9090
rect 42080 9230 42140 9250
rect 42080 9190 42090 9230
rect 42130 9190 42140 9230
rect 42080 9130 42140 9190
rect 42080 9090 42090 9130
rect 42130 9090 42140 9130
rect 42080 9030 42140 9090
rect 42190 9230 42250 9250
rect 42190 9190 42200 9230
rect 42240 9190 42250 9230
rect 42190 9130 42250 9190
rect 42190 9090 42200 9130
rect 42240 9090 42250 9130
rect 42070 9020 42150 9030
rect 42070 8960 42080 9020
rect 42140 8960 42150 9020
rect 42070 8950 42150 8960
rect 42190 8920 42250 9090
rect 42300 9230 42360 9250
rect 42300 9190 42310 9230
rect 42350 9190 42360 9230
rect 42300 9130 42360 9190
rect 42300 9090 42310 9130
rect 42350 9090 42360 9130
rect 42300 9030 42360 9090
rect 42410 9230 42470 9250
rect 42410 9190 42420 9230
rect 42460 9190 42470 9230
rect 42410 9130 42470 9190
rect 42410 9090 42420 9130
rect 42460 9090 42470 9130
rect 42290 9020 42370 9030
rect 42290 8960 42300 9020
rect 42360 8960 42370 9020
rect 42290 8950 42370 8960
rect 42410 8920 42470 9090
rect 42520 9230 42580 9250
rect 42520 9190 42530 9230
rect 42570 9190 42580 9230
rect 42520 9130 42580 9190
rect 42520 9090 42530 9130
rect 42570 9090 42580 9130
rect 42520 9030 42580 9090
rect 42630 9230 42690 9250
rect 42630 9190 42640 9230
rect 42680 9190 42690 9230
rect 42630 9130 42690 9190
rect 42630 9090 42640 9130
rect 42680 9090 42690 9130
rect 42510 9020 42590 9030
rect 42510 8960 42520 9020
rect 42580 8960 42590 9020
rect 42510 8950 42590 8960
rect 42630 8920 42690 9090
rect 42740 9230 42800 9250
rect 42740 9190 42750 9230
rect 42790 9190 42800 9230
rect 42740 9130 42800 9190
rect 42740 9090 42750 9130
rect 42790 9090 42800 9130
rect 42740 9030 42800 9090
rect 42850 9230 42910 9250
rect 42850 9190 42860 9230
rect 42900 9190 42910 9230
rect 42850 9130 42910 9190
rect 42850 9090 42860 9130
rect 42900 9090 42910 9130
rect 42730 9020 42810 9030
rect 42730 8960 42740 9020
rect 42800 8960 42810 9020
rect 42730 8950 42810 8960
rect 42850 8920 42910 9090
rect 42960 9230 43100 9250
rect 42960 9190 42970 9230
rect 43010 9190 43050 9230
rect 43090 9190 43100 9230
rect 42960 9130 43100 9190
rect 42960 9090 42970 9130
rect 43010 9090 43050 9130
rect 43090 9090 43100 9130
rect 42960 9070 43100 9090
rect 43460 9230 43600 9250
rect 43460 9190 43470 9230
rect 43510 9190 43550 9230
rect 43590 9190 43600 9230
rect 43460 9130 43600 9190
rect 43460 9090 43470 9130
rect 43510 9090 43550 9130
rect 43590 9090 43600 9130
rect 43460 9070 43600 9090
rect 42960 9030 43020 9070
rect 43540 9030 43600 9070
rect 43650 9230 43710 9250
rect 43650 9190 43660 9230
rect 43700 9190 43710 9230
rect 43650 9130 43710 9190
rect 43650 9090 43660 9130
rect 43700 9090 43710 9130
rect 42950 9020 43030 9030
rect 42950 8960 42960 9020
rect 43020 8960 43030 9020
rect 42950 8950 43030 8960
rect 43530 9020 43610 9030
rect 43530 8960 43540 9020
rect 43600 8960 43610 9020
rect 43530 8950 43610 8960
rect 39680 8850 39690 8910
rect 39750 8850 39760 8910
rect 39680 8840 39760 8850
rect 41740 8910 41820 8920
rect 41740 8850 41750 8910
rect 41810 8850 41820 8910
rect 41740 8840 41820 8850
rect 41960 8910 42040 8920
rect 41960 8850 41970 8910
rect 42030 8850 42040 8910
rect 41960 8840 42040 8850
rect 42180 8910 42260 8920
rect 42180 8850 42190 8910
rect 42250 8850 42260 8910
rect 42180 8840 42260 8850
rect 42400 8910 42480 8920
rect 42400 8850 42410 8910
rect 42470 8850 42480 8910
rect 42400 8840 42480 8850
rect 42620 8910 42700 8920
rect 42620 8850 42630 8910
rect 42690 8850 42700 8910
rect 42620 8840 42700 8850
rect 42840 8910 42920 8920
rect 43650 8910 43710 9090
rect 43760 9230 43820 9250
rect 43760 9190 43770 9230
rect 43810 9190 43820 9230
rect 43760 9130 43820 9190
rect 43760 9090 43770 9130
rect 43810 9090 43820 9130
rect 43760 9030 43820 9090
rect 43870 9230 43930 9250
rect 43870 9190 43880 9230
rect 43920 9190 43930 9230
rect 43870 9130 43930 9190
rect 43870 9090 43880 9130
rect 43920 9090 43930 9130
rect 43750 9020 43830 9030
rect 43750 8960 43760 9020
rect 43820 8960 43830 9020
rect 43750 8950 43830 8960
rect 43870 8910 43930 9090
rect 43980 9230 44040 9250
rect 43980 9190 43990 9230
rect 44030 9190 44040 9230
rect 43980 9130 44040 9190
rect 43980 9090 43990 9130
rect 44030 9090 44040 9130
rect 43980 9030 44040 9090
rect 44090 9230 44150 9250
rect 44090 9190 44100 9230
rect 44140 9190 44150 9230
rect 44090 9130 44150 9190
rect 44090 9090 44100 9130
rect 44140 9090 44150 9130
rect 43970 9020 44050 9030
rect 43970 8960 43980 9020
rect 44040 8960 44050 9020
rect 43970 8950 44050 8960
rect 44090 8910 44150 9090
rect 44200 9230 44260 9250
rect 44200 9190 44210 9230
rect 44250 9190 44260 9230
rect 44200 9130 44260 9190
rect 44200 9090 44210 9130
rect 44250 9090 44260 9130
rect 44200 9030 44260 9090
rect 44310 9230 44370 9250
rect 44310 9190 44320 9230
rect 44360 9190 44370 9230
rect 44310 9130 44370 9190
rect 44310 9090 44320 9130
rect 44360 9090 44370 9130
rect 44190 9020 44270 9030
rect 44190 8960 44200 9020
rect 44260 8960 44270 9020
rect 44190 8950 44270 8960
rect 44310 8910 44370 9090
rect 44420 9230 44480 9250
rect 44420 9190 44430 9230
rect 44470 9190 44480 9230
rect 44420 9130 44480 9190
rect 44420 9090 44430 9130
rect 44470 9090 44480 9130
rect 44420 9030 44480 9090
rect 44530 9230 44590 9250
rect 44530 9190 44540 9230
rect 44580 9190 44590 9230
rect 44530 9130 44590 9190
rect 44530 9090 44540 9130
rect 44580 9090 44590 9130
rect 44410 9020 44490 9030
rect 44410 8960 44420 9020
rect 44480 8960 44490 9020
rect 44410 8950 44490 8960
rect 44530 8910 44590 9090
rect 44640 9230 44700 9250
rect 44640 9190 44650 9230
rect 44690 9190 44700 9230
rect 44640 9130 44700 9190
rect 44640 9090 44650 9130
rect 44690 9090 44700 9130
rect 44640 9030 44700 9090
rect 44750 9230 44810 9250
rect 44750 9190 44760 9230
rect 44800 9190 44810 9230
rect 44750 9130 44810 9190
rect 44750 9090 44760 9130
rect 44800 9090 44810 9130
rect 44630 9020 44710 9030
rect 44630 8960 44640 9020
rect 44700 8960 44710 9020
rect 44630 8950 44710 8960
rect 44750 8910 44810 9090
rect 44860 9230 45000 9250
rect 44860 9190 44870 9230
rect 44910 9190 44950 9230
rect 44990 9190 45000 9230
rect 44860 9130 45000 9190
rect 44860 9090 44870 9130
rect 44910 9090 44950 9130
rect 44990 9090 45000 9130
rect 44860 9070 45000 9090
rect 44860 9030 44920 9070
rect 44850 9020 44930 9030
rect 44850 8960 44860 9020
rect 44920 8960 44930 9020
rect 44850 8950 44930 8960
rect 42840 8850 42850 8910
rect 42910 8850 42920 8910
rect 42840 8840 42920 8850
rect 43640 8900 43720 8910
rect 43640 8840 43650 8900
rect 43710 8840 43720 8900
rect 43640 8820 43720 8840
rect 43640 8760 43650 8820
rect 43710 8760 43720 8820
rect 43640 8740 43720 8760
rect 43640 8680 43650 8740
rect 43710 8680 43720 8740
rect 43640 8670 43720 8680
rect 43860 8900 43940 8910
rect 43860 8840 43870 8900
rect 43930 8840 43940 8900
rect 43860 8820 43940 8840
rect 43860 8760 43870 8820
rect 43930 8760 43940 8820
rect 43860 8740 43940 8760
rect 43860 8680 43870 8740
rect 43930 8680 43940 8740
rect 43860 8670 43940 8680
rect 44080 8900 44160 8910
rect 44080 8840 44090 8900
rect 44150 8840 44160 8900
rect 44080 8820 44160 8840
rect 44080 8760 44090 8820
rect 44150 8760 44160 8820
rect 44080 8740 44160 8760
rect 44080 8680 44090 8740
rect 44150 8680 44160 8740
rect 44080 8670 44160 8680
rect 44300 8900 44380 8910
rect 44300 8840 44310 8900
rect 44370 8840 44380 8900
rect 44300 8820 44380 8840
rect 44300 8760 44310 8820
rect 44370 8760 44380 8820
rect 44300 8740 44380 8760
rect 44300 8680 44310 8740
rect 44370 8680 44380 8740
rect 44300 8670 44380 8680
rect 44520 8900 44600 8910
rect 44520 8840 44530 8900
rect 44590 8840 44600 8900
rect 44520 8820 44600 8840
rect 44520 8760 44530 8820
rect 44590 8760 44600 8820
rect 44520 8740 44600 8760
rect 44520 8680 44530 8740
rect 44590 8680 44600 8740
rect 44520 8670 44600 8680
rect 44740 8900 44820 8910
rect 44740 8840 44750 8900
rect 44810 8840 44820 8900
rect 44740 8820 44820 8840
rect 44740 8760 44750 8820
rect 44810 8760 44820 8820
rect 44740 8740 44820 8760
rect 44740 8680 44750 8740
rect 44810 8680 44820 8740
rect 44740 8670 44820 8680
<< via1 >>
rect 39180 19130 39240 19190
rect 38800 19020 38860 19080
rect 38800 18940 38860 19000
rect 38800 18860 38860 18920
rect 38790 18050 38870 18420
rect 39180 18390 39240 18450
rect 39180 18310 39240 18370
rect 39180 18220 39240 18280
rect 39180 18130 39240 18190
rect 39180 18050 39240 18110
rect 39580 19020 39640 19080
rect 39580 18940 39640 19000
rect 39580 18860 39640 18920
rect 40690 19020 40750 19080
rect 40690 18940 40750 19000
rect 40690 18860 40750 18920
rect 38800 11120 38860 11180
rect 39470 13750 39530 13810
rect 40360 14660 40420 14720
rect 39580 12060 39640 12120
rect 39580 10740 39640 10800
rect 39690 14030 39750 14090
rect 39690 12290 39750 12350
rect 39470 10630 39530 10690
rect 38800 9300 38860 9360
rect 40630 13920 40690 13980
rect 48200 19130 48260 19190
rect 43250 19070 43310 19080
rect 43250 19030 43260 19070
rect 43260 19030 43300 19070
rect 43300 19030 43310 19070
rect 43250 19020 43310 19030
rect 43250 18990 43310 19000
rect 43250 18950 43260 18990
rect 43260 18950 43300 18990
rect 43300 18950 43310 18990
rect 43250 18940 43310 18950
rect 43250 18910 43310 18920
rect 43250 18870 43260 18910
rect 43260 18870 43300 18910
rect 43300 18870 43310 18910
rect 43250 18860 43310 18870
rect 45680 19020 45740 19080
rect 45680 18940 45740 19000
rect 45680 18860 45740 18920
rect 46790 19020 46850 19080
rect 46790 18940 46850 19000
rect 46790 18860 46850 18920
rect 47580 19020 47640 19080
rect 47580 18940 47640 19000
rect 47580 18860 47640 18920
rect 48200 18790 48260 18850
rect 47570 18050 47650 18420
rect 47960 18390 48020 18450
rect 47960 18310 48020 18370
rect 47960 18220 48020 18280
rect 47960 18130 48020 18190
rect 47960 18050 48020 18110
rect 48660 18090 48720 18150
rect 41150 16750 41210 16810
rect 41580 16750 41640 16810
rect 43250 16754 43310 16810
rect 43250 16750 43254 16754
rect 43254 16750 43310 16754
rect 45350 16750 45410 16810
rect 45350 14740 45410 14800
rect 47570 16680 47650 16760
rect 46360 15290 46420 15350
rect 46440 15290 46500 15350
rect 46520 15290 46580 15350
rect 46010 14740 46070 14800
rect 46250 14740 46310 14800
rect 44590 14660 44650 14720
rect 44680 14660 44740 14720
rect 44770 14660 44830 14720
rect 44860 14660 44920 14720
rect 44950 14660 45010 14720
rect 41150 14350 41210 14410
rect 41560 14350 41960 14402
rect 44600 14398 45000 14402
rect 44600 14360 44996 14398
rect 44996 14360 45000 14398
rect 44600 14350 45000 14360
rect 46160 14350 46220 14410
rect 41040 13920 41100 13980
rect 41090 13800 41150 13810
rect 41090 13760 41100 13800
rect 41100 13760 41140 13800
rect 41140 13760 41150 13800
rect 41090 13750 41150 13760
rect 45480 13840 45540 13850
rect 45480 13800 45490 13840
rect 45490 13800 45530 13840
rect 45530 13800 45540 13840
rect 45480 13790 45540 13800
rect 45480 13760 45540 13770
rect 45480 13720 45490 13760
rect 45490 13720 45530 13760
rect 45530 13720 45540 13760
rect 45480 13710 45540 13720
rect 41170 13630 41230 13640
rect 41170 13590 41180 13630
rect 41180 13590 41220 13630
rect 41220 13590 41230 13630
rect 41170 13580 41230 13590
rect 41330 13630 41390 13640
rect 41330 13590 41340 13630
rect 41340 13590 41380 13630
rect 41380 13590 41390 13630
rect 41330 13580 41390 13590
rect 41490 13630 41550 13640
rect 41490 13590 41500 13630
rect 41500 13590 41540 13630
rect 41540 13590 41550 13630
rect 41490 13580 41550 13590
rect 41650 13630 41710 13640
rect 41650 13590 41660 13630
rect 41660 13590 41700 13630
rect 41700 13590 41710 13630
rect 41650 13580 41710 13590
rect 41810 13630 41870 13640
rect 41810 13590 41820 13630
rect 41820 13590 41860 13630
rect 41860 13590 41870 13630
rect 41810 13580 41870 13590
rect 41970 13630 42030 13640
rect 41970 13590 41980 13630
rect 41980 13590 42020 13630
rect 42020 13590 42030 13630
rect 41970 13580 42030 13590
rect 42130 13630 42190 13640
rect 42130 13590 42140 13630
rect 42140 13590 42180 13630
rect 42180 13590 42190 13630
rect 42130 13580 42190 13590
rect 42290 13630 42350 13640
rect 42290 13590 42300 13630
rect 42300 13590 42340 13630
rect 42340 13590 42350 13630
rect 42290 13580 42350 13590
rect 42450 13630 42510 13640
rect 42450 13590 42460 13630
rect 42460 13590 42500 13630
rect 42500 13590 42510 13630
rect 42450 13580 42510 13590
rect 42610 13630 42670 13640
rect 42610 13590 42620 13630
rect 42620 13590 42660 13630
rect 42660 13590 42670 13630
rect 42610 13580 42670 13590
rect 42770 13630 42830 13640
rect 42770 13590 42780 13630
rect 42780 13590 42820 13630
rect 42820 13590 42830 13630
rect 42770 13580 42830 13590
rect 42930 13630 42990 13640
rect 42930 13590 42940 13630
rect 42940 13590 42980 13630
rect 42980 13590 42990 13630
rect 42930 13580 42990 13590
rect 43090 13630 43150 13640
rect 43090 13590 43100 13630
rect 43100 13590 43140 13630
rect 43140 13590 43150 13630
rect 43090 13580 43150 13590
rect 43250 13630 43310 13640
rect 43250 13590 43260 13630
rect 43260 13590 43300 13630
rect 43300 13590 43310 13630
rect 43250 13580 43310 13590
rect 43410 13630 43470 13640
rect 43410 13590 43420 13630
rect 43420 13590 43460 13630
rect 43460 13590 43470 13630
rect 43410 13580 43470 13590
rect 43570 13630 43630 13640
rect 43570 13590 43580 13630
rect 43580 13590 43620 13630
rect 43620 13590 43630 13630
rect 43570 13580 43630 13590
rect 43730 13630 43790 13640
rect 43730 13590 43740 13630
rect 43740 13590 43780 13630
rect 43780 13590 43790 13630
rect 43730 13580 43790 13590
rect 43890 13630 43950 13640
rect 43890 13590 43900 13630
rect 43900 13590 43940 13630
rect 43940 13590 43950 13630
rect 43890 13580 43950 13590
rect 44050 13630 44110 13640
rect 44050 13590 44060 13630
rect 44060 13590 44100 13630
rect 44100 13590 44110 13630
rect 44050 13580 44110 13590
rect 44210 13630 44270 13640
rect 44210 13590 44220 13630
rect 44220 13590 44260 13630
rect 44260 13590 44270 13630
rect 44210 13580 44270 13590
rect 44370 13630 44430 13640
rect 44370 13590 44380 13630
rect 44380 13590 44420 13630
rect 44420 13590 44430 13630
rect 44370 13580 44430 13590
rect 44530 13630 44590 13640
rect 44530 13590 44540 13630
rect 44540 13590 44580 13630
rect 44580 13590 44590 13630
rect 44530 13580 44590 13590
rect 44690 13630 44750 13640
rect 44690 13590 44700 13630
rect 44700 13590 44740 13630
rect 44740 13590 44750 13630
rect 44690 13580 44750 13590
rect 44850 13630 44910 13640
rect 44850 13590 44860 13630
rect 44860 13590 44900 13630
rect 44900 13590 44910 13630
rect 44850 13580 44910 13590
rect 45010 13630 45070 13640
rect 45010 13590 45020 13630
rect 45020 13590 45060 13630
rect 45060 13590 45070 13630
rect 45010 13580 45070 13590
rect 45170 13630 45230 13640
rect 45170 13590 45180 13630
rect 45180 13590 45220 13630
rect 45220 13590 45230 13630
rect 45170 13580 45230 13590
rect 41910 13470 41970 13530
rect 41910 13390 41970 13450
rect 41910 13360 41970 13370
rect 41910 13320 41920 13360
rect 41920 13320 41960 13360
rect 41960 13320 41970 13360
rect 41910 13310 41970 13320
rect 43170 13470 43230 13530
rect 43250 13470 43310 13530
rect 43330 13470 43390 13530
rect 43170 13390 43230 13450
rect 43250 13390 43310 13450
rect 43330 13390 43390 13450
rect 43170 13310 43230 13370
rect 43250 13310 43310 13370
rect 43330 13310 43390 13370
rect 40930 12720 40990 12730
rect 40930 12680 40940 12720
rect 40940 12680 40980 12720
rect 40980 12680 40990 12720
rect 40930 12670 40990 12680
rect 40930 12590 40990 12650
rect 40930 12510 40990 12570
rect 41170 12720 41230 12730
rect 41170 12680 41180 12720
rect 41180 12680 41220 12720
rect 41220 12680 41230 12720
rect 41170 12670 41230 12680
rect 41170 12590 41230 12650
rect 41170 12510 41230 12570
rect 41410 12720 41470 12730
rect 41410 12680 41420 12720
rect 41420 12680 41460 12720
rect 41460 12680 41470 12720
rect 41410 12670 41470 12680
rect 41410 12590 41470 12650
rect 41410 12510 41470 12570
rect 41650 12720 41710 12730
rect 41650 12680 41660 12720
rect 41660 12680 41700 12720
rect 41700 12680 41710 12720
rect 41650 12670 41710 12680
rect 41650 12590 41710 12650
rect 41650 12510 41710 12570
rect 42290 12720 42350 12730
rect 42290 12680 42300 12720
rect 42300 12680 42340 12720
rect 42340 12680 42350 12720
rect 42290 12670 42350 12680
rect 42290 12590 42350 12650
rect 42290 12510 42350 12570
rect 42530 12720 42590 12730
rect 42530 12680 42540 12720
rect 42540 12680 42580 12720
rect 42580 12680 42590 12720
rect 42530 12670 42590 12680
rect 42530 12590 42590 12650
rect 42530 12510 42590 12570
rect 42770 12720 42830 12730
rect 42770 12680 42780 12720
rect 42780 12680 42820 12720
rect 42820 12680 42830 12720
rect 42770 12670 42830 12680
rect 42770 12590 42830 12650
rect 42770 12510 42830 12570
rect 40750 12400 40810 12460
rect 41500 12400 41560 12460
rect 41720 12400 41780 12460
rect 41980 12400 42040 12460
rect 42200 12400 42260 12460
rect 42460 12400 42520 12460
rect 41433 12342 41485 12350
rect 41433 12308 41443 12342
rect 41443 12308 41477 12342
rect 41477 12308 41485 12342
rect 41433 12298 41485 12308
rect 41793 12342 41845 12350
rect 41793 12308 41803 12342
rect 41803 12308 41837 12342
rect 41837 12308 41845 12342
rect 41793 12298 41845 12308
rect 41913 12342 41965 12350
rect 41913 12308 41923 12342
rect 41923 12308 41957 12342
rect 41957 12308 41965 12342
rect 41913 12298 41965 12308
rect 42273 12342 42325 12350
rect 42273 12308 42283 12342
rect 42283 12308 42317 12342
rect 42317 12308 42325 12342
rect 42273 12298 42325 12308
rect 42393 12342 42445 12350
rect 42393 12308 42403 12342
rect 42403 12308 42437 12342
rect 42437 12308 42445 12342
rect 42393 12298 42445 12308
rect 42810 12320 42870 12330
rect 42810 12280 42820 12320
rect 42820 12280 42860 12320
rect 42860 12280 42870 12320
rect 42810 12270 42870 12280
rect 42810 12240 42870 12250
rect 42810 12200 42820 12240
rect 42820 12200 42860 12240
rect 42860 12200 42870 12240
rect 42810 12190 42870 12200
rect 41536 12112 41588 12122
rect 41536 12078 41544 12112
rect 41544 12078 41578 12112
rect 41578 12078 41588 12112
rect 41536 12070 41588 12078
rect 41694 12112 41746 12122
rect 41694 12078 41702 12112
rect 41702 12078 41736 12112
rect 41736 12078 41746 12112
rect 41694 12070 41746 12078
rect 41610 11960 41670 12020
rect 41370 11850 41430 11910
rect 40630 11580 40690 11640
rect 40710 11580 40770 11640
rect 41130 11580 41190 11640
rect 41370 11580 41430 11640
rect 40890 11510 40950 11520
rect 40890 11470 40900 11510
rect 40900 11470 40940 11510
rect 40940 11470 40950 11510
rect 40890 11460 40950 11470
rect 40650 11120 40710 11180
rect 42018 12112 42070 12122
rect 42018 12078 42026 12112
rect 42026 12078 42060 12112
rect 42060 12078 42070 12112
rect 42018 12070 42070 12078
rect 42172 12112 42224 12122
rect 42172 12078 42180 12112
rect 42180 12078 42214 12112
rect 42214 12078 42224 12112
rect 42172 12070 42224 12078
rect 42090 11960 42150 12020
rect 42496 12112 42548 12122
rect 42496 12078 42504 12112
rect 42504 12078 42538 12112
rect 42538 12078 42548 12112
rect 42496 12070 42548 12078
rect 42810 12160 42870 12170
rect 42810 12120 42820 12160
rect 42820 12120 42860 12160
rect 42860 12120 42870 12160
rect 42810 12110 42870 12120
rect 42570 11960 42630 12020
rect 41850 11850 41910 11910
rect 42330 11850 42390 11910
rect 41850 11580 41910 11640
rect 42090 11580 42150 11640
rect 42570 11580 42630 11640
rect 42750 11580 42810 11640
rect 41610 11510 41670 11520
rect 41610 11470 41620 11510
rect 41620 11470 41660 11510
rect 41660 11470 41670 11510
rect 41610 11460 41670 11470
rect 41370 11120 41430 11180
rect 42330 11510 42390 11520
rect 42330 11470 42340 11510
rect 42340 11470 42380 11510
rect 42380 11470 42390 11510
rect 42330 11460 42390 11470
rect 42090 11120 42150 11180
rect 42810 11120 42870 11180
rect 44590 13470 44650 13530
rect 44590 13390 44650 13450
rect 44590 13360 44650 13370
rect 44590 13320 44600 13360
rect 44600 13320 44640 13360
rect 44640 13320 44650 13360
rect 44590 13310 44650 13320
rect 43170 12270 43230 12330
rect 43250 12270 43310 12330
rect 43330 12270 43390 12330
rect 43170 12190 43230 12250
rect 43250 12190 43310 12250
rect 43330 12190 43390 12250
rect 43170 12110 43230 12170
rect 43250 12110 43310 12170
rect 43330 12110 43390 12170
rect 43730 12720 43790 12730
rect 43730 12680 43740 12720
rect 43740 12680 43780 12720
rect 43780 12680 43790 12720
rect 43730 12670 43790 12680
rect 43730 12590 43790 12650
rect 43730 12510 43790 12570
rect 43970 12720 44030 12730
rect 43970 12680 43980 12720
rect 43980 12680 44020 12720
rect 44020 12680 44030 12720
rect 43970 12670 44030 12680
rect 43970 12590 44030 12650
rect 43970 12510 44030 12570
rect 44210 12720 44270 12730
rect 44210 12680 44220 12720
rect 44220 12680 44260 12720
rect 44260 12680 44270 12720
rect 44210 12670 44270 12680
rect 44210 12590 44270 12650
rect 44210 12510 44270 12570
rect 44850 12720 44910 12730
rect 44850 12680 44860 12720
rect 44860 12680 44900 12720
rect 44900 12680 44910 12720
rect 44850 12670 44910 12680
rect 44850 12590 44910 12650
rect 44850 12510 44910 12570
rect 45090 12720 45150 12730
rect 45090 12680 45100 12720
rect 45100 12680 45140 12720
rect 45140 12680 45150 12720
rect 45090 12670 45150 12680
rect 45090 12590 45150 12650
rect 45090 12510 45150 12570
rect 45330 12720 45390 12730
rect 45330 12680 45340 12720
rect 45340 12680 45380 12720
rect 45380 12680 45390 12720
rect 45330 12670 45390 12680
rect 45330 12590 45390 12650
rect 45330 12510 45390 12570
rect 45570 12720 45630 12730
rect 45570 12680 45580 12720
rect 45580 12680 45620 12720
rect 45620 12680 45630 12720
rect 45570 12670 45630 12680
rect 45570 12590 45630 12650
rect 45570 12510 45630 12570
rect 44040 12400 44100 12460
rect 44300 12400 44360 12460
rect 44520 12400 44580 12460
rect 44780 12400 44840 12460
rect 45000 12400 45060 12460
rect 45750 12400 45810 12460
rect 43690 12320 43750 12330
rect 43690 12280 43700 12320
rect 43700 12280 43740 12320
rect 43740 12280 43750 12320
rect 43690 12270 43750 12280
rect 44115 12342 44167 12350
rect 44115 12308 44123 12342
rect 44123 12308 44157 12342
rect 44157 12308 44167 12342
rect 44115 12298 44167 12308
rect 44235 12342 44287 12350
rect 44235 12308 44243 12342
rect 44243 12308 44277 12342
rect 44277 12308 44287 12342
rect 44235 12298 44287 12308
rect 44595 12342 44647 12350
rect 44595 12308 44603 12342
rect 44603 12308 44637 12342
rect 44637 12308 44647 12342
rect 44595 12298 44647 12308
rect 44715 12342 44767 12350
rect 44715 12308 44723 12342
rect 44723 12308 44757 12342
rect 44757 12308 44767 12342
rect 44715 12298 44767 12308
rect 45075 12342 45127 12350
rect 45075 12308 45083 12342
rect 45083 12308 45117 12342
rect 45117 12308 45127 12342
rect 45075 12298 45127 12308
rect 46160 12290 46220 12350
rect 43690 12240 43750 12250
rect 43690 12200 43700 12240
rect 43700 12200 43740 12240
rect 43740 12200 43750 12240
rect 43690 12190 43750 12200
rect 43690 12160 43750 12170
rect 43690 12120 43700 12160
rect 43700 12120 43740 12160
rect 43740 12120 43750 12160
rect 43690 12110 43750 12120
rect 44012 12112 44064 12122
rect 44012 12078 44022 12112
rect 44022 12078 44056 12112
rect 44056 12078 44064 12112
rect 44012 12070 44064 12078
rect 43930 11960 43990 12020
rect 44336 12112 44388 12122
rect 44336 12078 44346 12112
rect 44346 12078 44380 12112
rect 44380 12078 44388 12112
rect 44336 12070 44388 12078
rect 44490 12112 44542 12122
rect 44490 12078 44500 12112
rect 44500 12078 44534 12112
rect 44534 12078 44542 12112
rect 44490 12070 44542 12078
rect 44410 11960 44470 12020
rect 44814 12112 44866 12122
rect 44814 12078 44824 12112
rect 44824 12078 44858 12112
rect 44858 12078 44866 12112
rect 44814 12070 44866 12078
rect 44972 12112 45024 12122
rect 44972 12078 44982 12112
rect 44982 12078 45016 12112
rect 45016 12078 45024 12112
rect 44972 12070 45024 12078
rect 44890 11960 44950 12020
rect 44170 11850 44230 11910
rect 44650 11850 44710 11910
rect 43750 11740 43810 11800
rect 43750 11660 43810 11720
rect 43750 11580 43810 11640
rect 43930 11740 43990 11800
rect 43930 11660 43990 11720
rect 43930 11580 43990 11640
rect 44170 11740 44230 11800
rect 44170 11660 44230 11720
rect 44170 11580 44230 11640
rect 44410 11740 44470 11800
rect 44410 11660 44470 11720
rect 44410 11580 44470 11640
rect 44650 11740 44710 11800
rect 44650 11660 44710 11720
rect 44650 11580 44710 11640
rect 43070 11120 43130 11180
rect 43430 11120 43490 11180
rect 40530 11010 40590 11070
rect 40530 10930 40590 10990
rect 40530 10850 40590 10910
rect 40770 11010 40830 11070
rect 40770 10930 40830 10990
rect 40770 10850 40830 10910
rect 41010 11010 41070 11070
rect 41010 10930 41070 10990
rect 41010 10850 41070 10910
rect 41250 11010 41310 11070
rect 41250 10930 41310 10990
rect 41250 10850 41310 10910
rect 41490 11010 41550 11070
rect 41490 10930 41550 10990
rect 41490 10850 41550 10910
rect 41730 11010 41790 11070
rect 41730 10930 41790 10990
rect 41730 10850 41790 10910
rect 41970 11010 42030 11070
rect 41970 10930 42030 10990
rect 41970 10850 42030 10910
rect 42210 11010 42270 11070
rect 42210 10930 42270 10990
rect 42210 10850 42270 10910
rect 42450 11010 42510 11070
rect 42450 10930 42510 10990
rect 42450 10850 42510 10910
rect 42690 11010 42750 11070
rect 42690 10930 42750 10990
rect 42690 10850 42750 10910
rect 42930 11010 42990 11070
rect 42930 10930 42990 10990
rect 42930 10850 42990 10910
rect 41810 10740 41870 10800
rect 43250 10740 43310 10800
rect 42170 10630 42230 10690
rect 41900 10350 41960 10360
rect 41900 10310 41910 10350
rect 41910 10310 41950 10350
rect 41950 10310 41960 10350
rect 41900 10300 41960 10310
rect 42080 10350 42140 10360
rect 42080 10310 42090 10350
rect 42090 10310 42130 10350
rect 42130 10310 42140 10350
rect 42080 10300 42140 10310
rect 42530 10520 42590 10580
rect 42260 10350 42320 10360
rect 42260 10310 42270 10350
rect 42270 10310 42310 10350
rect 42310 10310 42320 10350
rect 42260 10300 42320 10310
rect 42440 10350 42500 10360
rect 42440 10310 42450 10350
rect 42450 10310 42490 10350
rect 42490 10310 42500 10350
rect 42440 10300 42500 10310
rect 42890 10410 42950 10470
rect 42620 10350 42680 10360
rect 42620 10310 42630 10350
rect 42630 10310 42670 10350
rect 42670 10310 42680 10350
rect 42620 10300 42680 10310
rect 42800 10350 42860 10360
rect 42800 10310 42810 10350
rect 42810 10310 42850 10350
rect 42850 10310 42860 10350
rect 42800 10300 42860 10310
rect 42980 10350 43040 10360
rect 42980 10310 42990 10350
rect 42990 10310 43030 10350
rect 43030 10310 43040 10350
rect 42980 10300 43040 10310
rect 43160 10350 43220 10360
rect 43160 10310 43170 10350
rect 43170 10310 43210 10350
rect 43210 10310 43220 10350
rect 43160 10300 43220 10310
rect 43690 11120 43750 11180
rect 44170 11510 44230 11520
rect 44170 11470 44180 11510
rect 44180 11470 44220 11510
rect 44220 11470 44230 11510
rect 44170 11460 44230 11470
rect 44410 11120 44470 11180
rect 45130 11850 45190 11910
rect 45130 11740 45190 11800
rect 45130 11660 45190 11720
rect 45130 11580 45190 11640
rect 45370 11740 45430 11800
rect 45370 11660 45430 11720
rect 45370 11580 45430 11640
rect 45790 11740 45850 11800
rect 45790 11660 45850 11720
rect 45790 11580 45850 11640
rect 44890 11510 44950 11520
rect 44890 11470 44900 11510
rect 44900 11470 44940 11510
rect 44940 11470 44950 11510
rect 44890 11460 44950 11470
rect 45130 11120 45190 11180
rect 45610 11510 45670 11520
rect 45610 11470 45620 11510
rect 45620 11470 45660 11510
rect 45660 11470 45670 11510
rect 45610 11460 45670 11470
rect 45850 11120 45910 11180
rect 43570 11010 43630 11070
rect 43570 10930 43630 10990
rect 43570 10850 43630 10910
rect 43810 11010 43870 11070
rect 43810 10930 43870 10990
rect 43810 10850 43870 10910
rect 44050 11010 44110 11070
rect 44050 10930 44110 10990
rect 44050 10850 44110 10910
rect 44290 11010 44350 11070
rect 44290 10930 44350 10990
rect 44290 10850 44350 10910
rect 44530 11010 44590 11070
rect 44530 10930 44590 10990
rect 44530 10850 44590 10910
rect 44770 11010 44830 11070
rect 44770 10930 44830 10990
rect 44770 10850 44830 10910
rect 45010 11010 45070 11070
rect 45010 10930 45070 10990
rect 45010 10850 45070 10910
rect 45250 11010 45310 11070
rect 45250 10930 45310 10990
rect 45250 10850 45310 10910
rect 45490 11010 45550 11070
rect 45490 10930 45550 10990
rect 45490 10850 45550 10910
rect 45730 11010 45790 11070
rect 45730 10930 45790 10990
rect 45730 10850 45790 10910
rect 44690 10740 44750 10800
rect 44330 10630 44390 10690
rect 43970 10520 44030 10580
rect 43610 10410 43670 10470
rect 43340 10350 43400 10360
rect 43340 10310 43350 10350
rect 43350 10310 43390 10350
rect 43390 10310 43400 10350
rect 43340 10300 43400 10310
rect 43430 10300 43490 10360
rect 43520 10350 43580 10360
rect 43520 10310 43530 10350
rect 43530 10310 43570 10350
rect 43570 10310 43580 10350
rect 43520 10300 43580 10310
rect 43700 10350 43760 10360
rect 43700 10310 43710 10350
rect 43710 10310 43750 10350
rect 43750 10310 43760 10350
rect 43700 10300 43760 10310
rect 43880 10350 43940 10360
rect 43880 10310 43890 10350
rect 43890 10310 43930 10350
rect 43930 10310 43940 10350
rect 43880 10300 43940 10310
rect 44060 10350 44120 10360
rect 44060 10310 44070 10350
rect 44070 10310 44110 10350
rect 44110 10310 44120 10350
rect 44060 10300 44120 10310
rect 44240 10350 44300 10360
rect 44240 10310 44250 10350
rect 44250 10310 44290 10350
rect 44290 10310 44300 10350
rect 44240 10300 44300 10310
rect 44420 10350 44480 10360
rect 44420 10310 44430 10350
rect 44430 10310 44470 10350
rect 44470 10310 44480 10350
rect 44420 10300 44480 10310
rect 44600 10350 44660 10360
rect 44600 10310 44610 10350
rect 44610 10310 44650 10350
rect 44650 10310 44660 10350
rect 44600 10300 44660 10310
rect 45720 10630 45780 10690
rect 45250 10520 45310 10580
rect 45600 10150 45660 10160
rect 45600 10110 45610 10150
rect 45610 10110 45650 10150
rect 45650 10110 45660 10150
rect 45600 10100 45660 10110
rect 45970 11010 46030 11070
rect 45970 10930 46030 10990
rect 45970 10850 46030 10910
rect 46250 12060 46310 12120
rect 46790 14030 46850 14090
rect 46360 11740 46420 11800
rect 46440 11740 46500 11800
rect 46520 11740 46580 11800
rect 46360 11660 46420 11720
rect 46440 11660 46500 11720
rect 46520 11660 46580 11720
rect 46360 11580 46420 11640
rect 46440 11580 46500 11640
rect 46520 11580 46580 11640
rect 47960 15990 48020 16050
rect 48130 17390 48190 17450
rect 48800 16690 48860 16750
rect 48800 15290 48860 15350
rect 48660 13920 48720 13980
rect 47580 11120 47640 11180
rect 46250 10520 46310 10580
rect 46160 10410 46220 10470
rect 45840 10150 45900 10160
rect 45840 10110 45850 10150
rect 45850 10110 45890 10150
rect 45890 10110 45900 10150
rect 45840 10100 45900 10110
rect 45250 9760 45310 9820
rect 45720 9810 45780 9820
rect 45720 9770 45730 9810
rect 45730 9770 45770 9810
rect 45770 9770 45780 9810
rect 45720 9760 45780 9770
rect 41630 9610 41690 9620
rect 41630 9570 41640 9610
rect 41640 9570 41680 9610
rect 41680 9570 41690 9610
rect 41630 9560 41690 9570
rect 41630 9480 41690 9540
rect 41630 9400 41690 9460
rect 41990 9610 42050 9620
rect 41990 9570 42000 9610
rect 42000 9570 42040 9610
rect 42040 9570 42050 9610
rect 41990 9560 42050 9570
rect 41990 9480 42050 9540
rect 41990 9400 42050 9460
rect 42350 9610 42410 9620
rect 42350 9570 42360 9610
rect 42360 9570 42400 9610
rect 42400 9570 42410 9610
rect 42350 9560 42410 9570
rect 42350 9480 42410 9540
rect 42350 9400 42410 9460
rect 42710 9610 42770 9620
rect 42710 9570 42720 9610
rect 42720 9570 42760 9610
rect 42760 9570 42770 9610
rect 42710 9560 42770 9570
rect 42710 9480 42770 9540
rect 42710 9400 42770 9460
rect 43070 9610 43130 9620
rect 43070 9570 43080 9610
rect 43080 9570 43120 9610
rect 43120 9570 43130 9610
rect 43070 9560 43130 9570
rect 43070 9480 43130 9540
rect 43070 9400 43130 9460
rect 43430 9610 43490 9620
rect 43430 9570 43440 9610
rect 43440 9570 43480 9610
rect 43480 9570 43490 9610
rect 43430 9560 43490 9570
rect 43430 9480 43490 9540
rect 43430 9400 43490 9460
rect 43790 9610 43850 9620
rect 43790 9570 43800 9610
rect 43800 9570 43840 9610
rect 43840 9570 43850 9610
rect 43790 9560 43850 9570
rect 43790 9480 43850 9540
rect 43790 9400 43850 9460
rect 44150 9610 44210 9620
rect 44150 9570 44160 9610
rect 44160 9570 44200 9610
rect 44200 9570 44210 9610
rect 44150 9560 44210 9570
rect 44150 9480 44210 9540
rect 44150 9400 44210 9460
rect 44510 9610 44570 9620
rect 44510 9570 44520 9610
rect 44520 9570 44560 9610
rect 44560 9570 44570 9610
rect 44510 9560 44570 9570
rect 44510 9480 44570 9540
rect 44510 9400 44570 9460
rect 44870 9610 44930 9620
rect 44870 9570 44880 9610
rect 44880 9570 44920 9610
rect 44920 9570 44930 9610
rect 44870 9560 44930 9570
rect 44870 9480 44930 9540
rect 44870 9400 44930 9460
rect 45500 9560 45560 9620
rect 45500 9480 45560 9540
rect 45500 9400 45560 9460
rect 45940 9560 46000 9620
rect 45940 9480 46000 9540
rect 45940 9400 46000 9460
rect 41808 9342 41860 9350
rect 41808 9308 41818 9342
rect 41818 9308 41852 9342
rect 41852 9308 41860 9342
rect 41808 9298 41860 9308
rect 41918 9342 41970 9350
rect 41918 9308 41928 9342
rect 41928 9308 41962 9342
rect 41962 9308 41970 9342
rect 41918 9298 41970 9308
rect 42028 9342 42080 9350
rect 42028 9308 42038 9342
rect 42038 9308 42072 9342
rect 42072 9308 42080 9342
rect 42028 9298 42080 9308
rect 42138 9342 42190 9350
rect 42138 9308 42148 9342
rect 42148 9308 42182 9342
rect 42182 9308 42190 9342
rect 42138 9298 42190 9308
rect 42248 9342 42300 9350
rect 42248 9308 42258 9342
rect 42258 9308 42292 9342
rect 42292 9308 42300 9342
rect 42248 9298 42300 9308
rect 42358 9342 42410 9350
rect 42358 9308 42368 9342
rect 42368 9308 42402 9342
rect 42402 9308 42410 9342
rect 42358 9298 42410 9308
rect 42468 9342 42520 9350
rect 42468 9308 42478 9342
rect 42478 9308 42512 9342
rect 42512 9308 42520 9342
rect 42468 9298 42520 9308
rect 42578 9342 42630 9350
rect 42578 9308 42588 9342
rect 42588 9308 42622 9342
rect 42622 9308 42630 9342
rect 42578 9298 42630 9308
rect 42688 9342 42740 9350
rect 42688 9308 42698 9342
rect 42698 9308 42732 9342
rect 42732 9308 42740 9342
rect 42688 9298 42740 9308
rect 42798 9342 42850 9350
rect 42798 9308 42808 9342
rect 42808 9308 42842 9342
rect 42842 9308 42850 9342
rect 42798 9298 42850 9308
rect 43708 9342 43760 9350
rect 43708 9308 43718 9342
rect 43718 9308 43752 9342
rect 43752 9308 43760 9342
rect 43708 9298 43760 9308
rect 43818 9342 43870 9350
rect 43818 9308 43828 9342
rect 43828 9308 43862 9342
rect 43862 9308 43870 9342
rect 43818 9298 43870 9308
rect 43928 9342 43980 9350
rect 43928 9308 43938 9342
rect 43938 9308 43972 9342
rect 43972 9308 43980 9342
rect 43928 9298 43980 9308
rect 44038 9342 44090 9350
rect 44038 9308 44048 9342
rect 44048 9308 44082 9342
rect 44082 9308 44090 9342
rect 44038 9298 44090 9308
rect 44148 9342 44200 9350
rect 44148 9308 44158 9342
rect 44158 9308 44192 9342
rect 44192 9308 44200 9342
rect 44148 9298 44200 9308
rect 44258 9342 44310 9350
rect 44258 9308 44268 9342
rect 44268 9308 44302 9342
rect 44302 9308 44310 9342
rect 44258 9298 44310 9308
rect 44368 9342 44420 9350
rect 44368 9308 44378 9342
rect 44378 9308 44412 9342
rect 44412 9308 44420 9342
rect 44368 9298 44420 9308
rect 44478 9342 44530 9350
rect 44478 9308 44488 9342
rect 44488 9308 44522 9342
rect 44522 9308 44530 9342
rect 44478 9298 44530 9308
rect 44588 9342 44640 9350
rect 44588 9308 44598 9342
rect 44598 9308 44632 9342
rect 44632 9308 44640 9342
rect 44588 9298 44640 9308
rect 44698 9342 44750 9350
rect 44698 9308 44708 9342
rect 44708 9308 44742 9342
rect 44742 9308 44750 9342
rect 44698 9298 44750 9308
rect 41640 9010 41700 9020
rect 41640 8970 41650 9010
rect 41650 8970 41690 9010
rect 41690 8970 41700 9010
rect 41640 8960 41700 8970
rect 41860 8960 41920 9020
rect 42080 8960 42140 9020
rect 42300 8960 42360 9020
rect 42520 8960 42580 9020
rect 42740 8960 42800 9020
rect 42960 9010 43020 9020
rect 42960 8970 42970 9010
rect 42970 8970 43010 9010
rect 43010 8970 43020 9010
rect 42960 8960 43020 8970
rect 43540 9010 43600 9020
rect 43540 8970 43550 9010
rect 43550 8970 43590 9010
rect 43590 8970 43600 9010
rect 43540 8960 43600 8970
rect 39690 8850 39750 8910
rect 41750 8850 41810 8910
rect 41970 8850 42030 8910
rect 42190 8850 42250 8910
rect 42410 8850 42470 8910
rect 42630 8850 42690 8910
rect 43760 8960 43820 9020
rect 43980 8960 44040 9020
rect 44200 8960 44260 9020
rect 44420 8960 44480 9020
rect 44640 8960 44700 9020
rect 44860 9010 44920 9020
rect 44860 8970 44870 9010
rect 44870 8970 44910 9010
rect 44910 8970 44920 9010
rect 44860 8960 44920 8970
rect 42850 8850 42910 8910
rect 43650 8840 43710 8900
rect 43650 8760 43710 8820
rect 43650 8680 43710 8740
rect 43870 8840 43930 8900
rect 43870 8760 43930 8820
rect 43870 8680 43930 8740
rect 44090 8840 44150 8900
rect 44090 8760 44150 8820
rect 44090 8680 44150 8740
rect 44310 8840 44370 8900
rect 44310 8760 44370 8820
rect 44310 8680 44370 8740
rect 44530 8840 44590 8900
rect 44530 8760 44590 8820
rect 44530 8680 44590 8740
rect 44750 8840 44810 8900
rect 44750 8760 44810 8820
rect 44750 8680 44810 8740
<< metal2 >>
rect 39170 19190 48270 19200
rect 39170 19130 39180 19190
rect 39240 19130 48200 19190
rect 48260 19130 48270 19190
rect 39170 19120 48270 19130
rect 38790 19080 47650 19090
rect 38790 19020 38800 19080
rect 38860 19020 39580 19080
rect 39640 19020 40690 19080
rect 40750 19020 43250 19080
rect 43310 19020 45680 19080
rect 45740 19020 46790 19080
rect 46850 19020 47580 19080
rect 47640 19020 47650 19080
rect 38790 19000 47650 19020
rect 38790 18940 38800 19000
rect 38860 18940 39580 19000
rect 39640 18940 40690 19000
rect 40750 18940 43250 19000
rect 43310 18940 45680 19000
rect 45740 18940 46790 19000
rect 46850 18940 47580 19000
rect 47640 18940 47650 19000
rect 38790 18920 47650 18940
rect 38790 18860 38800 18920
rect 38860 18860 39580 18920
rect 39640 18860 40690 18920
rect 40750 18860 43250 18920
rect 43310 18860 45680 18920
rect 45740 18860 46790 18920
rect 46850 18860 47580 18920
rect 47640 18860 47650 18920
rect 38790 18850 47650 18860
rect 48190 18850 48270 18860
rect 48190 18790 48200 18850
rect 48260 18790 48270 18850
rect 48190 18780 48270 18790
rect 38770 18450 39250 18460
rect 38770 18420 39180 18450
rect 38770 18050 38790 18420
rect 38870 18390 39180 18420
rect 39240 18390 39250 18450
rect 38870 18370 39250 18390
rect 38870 18310 39180 18370
rect 39240 18310 39250 18370
rect 38870 18280 39250 18310
rect 38870 18220 39180 18280
rect 39240 18220 39250 18280
rect 38870 18190 39250 18220
rect 38870 18130 39180 18190
rect 39240 18130 39250 18190
rect 38870 18110 39250 18130
rect 38870 18050 39180 18110
rect 39240 18050 39250 18110
rect 38770 18030 39250 18050
rect 47550 18450 48030 18460
rect 47550 18420 47960 18450
rect 47550 18050 47570 18420
rect 47650 18390 47960 18420
rect 48020 18390 48030 18450
rect 47650 18370 48030 18390
rect 47650 18310 47960 18370
rect 48020 18310 48030 18370
rect 47650 18280 48030 18310
rect 47650 18220 47960 18280
rect 48020 18220 48030 18280
rect 47650 18190 48030 18220
rect 47650 18130 47960 18190
rect 48020 18130 48030 18190
rect 47650 18110 48030 18130
rect 47650 18050 47960 18110
rect 48020 18050 48030 18110
rect 48640 18150 48740 18170
rect 48640 18090 48660 18150
rect 48720 18090 48740 18150
rect 48640 18070 48740 18090
rect 47550 18030 48030 18050
rect 48120 17450 48200 17460
rect 48120 17390 48130 17450
rect 48190 17390 48200 17450
rect 48120 17380 48200 17390
rect 41140 16810 41650 16820
rect 41140 16750 41150 16810
rect 41210 16750 41580 16810
rect 41640 16750 41650 16810
rect 41140 16740 41650 16750
rect 43240 16810 45420 16820
rect 43240 16750 43250 16810
rect 43310 16750 45350 16810
rect 45410 16750 45420 16810
rect 43240 16740 45420 16750
rect 47560 16760 48880 16770
rect 47560 16680 47570 16760
rect 47650 16750 48880 16760
rect 47650 16690 48800 16750
rect 48860 16690 48880 16750
rect 47650 16680 48880 16690
rect 47560 16670 48880 16680
rect 47950 16050 49070 16060
rect 47950 15990 47960 16050
rect 48020 15990 49000 16050
rect 49060 15990 49070 16050
rect 47950 15980 49070 15990
rect 46350 15350 48880 15370
rect 46350 15290 46360 15350
rect 46420 15290 46440 15350
rect 46500 15290 46520 15350
rect 46580 15290 48800 15350
rect 48860 15290 48880 15350
rect 46350 15270 48880 15290
rect 45340 14800 46320 14810
rect 45340 14740 45350 14800
rect 45410 14740 46010 14800
rect 46070 14740 46250 14800
rect 46310 14740 46320 14800
rect 45340 14730 46320 14740
rect 40350 14720 45020 14730
rect 40350 14660 40360 14720
rect 40420 14660 44590 14720
rect 44650 14660 44680 14720
rect 44740 14660 44770 14720
rect 44830 14660 44860 14720
rect 44920 14660 44950 14720
rect 45010 14660 45020 14720
rect 40350 14650 45020 14660
rect 41140 14410 41980 14420
rect 41140 14350 41150 14410
rect 41210 14402 41980 14410
rect 41210 14350 41560 14402
rect 41960 14350 41980 14402
rect 41140 14340 41980 14350
rect 44580 14410 46230 14420
rect 44580 14402 46160 14410
rect 44580 14350 44600 14402
rect 45000 14350 46160 14402
rect 46220 14350 46230 14410
rect 44580 14340 46230 14350
rect 39680 14090 46860 14100
rect 39680 14030 39690 14090
rect 39750 14030 46790 14090
rect 46850 14030 46860 14090
rect 39680 14020 46860 14030
rect 40620 13980 48730 13990
rect 40620 13920 40630 13980
rect 40690 13920 41040 13980
rect 41100 13920 48660 13980
rect 48720 13920 48730 13980
rect 40620 13910 48730 13920
rect 45470 13850 45550 13860
rect 39460 13810 41160 13820
rect 39460 13750 39470 13810
rect 39530 13750 41090 13810
rect 41150 13750 41160 13810
rect 39460 13740 41160 13750
rect 45470 13790 45480 13850
rect 45540 13790 45550 13850
rect 45470 13770 45550 13790
rect 45470 13710 45480 13770
rect 45540 13710 45550 13770
rect 45470 13700 45550 13710
rect 41160 13640 41240 13650
rect 41160 13580 41170 13640
rect 41230 13630 41240 13640
rect 41320 13640 41400 13650
rect 41320 13630 41330 13640
rect 41230 13590 41330 13630
rect 41230 13580 41240 13590
rect 41160 13570 41240 13580
rect 41320 13580 41330 13590
rect 41390 13630 41400 13640
rect 41480 13640 41560 13650
rect 41480 13630 41490 13640
rect 41390 13590 41490 13630
rect 41390 13580 41400 13590
rect 41320 13570 41400 13580
rect 41480 13580 41490 13590
rect 41550 13630 41560 13640
rect 41640 13640 41720 13650
rect 41640 13630 41650 13640
rect 41550 13590 41650 13630
rect 41550 13580 41560 13590
rect 41480 13570 41560 13580
rect 41640 13580 41650 13590
rect 41710 13630 41720 13640
rect 41800 13640 41880 13650
rect 41800 13630 41810 13640
rect 41710 13590 41810 13630
rect 41710 13580 41720 13590
rect 41640 13570 41720 13580
rect 41800 13580 41810 13590
rect 41870 13630 41880 13640
rect 41960 13640 42040 13650
rect 41960 13630 41970 13640
rect 41870 13590 41970 13630
rect 41870 13580 41880 13590
rect 41800 13570 41880 13580
rect 41960 13580 41970 13590
rect 42030 13630 42040 13640
rect 42120 13640 42200 13650
rect 42120 13630 42130 13640
rect 42030 13590 42130 13630
rect 42030 13580 42040 13590
rect 41960 13570 42040 13580
rect 42120 13580 42130 13590
rect 42190 13630 42200 13640
rect 42280 13640 42360 13650
rect 42280 13630 42290 13640
rect 42190 13590 42290 13630
rect 42190 13580 42200 13590
rect 42120 13570 42200 13580
rect 42280 13580 42290 13590
rect 42350 13630 42360 13640
rect 42440 13640 42520 13650
rect 42440 13630 42450 13640
rect 42350 13590 42450 13630
rect 42350 13580 42360 13590
rect 42280 13570 42360 13580
rect 42440 13580 42450 13590
rect 42510 13630 42520 13640
rect 42600 13640 42680 13650
rect 42600 13630 42610 13640
rect 42510 13590 42610 13630
rect 42510 13580 42520 13590
rect 42440 13570 42520 13580
rect 42600 13580 42610 13590
rect 42670 13630 42680 13640
rect 42760 13640 42840 13650
rect 42760 13630 42770 13640
rect 42670 13590 42770 13630
rect 42670 13580 42680 13590
rect 42600 13570 42680 13580
rect 42760 13580 42770 13590
rect 42830 13630 42840 13640
rect 42920 13640 43000 13650
rect 42920 13630 42930 13640
rect 42830 13590 42930 13630
rect 42830 13580 42840 13590
rect 42760 13570 42840 13580
rect 42920 13580 42930 13590
rect 42990 13630 43000 13640
rect 43080 13640 43160 13650
rect 43080 13630 43090 13640
rect 42990 13590 43090 13630
rect 42990 13580 43000 13590
rect 42920 13570 43000 13580
rect 43080 13580 43090 13590
rect 43150 13580 43160 13640
rect 43080 13570 43160 13580
rect 43240 13640 43320 13650
rect 43240 13580 43250 13640
rect 43310 13630 43320 13640
rect 43400 13640 43480 13650
rect 43400 13630 43410 13640
rect 43310 13590 43410 13630
rect 43310 13580 43320 13590
rect 43240 13570 43320 13580
rect 43400 13580 43410 13590
rect 43470 13630 43480 13640
rect 43560 13640 43640 13650
rect 43560 13630 43570 13640
rect 43470 13590 43570 13630
rect 43470 13580 43480 13590
rect 43400 13570 43480 13580
rect 43560 13580 43570 13590
rect 43630 13630 43640 13640
rect 43720 13640 43800 13650
rect 43720 13630 43730 13640
rect 43630 13590 43730 13630
rect 43630 13580 43640 13590
rect 43560 13570 43640 13580
rect 43720 13580 43730 13590
rect 43790 13630 43800 13640
rect 43880 13640 43960 13650
rect 43880 13630 43890 13640
rect 43790 13590 43890 13630
rect 43790 13580 43800 13590
rect 43720 13570 43800 13580
rect 43880 13580 43890 13590
rect 43950 13630 43960 13640
rect 44040 13640 44120 13650
rect 44040 13630 44050 13640
rect 43950 13590 44050 13630
rect 43950 13580 43960 13590
rect 43880 13570 43960 13580
rect 44040 13580 44050 13590
rect 44110 13630 44120 13640
rect 44200 13640 44280 13650
rect 44200 13630 44210 13640
rect 44110 13590 44210 13630
rect 44110 13580 44120 13590
rect 44040 13570 44120 13580
rect 44200 13580 44210 13590
rect 44270 13630 44280 13640
rect 44360 13640 44440 13650
rect 44360 13630 44370 13640
rect 44270 13590 44370 13630
rect 44270 13580 44280 13590
rect 44200 13570 44280 13580
rect 44360 13580 44370 13590
rect 44430 13630 44440 13640
rect 44520 13640 44600 13650
rect 44520 13630 44530 13640
rect 44430 13590 44530 13630
rect 44430 13580 44440 13590
rect 44360 13570 44440 13580
rect 44520 13580 44530 13590
rect 44590 13630 44600 13640
rect 44680 13640 44760 13650
rect 44680 13630 44690 13640
rect 44590 13590 44690 13630
rect 44590 13580 44600 13590
rect 44520 13570 44600 13580
rect 44680 13580 44690 13590
rect 44750 13630 44760 13640
rect 44840 13640 44920 13650
rect 44840 13630 44850 13640
rect 44750 13590 44850 13630
rect 44750 13580 44760 13590
rect 44680 13570 44760 13580
rect 44840 13580 44850 13590
rect 44910 13630 44920 13640
rect 45000 13640 45080 13650
rect 45000 13630 45010 13640
rect 44910 13590 45010 13630
rect 44910 13580 44920 13590
rect 44840 13570 44920 13580
rect 45000 13580 45010 13590
rect 45070 13630 45080 13640
rect 45160 13640 45240 13650
rect 45160 13630 45170 13640
rect 45070 13590 45170 13630
rect 45070 13580 45080 13590
rect 45000 13570 45080 13580
rect 45160 13580 45170 13590
rect 45230 13580 45240 13640
rect 45160 13570 45240 13580
rect 41900 13530 44660 13540
rect 41900 13470 41910 13530
rect 41970 13470 43170 13530
rect 43230 13470 43250 13530
rect 43310 13470 43330 13530
rect 43390 13470 44590 13530
rect 44650 13470 44660 13530
rect 41900 13450 44660 13470
rect 41900 13390 41910 13450
rect 41970 13390 43170 13450
rect 43230 13390 43250 13450
rect 43310 13390 43330 13450
rect 43390 13390 44590 13450
rect 44650 13390 44660 13450
rect 41900 13370 44660 13390
rect 41900 13310 41910 13370
rect 41970 13310 43170 13370
rect 43230 13310 43250 13370
rect 43310 13310 43330 13370
rect 43390 13310 44590 13370
rect 44650 13310 44660 13370
rect 41900 13300 44660 13310
rect 40920 12730 45640 12740
rect 40920 12670 40930 12730
rect 40990 12670 41170 12730
rect 41230 12670 41410 12730
rect 41470 12670 41650 12730
rect 41710 12670 42290 12730
rect 42350 12670 42530 12730
rect 42590 12670 42770 12730
rect 42830 12670 43730 12730
rect 43790 12670 43970 12730
rect 44030 12670 44210 12730
rect 44270 12670 44850 12730
rect 44910 12670 45090 12730
rect 45150 12670 45330 12730
rect 45390 12670 45570 12730
rect 45630 12670 45640 12730
rect 40920 12650 45640 12670
rect 40920 12590 40930 12650
rect 40990 12590 41170 12650
rect 41230 12590 41410 12650
rect 41470 12590 41650 12650
rect 41710 12590 42290 12650
rect 42350 12590 42530 12650
rect 42590 12590 42770 12650
rect 42830 12590 43730 12650
rect 43790 12590 43970 12650
rect 44030 12590 44210 12650
rect 44270 12590 44850 12650
rect 44910 12590 45090 12650
rect 45150 12590 45330 12650
rect 45390 12590 45570 12650
rect 45630 12590 45640 12650
rect 40920 12570 45640 12590
rect 40920 12510 40930 12570
rect 40990 12510 41170 12570
rect 41230 12510 41410 12570
rect 41470 12510 41650 12570
rect 41710 12510 42290 12570
rect 42350 12510 42530 12570
rect 42590 12510 42770 12570
rect 42830 12510 43730 12570
rect 43790 12510 43970 12570
rect 44030 12510 44210 12570
rect 44270 12510 44850 12570
rect 44910 12510 45090 12570
rect 45150 12510 45330 12570
rect 45390 12510 45570 12570
rect 45630 12510 45640 12570
rect 40920 12500 45640 12510
rect 40740 12460 42530 12470
rect 40740 12400 40750 12460
rect 40810 12400 41500 12460
rect 41560 12400 41720 12460
rect 41780 12400 41980 12460
rect 42040 12400 42200 12460
rect 42260 12400 42460 12460
rect 42520 12400 42530 12460
rect 40740 12390 42530 12400
rect 44030 12460 45820 12470
rect 44030 12400 44040 12460
rect 44100 12400 44300 12460
rect 44360 12400 44520 12460
rect 44580 12400 44780 12460
rect 44840 12400 45000 12460
rect 45060 12400 45750 12460
rect 45810 12400 45820 12460
rect 44030 12390 45820 12400
rect 39680 12350 42449 12360
rect 39680 12290 39690 12350
rect 39750 12298 41433 12350
rect 41485 12298 41793 12350
rect 41845 12298 41913 12350
rect 41965 12298 42273 12350
rect 42325 12298 42393 12350
rect 42445 12298 42449 12350
rect 44111 12350 46230 12360
rect 39750 12290 42449 12298
rect 42800 12330 43760 12340
rect 39680 12280 39760 12290
rect 42800 12270 42810 12330
rect 42870 12270 43170 12330
rect 43230 12270 43250 12330
rect 43310 12270 43330 12330
rect 43390 12270 43690 12330
rect 43750 12270 43760 12330
rect 44111 12298 44115 12350
rect 44167 12298 44235 12350
rect 44287 12298 44595 12350
rect 44647 12298 44715 12350
rect 44767 12298 45075 12350
rect 45127 12298 46160 12350
rect 44111 12290 46160 12298
rect 46220 12290 46230 12350
rect 46150 12280 46230 12290
rect 42800 12250 43760 12270
rect 42800 12190 42810 12250
rect 42870 12190 43170 12250
rect 43230 12190 43250 12250
rect 43310 12190 43330 12250
rect 43390 12190 43690 12250
rect 43750 12190 43760 12250
rect 42800 12170 43760 12190
rect 39570 12122 42550 12130
rect 39570 12120 41536 12122
rect 39570 12060 39580 12120
rect 39640 12070 41536 12120
rect 41588 12070 41694 12122
rect 41746 12070 42018 12122
rect 42070 12070 42172 12122
rect 42224 12070 42496 12122
rect 42548 12070 42550 12122
rect 42800 12110 42810 12170
rect 42870 12110 43170 12170
rect 43230 12110 43250 12170
rect 43310 12110 43330 12170
rect 43390 12110 43690 12170
rect 43750 12110 43760 12170
rect 42800 12100 43760 12110
rect 44010 12122 46320 12130
rect 39640 12060 42550 12070
rect 44010 12070 44012 12122
rect 44064 12070 44336 12122
rect 44388 12070 44490 12122
rect 44542 12070 44814 12122
rect 44866 12070 44972 12122
rect 45024 12120 46320 12122
rect 45024 12070 46250 12120
rect 44010 12060 46250 12070
rect 46310 12060 46320 12120
rect 39570 12050 39650 12060
rect 46240 12050 46320 12060
rect 41600 12020 42640 12030
rect 41600 11960 41610 12020
rect 41670 11960 42090 12020
rect 42150 11960 42570 12020
rect 42630 11960 42640 12020
rect 41600 11950 42640 11960
rect 43920 12020 44960 12030
rect 43920 11960 43930 12020
rect 43990 11960 44410 12020
rect 44470 11960 44890 12020
rect 44950 11960 44960 12020
rect 43920 11950 44960 11960
rect 41360 11910 42400 11920
rect 41360 11850 41370 11910
rect 41430 11850 41850 11910
rect 41910 11850 42330 11910
rect 42390 11850 42400 11910
rect 41360 11840 42400 11850
rect 44160 11910 45200 11920
rect 44160 11850 44170 11910
rect 44230 11850 44650 11910
rect 44710 11850 45130 11910
rect 45190 11850 45200 11910
rect 44160 11840 45200 11850
rect 43740 11800 46590 11810
rect 43740 11740 43750 11800
rect 43810 11740 43930 11800
rect 43990 11740 44170 11800
rect 44230 11740 44410 11800
rect 44470 11740 44650 11800
rect 44710 11740 45130 11800
rect 45190 11740 45370 11800
rect 45430 11740 45790 11800
rect 45850 11740 46360 11800
rect 46420 11740 46440 11800
rect 46500 11740 46520 11800
rect 46580 11740 46590 11800
rect 43740 11720 46590 11740
rect 43740 11660 43750 11720
rect 43810 11660 43930 11720
rect 43990 11660 44170 11720
rect 44230 11660 44410 11720
rect 44470 11660 44650 11720
rect 44710 11660 45130 11720
rect 45190 11660 45370 11720
rect 45430 11660 45790 11720
rect 45850 11660 46360 11720
rect 46420 11660 46440 11720
rect 46500 11660 46520 11720
rect 46580 11660 46590 11720
rect 40620 11640 42820 11650
rect 40620 11580 40630 11640
rect 40690 11580 40710 11640
rect 40770 11580 41130 11640
rect 41190 11580 41370 11640
rect 41430 11580 41850 11640
rect 41910 11580 42090 11640
rect 42150 11580 42570 11640
rect 42630 11580 42750 11640
rect 42810 11580 42820 11640
rect 40620 11570 42820 11580
rect 43740 11640 46590 11660
rect 43740 11580 43750 11640
rect 43810 11580 43930 11640
rect 43990 11580 44170 11640
rect 44230 11580 44410 11640
rect 44470 11580 44650 11640
rect 44710 11580 45130 11640
rect 45190 11580 45370 11640
rect 45430 11580 45790 11640
rect 45850 11580 46360 11640
rect 46420 11580 46440 11640
rect 46500 11580 46520 11640
rect 46580 11580 46590 11640
rect 43740 11570 46590 11580
rect 40880 11520 40960 11530
rect 40880 11460 40890 11520
rect 40950 11510 40960 11520
rect 41600 11520 41680 11530
rect 41600 11510 41610 11520
rect 40950 11470 41610 11510
rect 40950 11460 40960 11470
rect 40880 11450 40960 11460
rect 41600 11460 41610 11470
rect 41670 11510 41680 11520
rect 42320 11520 42400 11530
rect 42320 11510 42330 11520
rect 41670 11470 42330 11510
rect 41670 11460 41680 11470
rect 41600 11450 41680 11460
rect 42320 11460 42330 11470
rect 42390 11460 42400 11520
rect 42320 11450 42400 11460
rect 44160 11520 44240 11530
rect 44160 11460 44170 11520
rect 44230 11510 44240 11520
rect 44880 11520 44960 11530
rect 44880 11510 44890 11520
rect 44230 11470 44890 11510
rect 44230 11460 44240 11470
rect 44160 11450 44240 11460
rect 44880 11460 44890 11470
rect 44950 11510 44960 11520
rect 45600 11520 45680 11530
rect 45600 11510 45610 11520
rect 44950 11470 45610 11510
rect 44950 11460 44960 11470
rect 44880 11450 44960 11460
rect 45600 11460 45610 11470
rect 45670 11460 45680 11520
rect 45600 11450 45680 11460
rect 41370 11190 41430 11220
rect 45130 11190 45190 11230
rect 38790 11180 43140 11190
rect 38790 11120 38800 11180
rect 38860 11120 40650 11180
rect 40710 11120 41370 11180
rect 41430 11120 42090 11180
rect 42150 11120 42810 11180
rect 42870 11120 43070 11180
rect 43130 11120 43140 11180
rect 38790 11110 43140 11120
rect 43420 11180 47650 11190
rect 43420 11120 43430 11180
rect 43490 11120 43690 11180
rect 43750 11120 44410 11180
rect 44470 11120 45130 11180
rect 45190 11120 45850 11180
rect 45910 11120 47580 11180
rect 47640 11120 47650 11180
rect 43420 11110 47650 11120
rect 40520 11070 46040 11080
rect 40520 11010 40530 11070
rect 40590 11010 40770 11070
rect 40830 11010 41010 11070
rect 41070 11010 41250 11070
rect 41310 11010 41490 11070
rect 41550 11010 41730 11070
rect 41790 11010 41970 11070
rect 42030 11010 42210 11070
rect 42270 11010 42450 11070
rect 42510 11010 42690 11070
rect 42750 11010 42930 11070
rect 42990 11010 43570 11070
rect 43630 11010 43810 11070
rect 43870 11010 44050 11070
rect 44110 11010 44290 11070
rect 44350 11010 44530 11070
rect 44590 11010 44770 11070
rect 44830 11010 45010 11070
rect 45070 11010 45250 11070
rect 45310 11010 45490 11070
rect 45550 11010 45730 11070
rect 45790 11010 45970 11070
rect 46030 11010 46040 11070
rect 40520 10990 46040 11010
rect 40520 10930 40530 10990
rect 40590 10930 40770 10990
rect 40830 10930 41010 10990
rect 41070 10930 41250 10990
rect 41310 10930 41490 10990
rect 41550 10930 41730 10990
rect 41790 10930 41970 10990
rect 42030 10930 42210 10990
rect 42270 10930 42450 10990
rect 42510 10930 42690 10990
rect 42750 10930 42930 10990
rect 42990 10930 43570 10990
rect 43630 10930 43810 10990
rect 43870 10930 44050 10990
rect 44110 10930 44290 10990
rect 44350 10930 44530 10990
rect 44590 10930 44770 10990
rect 44830 10930 45010 10990
rect 45070 10930 45250 10990
rect 45310 10930 45490 10990
rect 45550 10930 45730 10990
rect 45790 10930 45970 10990
rect 46030 10930 46040 10990
rect 40520 10910 46040 10930
rect 40520 10850 40530 10910
rect 40590 10850 40770 10910
rect 40830 10850 41010 10910
rect 41070 10850 41250 10910
rect 41310 10850 41490 10910
rect 41550 10850 41730 10910
rect 41790 10850 41970 10910
rect 42030 10850 42210 10910
rect 42270 10850 42450 10910
rect 42510 10850 42690 10910
rect 42750 10850 42930 10910
rect 42990 10850 43570 10910
rect 43630 10850 43810 10910
rect 43870 10850 44050 10910
rect 44110 10850 44290 10910
rect 44350 10850 44530 10910
rect 44590 10850 44770 10910
rect 44830 10850 45010 10910
rect 45070 10850 45250 10910
rect 45310 10850 45490 10910
rect 45550 10850 45730 10910
rect 45790 10850 45970 10910
rect 46030 10850 46040 10910
rect 40520 10840 46040 10850
rect 39570 10800 44760 10810
rect 39570 10740 39580 10800
rect 39640 10740 41810 10800
rect 41870 10740 43250 10800
rect 43310 10740 44690 10800
rect 44750 10740 44760 10800
rect 39570 10730 44760 10740
rect 39460 10690 45790 10700
rect 39460 10630 39470 10690
rect 39530 10630 42170 10690
rect 42230 10630 44330 10690
rect 44390 10630 45720 10690
rect 45780 10630 45790 10690
rect 39460 10620 45790 10630
rect 42520 10580 46320 10590
rect 42520 10520 42530 10580
rect 42590 10520 43970 10580
rect 44030 10520 45250 10580
rect 45310 10520 46250 10580
rect 46310 10520 46320 10580
rect 42520 10510 46320 10520
rect 42880 10470 46230 10480
rect 42880 10410 42890 10470
rect 42950 10410 43610 10470
rect 43670 10410 46160 10470
rect 46220 10410 46230 10470
rect 42880 10400 46230 10410
rect 41900 10360 44660 10370
rect 41960 10300 42080 10360
rect 42140 10300 42260 10360
rect 42320 10300 42440 10360
rect 42500 10300 42620 10360
rect 42680 10300 42800 10360
rect 42860 10300 42980 10360
rect 43040 10300 43160 10360
rect 43220 10300 43340 10360
rect 43400 10300 43430 10360
rect 43490 10300 43520 10360
rect 43580 10300 43700 10360
rect 43760 10300 43880 10360
rect 43940 10300 44060 10360
rect 44120 10300 44240 10360
rect 44300 10300 44420 10360
rect 44480 10300 44600 10360
rect 41900 10290 44660 10300
rect 45590 10160 45910 10170
rect 45590 10100 45600 10160
rect 45660 10100 45840 10160
rect 45900 10100 45910 10160
rect 45590 10090 45910 10100
rect 45240 9820 45320 9830
rect 45240 9760 45250 9820
rect 45310 9810 45320 9820
rect 45710 9820 45790 9830
rect 45710 9810 45720 9820
rect 45310 9770 45720 9810
rect 45310 9760 45320 9770
rect 45240 9750 45320 9760
rect 45710 9760 45720 9770
rect 45780 9760 45790 9820
rect 45710 9750 45790 9760
rect 41620 9620 46010 9630
rect 41620 9560 41630 9620
rect 41690 9560 41990 9620
rect 42050 9560 42350 9620
rect 42410 9560 42710 9620
rect 42770 9560 43070 9620
rect 43130 9560 43430 9620
rect 43490 9560 43790 9620
rect 43850 9560 44150 9620
rect 44210 9560 44510 9620
rect 44570 9560 44870 9620
rect 44930 9560 45500 9620
rect 45560 9560 45940 9620
rect 46000 9560 46010 9620
rect 41620 9540 46010 9560
rect 41620 9480 41630 9540
rect 41690 9480 41990 9540
rect 42050 9480 42350 9540
rect 42410 9480 42710 9540
rect 42770 9480 43070 9540
rect 43130 9480 43430 9540
rect 43490 9480 43790 9540
rect 43850 9480 44150 9540
rect 44210 9480 44510 9540
rect 44570 9480 44870 9540
rect 44930 9480 45500 9540
rect 45560 9480 45940 9540
rect 46000 9480 46010 9540
rect 41620 9460 46010 9480
rect 41620 9400 41630 9460
rect 41690 9400 41990 9460
rect 42050 9400 42350 9460
rect 42410 9400 42710 9460
rect 42770 9400 43070 9460
rect 43130 9400 43430 9460
rect 43490 9400 43790 9460
rect 43850 9400 44150 9460
rect 44210 9400 44510 9460
rect 44570 9400 44870 9460
rect 44930 9400 45500 9460
rect 45560 9400 45940 9460
rect 46000 9400 46010 9460
rect 41620 9390 46010 9400
rect 38790 9300 38800 9360
rect 38860 9350 44754 9360
rect 38860 9300 41808 9350
rect 38790 9298 41808 9300
rect 41860 9298 41918 9350
rect 41970 9298 42028 9350
rect 42080 9298 42138 9350
rect 42190 9298 42248 9350
rect 42300 9298 42358 9350
rect 42410 9298 42468 9350
rect 42520 9298 42578 9350
rect 42630 9298 42688 9350
rect 42740 9298 42798 9350
rect 42850 9298 43708 9350
rect 43760 9298 43818 9350
rect 43870 9298 43928 9350
rect 43980 9298 44038 9350
rect 44090 9298 44148 9350
rect 44200 9298 44258 9350
rect 44310 9298 44368 9350
rect 44420 9298 44478 9350
rect 44530 9298 44588 9350
rect 44640 9298 44698 9350
rect 44750 9298 44754 9350
rect 38790 9290 44754 9298
rect 41630 9020 44930 9030
rect 41630 8960 41640 9020
rect 41700 8960 41860 9020
rect 41920 8960 42080 9020
rect 42140 8960 42300 9020
rect 42360 8960 42520 9020
rect 42580 8960 42740 9020
rect 42800 8960 42960 9020
rect 43020 8960 43540 9020
rect 43600 8960 43760 9020
rect 43820 8960 43980 9020
rect 44040 8960 44200 9020
rect 44260 8960 44420 9020
rect 44480 8960 44640 9020
rect 44700 8960 44860 9020
rect 44920 8960 44930 9020
rect 41630 8950 44930 8960
rect 39680 8910 42920 8920
rect 39680 8850 39690 8910
rect 39750 8850 41750 8910
rect 41810 8850 41970 8910
rect 42030 8850 42190 8910
rect 42250 8850 42410 8910
rect 42470 8850 42630 8910
rect 42690 8850 42850 8910
rect 42910 8850 42920 8910
rect 39680 8840 42920 8850
rect 43640 8900 44820 8910
rect 43640 8840 43650 8900
rect 43710 8840 43870 8900
rect 43930 8840 44090 8900
rect 44150 8840 44310 8900
rect 44370 8840 44530 8900
rect 44590 8840 44750 8900
rect 44810 8840 44820 8900
rect 43640 8820 44820 8840
rect 43640 8760 43650 8820
rect 43710 8760 43870 8820
rect 43930 8760 44090 8820
rect 44150 8760 44310 8820
rect 44370 8760 44530 8820
rect 44590 8760 44750 8820
rect 44810 8760 44820 8820
rect 43640 8740 44820 8760
rect 43640 8680 43650 8740
rect 43710 8680 43870 8740
rect 43930 8680 44090 8740
rect 44150 8680 44310 8740
rect 44370 8680 44530 8740
rect 44590 8680 44750 8740
rect 44810 8680 44820 8740
rect 43640 8670 44820 8680
<< via2 >>
rect 48200 18790 48260 18850
rect 48660 18090 48720 18150
rect 48130 17390 48190 17450
rect 48800 16690 48860 16750
rect 49000 15990 49060 16050
rect 48800 15290 48860 15350
<< metal3 >>
rect 49120 18870 49580 19040
rect 49820 18870 50280 19040
rect 50520 18870 50980 19040
rect 51220 18870 51680 19040
rect 51920 18870 52380 19040
rect 52620 18870 53080 19040
rect 53320 18870 53780 19040
rect 54020 18870 54480 19040
rect 54720 18870 55180 19040
rect 55420 18870 55880 19040
rect 49120 18860 55880 18870
rect 48190 18850 55880 18860
rect 48190 18790 48200 18850
rect 48260 18790 55880 18850
rect 48190 18780 55880 18790
rect 49120 18770 55880 18780
rect 49120 18580 49580 18770
rect 49820 18580 50280 18770
rect 50520 18580 50980 18770
rect 51220 18580 51680 18770
rect 51920 18580 52380 18770
rect 52620 18580 53080 18770
rect 53320 18580 53780 18770
rect 54020 18580 54480 18770
rect 54720 18580 55180 18770
rect 55420 18580 55880 18770
rect 55600 18340 55700 18580
rect 49120 18170 49580 18340
rect 49820 18170 50280 18340
rect 50520 18170 50980 18340
rect 51220 18170 51680 18340
rect 51920 18170 52380 18340
rect 52620 18170 53080 18340
rect 53320 18170 53780 18340
rect 54020 18170 54480 18340
rect 54720 18170 55180 18340
rect 55420 18170 55880 18340
rect 48640 18160 48740 18170
rect 48640 18080 48650 18160
rect 48730 18080 48740 18160
rect 48640 18070 48740 18080
rect 49120 18070 55880 18170
rect 49120 17880 49580 18070
rect 49820 17880 50280 18070
rect 50520 17880 50980 18070
rect 51220 17880 51680 18070
rect 51920 17880 52380 18070
rect 52620 17880 53080 18070
rect 53320 17880 53780 18070
rect 54020 17880 54480 18070
rect 54720 17880 55180 18070
rect 55420 17880 55880 18070
rect 49120 17470 49580 17640
rect 49820 17470 50280 17640
rect 50520 17470 50980 17640
rect 51220 17470 51680 17640
rect 51920 17470 52380 17640
rect 52620 17470 53080 17640
rect 53320 17470 53780 17640
rect 54020 17470 54480 17640
rect 54720 17470 55180 17640
rect 55420 17470 55880 17640
rect 49120 17460 55880 17470
rect 48120 17450 55880 17460
rect 48120 17390 48130 17450
rect 48190 17390 55880 17450
rect 48120 17380 55880 17390
rect 49120 17370 55880 17380
rect 49120 17180 49580 17370
rect 49820 17180 50280 17370
rect 50520 17180 50980 17370
rect 51220 17180 51680 17370
rect 51920 17180 52380 17370
rect 52620 17180 53080 17370
rect 53320 17180 53780 17370
rect 54020 17180 54480 17370
rect 54720 17180 55180 17370
rect 55420 17180 55880 17370
rect 55600 16940 55700 17180
rect 49120 16770 49580 16940
rect 49820 16770 50280 16940
rect 50520 16770 50980 16940
rect 51220 16770 51680 16940
rect 51920 16770 52380 16940
rect 52620 16770 53080 16940
rect 53320 16770 53780 16940
rect 54020 16770 54480 16940
rect 54720 16770 55180 16940
rect 55420 16770 55880 16940
rect 48780 16760 48880 16770
rect 48780 16680 48790 16760
rect 48870 16680 48880 16760
rect 48780 16670 48880 16680
rect 49120 16670 55880 16770
rect 49120 16480 49580 16670
rect 49820 16480 50280 16670
rect 50520 16480 50980 16670
rect 51220 16480 51680 16670
rect 51920 16480 52380 16670
rect 52620 16480 53080 16670
rect 53320 16480 53780 16670
rect 54020 16480 54480 16670
rect 54720 16480 55180 16670
rect 55420 16480 55880 16670
rect 49120 16070 49580 16240
rect 49820 16070 50280 16240
rect 50520 16070 50980 16240
rect 51220 16070 51680 16240
rect 51920 16070 52380 16240
rect 52620 16070 53080 16240
rect 53320 16070 53780 16240
rect 54020 16070 54480 16240
rect 54720 16070 55180 16240
rect 55420 16070 55880 16240
rect 49120 16060 55880 16070
rect 48990 16050 55880 16060
rect 48990 15990 49000 16050
rect 49060 15990 55880 16050
rect 48990 15980 55880 15990
rect 49120 15970 55880 15980
rect 49120 15780 49580 15970
rect 49820 15780 50280 15970
rect 50520 15780 50980 15970
rect 51220 15780 51680 15970
rect 51920 15780 52380 15970
rect 52620 15780 53080 15970
rect 53320 15780 53780 15970
rect 54020 15780 54480 15970
rect 54720 15780 55180 15970
rect 55420 15780 55880 15970
rect 55600 15540 55700 15780
rect 49120 15370 49580 15540
rect 49820 15370 50280 15540
rect 50520 15370 50980 15540
rect 51220 15370 51680 15540
rect 51920 15370 52380 15540
rect 52620 15370 53080 15540
rect 53320 15370 53780 15540
rect 54020 15370 54480 15540
rect 54720 15370 55180 15540
rect 55420 15370 55880 15540
rect 48780 15360 48880 15370
rect 48780 15280 48790 15360
rect 48870 15280 48880 15360
rect 48780 15270 48880 15280
rect 49120 15270 55880 15370
rect 49120 15080 49580 15270
rect 49820 15080 50280 15270
rect 50520 15080 50980 15270
rect 51220 15080 51680 15270
rect 51920 15080 52380 15270
rect 52620 15080 53080 15270
rect 53320 15080 53780 15270
rect 54020 15080 54480 15270
rect 54720 15080 55180 15270
rect 55420 15080 55880 15270
<< via3 >>
rect 48650 18150 48730 18160
rect 48650 18090 48660 18150
rect 48660 18090 48720 18150
rect 48720 18090 48730 18150
rect 48650 18080 48730 18090
rect 48790 16750 48870 16760
rect 48790 16690 48800 16750
rect 48800 16690 48860 16750
rect 48860 16690 48870 16750
rect 48790 16680 48870 16690
rect 48790 15350 48870 15360
rect 48790 15290 48800 15350
rect 48800 15290 48860 15350
rect 48860 15290 48870 15350
rect 48790 15280 48870 15290
<< mimcap >>
rect 49150 18860 49550 19010
rect 49150 18780 49320 18860
rect 49400 18780 49550 18860
rect 49150 18610 49550 18780
rect 49850 18860 50250 19010
rect 49850 18780 50010 18860
rect 50090 18780 50250 18860
rect 49850 18610 50250 18780
rect 50550 18860 50950 19010
rect 50550 18780 50710 18860
rect 50790 18780 50950 18860
rect 50550 18610 50950 18780
rect 51250 18860 51650 19010
rect 51250 18780 51410 18860
rect 51490 18780 51650 18860
rect 51250 18610 51650 18780
rect 51950 18860 52350 19010
rect 51950 18780 52110 18860
rect 52190 18780 52350 18860
rect 51950 18610 52350 18780
rect 52650 18860 53050 19010
rect 52650 18780 52810 18860
rect 52890 18780 53050 18860
rect 52650 18610 53050 18780
rect 53350 18860 53750 19010
rect 53350 18780 53510 18860
rect 53590 18780 53750 18860
rect 53350 18610 53750 18780
rect 54050 18860 54450 19010
rect 54050 18780 54210 18860
rect 54290 18780 54450 18860
rect 54050 18610 54450 18780
rect 54750 18860 55150 19010
rect 54750 18780 54910 18860
rect 54990 18780 55150 18860
rect 54750 18610 55150 18780
rect 55450 18860 55850 19010
rect 55450 18780 55610 18860
rect 55690 18780 55850 18860
rect 55450 18610 55850 18780
rect 49150 18160 49550 18310
rect 49150 18080 49320 18160
rect 49400 18080 49550 18160
rect 49150 17910 49550 18080
rect 49850 18160 50250 18310
rect 49850 18080 50010 18160
rect 50090 18080 50250 18160
rect 49850 17910 50250 18080
rect 50550 18160 50950 18310
rect 50550 18080 50710 18160
rect 50790 18080 50950 18160
rect 50550 17910 50950 18080
rect 51250 18160 51650 18310
rect 51250 18080 51410 18160
rect 51490 18080 51650 18160
rect 51250 17910 51650 18080
rect 51950 18160 52350 18310
rect 51950 18080 52110 18160
rect 52190 18080 52350 18160
rect 51950 17910 52350 18080
rect 52650 18160 53050 18310
rect 52650 18080 52810 18160
rect 52890 18080 53050 18160
rect 52650 17910 53050 18080
rect 53350 18160 53750 18310
rect 53350 18080 53510 18160
rect 53590 18080 53750 18160
rect 53350 17910 53750 18080
rect 54050 18160 54450 18310
rect 54050 18080 54210 18160
rect 54290 18080 54450 18160
rect 54050 17910 54450 18080
rect 54750 18160 55150 18310
rect 54750 18080 54910 18160
rect 54990 18080 55150 18160
rect 54750 17910 55150 18080
rect 55450 18160 55850 18310
rect 55450 18080 55610 18160
rect 55690 18080 55850 18160
rect 55450 17910 55850 18080
rect 49150 17460 49550 17610
rect 49150 17380 49320 17460
rect 49400 17380 49550 17460
rect 49150 17210 49550 17380
rect 49850 17460 50250 17610
rect 49850 17380 50010 17460
rect 50090 17380 50250 17460
rect 49850 17210 50250 17380
rect 50550 17460 50950 17610
rect 50550 17380 50710 17460
rect 50790 17380 50950 17460
rect 50550 17210 50950 17380
rect 51250 17460 51650 17610
rect 51250 17380 51410 17460
rect 51490 17380 51650 17460
rect 51250 17210 51650 17380
rect 51950 17460 52350 17610
rect 51950 17380 52110 17460
rect 52190 17380 52350 17460
rect 51950 17210 52350 17380
rect 52650 17460 53050 17610
rect 52650 17380 52810 17460
rect 52890 17380 53050 17460
rect 52650 17210 53050 17380
rect 53350 17460 53750 17610
rect 53350 17380 53510 17460
rect 53590 17380 53750 17460
rect 53350 17210 53750 17380
rect 54050 17460 54450 17610
rect 54050 17380 54210 17460
rect 54290 17380 54450 17460
rect 54050 17210 54450 17380
rect 54750 17460 55150 17610
rect 54750 17380 54910 17460
rect 54990 17380 55150 17460
rect 54750 17210 55150 17380
rect 55450 17460 55850 17610
rect 55450 17380 55610 17460
rect 55690 17380 55850 17460
rect 55450 17210 55850 17380
rect 49150 16760 49550 16910
rect 49150 16680 49320 16760
rect 49400 16680 49550 16760
rect 49150 16510 49550 16680
rect 49850 16760 50250 16910
rect 49850 16680 50010 16760
rect 50090 16680 50250 16760
rect 49850 16510 50250 16680
rect 50550 16760 50950 16910
rect 50550 16680 50710 16760
rect 50790 16680 50950 16760
rect 50550 16510 50950 16680
rect 51250 16760 51650 16910
rect 51250 16680 51410 16760
rect 51490 16680 51650 16760
rect 51250 16510 51650 16680
rect 51950 16760 52350 16910
rect 51950 16680 52110 16760
rect 52190 16680 52350 16760
rect 51950 16510 52350 16680
rect 52650 16760 53050 16910
rect 52650 16680 52810 16760
rect 52890 16680 53050 16760
rect 52650 16510 53050 16680
rect 53350 16760 53750 16910
rect 53350 16680 53510 16760
rect 53590 16680 53750 16760
rect 53350 16510 53750 16680
rect 54050 16760 54450 16910
rect 54050 16680 54210 16760
rect 54290 16680 54450 16760
rect 54050 16510 54450 16680
rect 54750 16760 55150 16910
rect 54750 16680 54910 16760
rect 54990 16680 55150 16760
rect 54750 16510 55150 16680
rect 55450 16760 55850 16910
rect 55450 16680 55610 16760
rect 55690 16680 55850 16760
rect 55450 16510 55850 16680
rect 49150 16060 49550 16210
rect 49150 15980 49320 16060
rect 49400 15980 49550 16060
rect 49150 15810 49550 15980
rect 49850 16060 50250 16210
rect 49850 15980 50010 16060
rect 50090 15980 50250 16060
rect 49850 15810 50250 15980
rect 50550 16060 50950 16210
rect 50550 15980 50710 16060
rect 50790 15980 50950 16060
rect 50550 15810 50950 15980
rect 51250 16060 51650 16210
rect 51250 15980 51410 16060
rect 51490 15980 51650 16060
rect 51250 15810 51650 15980
rect 51950 16060 52350 16210
rect 51950 15980 52110 16060
rect 52190 15980 52350 16060
rect 51950 15810 52350 15980
rect 52650 16060 53050 16210
rect 52650 15980 52810 16060
rect 52890 15980 53050 16060
rect 52650 15810 53050 15980
rect 53350 16060 53750 16210
rect 53350 15980 53510 16060
rect 53590 15980 53750 16060
rect 53350 15810 53750 15980
rect 54050 16060 54450 16210
rect 54050 15980 54210 16060
rect 54290 15980 54450 16060
rect 54050 15810 54450 15980
rect 54750 16060 55150 16210
rect 54750 15980 54910 16060
rect 54990 15980 55150 16060
rect 54750 15810 55150 15980
rect 55450 16060 55850 16210
rect 55450 15980 55610 16060
rect 55690 15980 55850 16060
rect 55450 15810 55850 15980
rect 49150 15360 49550 15510
rect 49150 15280 49320 15360
rect 49400 15280 49550 15360
rect 49150 15110 49550 15280
rect 49850 15360 50250 15510
rect 49850 15280 50010 15360
rect 50090 15280 50250 15360
rect 49850 15110 50250 15280
rect 50550 15360 50950 15510
rect 50550 15280 50710 15360
rect 50790 15280 50950 15360
rect 50550 15110 50950 15280
rect 51250 15360 51650 15510
rect 51250 15280 51410 15360
rect 51490 15280 51650 15360
rect 51250 15110 51650 15280
rect 51950 15360 52350 15510
rect 51950 15280 52110 15360
rect 52190 15280 52350 15360
rect 51950 15110 52350 15280
rect 52650 15360 53050 15510
rect 52650 15280 52810 15360
rect 52890 15280 53050 15360
rect 52650 15110 53050 15280
rect 53350 15360 53750 15510
rect 53350 15280 53510 15360
rect 53590 15280 53750 15360
rect 53350 15110 53750 15280
rect 54050 15360 54450 15510
rect 54050 15280 54210 15360
rect 54290 15280 54450 15360
rect 54050 15110 54450 15280
rect 54750 15360 55150 15510
rect 54750 15280 54910 15360
rect 54990 15280 55150 15360
rect 54750 15110 55150 15280
rect 55450 15360 55850 15510
rect 55450 15280 55610 15360
rect 55690 15280 55850 15360
rect 55450 15110 55850 15280
<< mimcapcontact >>
rect 49320 18780 49400 18860
rect 50010 18780 50090 18860
rect 50710 18780 50790 18860
rect 51410 18780 51490 18860
rect 52110 18780 52190 18860
rect 52810 18780 52890 18860
rect 53510 18780 53590 18860
rect 54210 18780 54290 18860
rect 54910 18780 54990 18860
rect 55610 18780 55690 18860
rect 49320 18080 49400 18160
rect 50010 18080 50090 18160
rect 50710 18080 50790 18160
rect 51410 18080 51490 18160
rect 52110 18080 52190 18160
rect 52810 18080 52890 18160
rect 53510 18080 53590 18160
rect 54210 18080 54290 18160
rect 54910 18080 54990 18160
rect 55610 18080 55690 18160
rect 49320 17380 49400 17460
rect 50010 17380 50090 17460
rect 50710 17380 50790 17460
rect 51410 17380 51490 17460
rect 52110 17380 52190 17460
rect 52810 17380 52890 17460
rect 53510 17380 53590 17460
rect 54210 17380 54290 17460
rect 54910 17380 54990 17460
rect 55610 17380 55690 17460
rect 49320 16680 49400 16760
rect 50010 16680 50090 16760
rect 50710 16680 50790 16760
rect 51410 16680 51490 16760
rect 52110 16680 52190 16760
rect 52810 16680 52890 16760
rect 53510 16680 53590 16760
rect 54210 16680 54290 16760
rect 54910 16680 54990 16760
rect 55610 16680 55690 16760
rect 49320 15980 49400 16060
rect 50010 15980 50090 16060
rect 50710 15980 50790 16060
rect 51410 15980 51490 16060
rect 52110 15980 52190 16060
rect 52810 15980 52890 16060
rect 53510 15980 53590 16060
rect 54210 15980 54290 16060
rect 54910 15980 54990 16060
rect 55610 15980 55690 16060
rect 49320 15280 49400 15360
rect 50010 15280 50090 15360
rect 50710 15280 50790 15360
rect 51410 15280 51490 15360
rect 52110 15280 52190 15360
rect 52810 15280 52890 15360
rect 53510 15280 53590 15360
rect 54210 15280 54290 15360
rect 54910 15280 54990 15360
rect 55610 15280 55690 15360
<< metal4 >>
rect 49310 18860 55700 18870
rect 49310 18780 49320 18860
rect 49400 18780 50010 18860
rect 50090 18780 50710 18860
rect 50790 18780 51410 18860
rect 51490 18780 52110 18860
rect 52190 18780 52810 18860
rect 52890 18780 53510 18860
rect 53590 18780 54210 18860
rect 54290 18780 54910 18860
rect 54990 18780 55610 18860
rect 55690 18780 55700 18860
rect 49310 18770 55700 18780
rect 55600 18170 55700 18770
rect 48640 18160 55700 18170
rect 48640 18080 48650 18160
rect 48730 18080 49320 18160
rect 49400 18080 50010 18160
rect 50090 18080 50710 18160
rect 50790 18080 51410 18160
rect 51490 18080 52110 18160
rect 52190 18080 52810 18160
rect 52890 18080 53510 18160
rect 53590 18080 54210 18160
rect 54290 18080 54910 18160
rect 54990 18080 55610 18160
rect 55690 18080 55700 18160
rect 48640 18070 55700 18080
rect 49310 17460 55700 17470
rect 49310 17380 49320 17460
rect 49400 17380 50010 17460
rect 50090 17380 50710 17460
rect 50790 17380 51410 17460
rect 51490 17380 52110 17460
rect 52190 17380 52810 17460
rect 52890 17380 53510 17460
rect 53590 17380 54210 17460
rect 54290 17380 54910 17460
rect 54990 17380 55610 17460
rect 55690 17380 55700 17460
rect 49310 17370 55700 17380
rect 55600 16770 55700 17370
rect 48780 16760 55700 16770
rect 48780 16680 48790 16760
rect 48870 16680 49320 16760
rect 49400 16680 50010 16760
rect 50090 16680 50710 16760
rect 50790 16680 51410 16760
rect 51490 16680 52110 16760
rect 52190 16680 52810 16760
rect 52890 16680 53510 16760
rect 53590 16680 54210 16760
rect 54290 16680 54910 16760
rect 54990 16680 55610 16760
rect 55690 16680 55700 16760
rect 48780 16670 55700 16680
rect 49310 16060 55700 16070
rect 49310 15980 49320 16060
rect 49400 15980 50010 16060
rect 50090 15980 50710 16060
rect 50790 15980 51410 16060
rect 51490 15980 52110 16060
rect 52190 15980 52810 16060
rect 52890 15980 53510 16060
rect 53590 15980 54210 16060
rect 54290 15980 54910 16060
rect 54990 15980 55610 16060
rect 55690 15980 55700 16060
rect 49310 15970 55700 15980
rect 55600 15370 55700 15970
rect 48780 15360 55700 15370
rect 48780 15280 48790 15360
rect 48870 15280 49320 15360
rect 49400 15280 50010 15360
rect 50090 15280 50710 15360
rect 50790 15280 51410 15360
rect 51490 15280 52110 15360
rect 52190 15280 52810 15360
rect 52890 15280 53510 15360
rect 53590 15280 54210 15360
rect 54290 15280 54910 15360
rect 54990 15280 55610 15360
rect 55690 15280 55700 15360
rect 48780 15270 55700 15280
<< labels >>
flabel metal2 43290 9290 43290 9290 5 FreeSans 1600 0 0 -800 PFET_GATE
<< end >>
