magic
tech sky130A
magscale 1 2
timestamp 1757109784
<< nwell >>
rect 19300 11490 22740 12800
rect 22997 11427 23989 13767
rect 22997 9057 23989 11167
<< nmos >>
rect 19540 10960 19570 11060
rect 19670 10960 19700 11060
rect 19800 10960 19830 11060
rect 19930 10960 19960 11060
rect 20060 10960 20090 11060
rect 20190 10960 20220 11060
rect 20680 10960 20710 11060
rect 20810 10960 20840 11060
rect 20940 10960 20970 11060
rect 21070 10960 21100 11060
rect 21200 10960 21230 11060
rect 21330 10960 21360 11060
rect 21820 10960 21850 11060
rect 21950 10960 21980 11060
rect 22080 10960 22110 11060
rect 22210 10960 22240 11060
rect 22340 10960 22370 11060
rect 22470 10960 22500 11060
rect 19490 10270 19590 10520
rect 19690 10270 19790 10520
rect 19890 10270 19990 10520
rect 20090 10270 20190 10520
rect 20290 10270 20390 10520
rect 20490 10270 20590 10520
rect 20690 10270 20790 10520
rect 20890 10270 20990 10520
rect 21090 10270 21190 10520
rect 21290 10270 21390 10520
<< pmos >>
rect 19610 12190 19710 12690
rect 19810 12190 19910 12690
rect 20010 12190 20110 12690
rect 20210 12190 20310 12690
rect 20410 12190 20510 12690
rect 20610 12190 20710 12690
rect 20810 12190 20910 12690
rect 21010 12190 21110 12690
rect 21210 12190 21310 12690
rect 21410 12190 21510 12690
rect 19540 11540 19570 11740
rect 19670 11540 19700 11740
rect 19800 11540 19830 11740
rect 19930 11540 19960 11740
rect 20060 11540 20090 11740
rect 20190 11540 20220 11740
rect 20680 11540 20710 11740
rect 20810 11540 20840 11740
rect 20940 11540 20970 11740
rect 21070 11540 21100 11740
rect 21200 11540 21230 11740
rect 21330 11540 21360 11740
rect 21820 11540 21850 11740
rect 21950 11540 21980 11740
rect 22080 11540 22110 11740
rect 22210 11540 22240 11740
rect 22340 11540 22370 11740
rect 22470 11540 22500 11740
<< ndiff >>
rect 19440 11030 19540 11060
rect 19440 10990 19470 11030
rect 19510 10990 19540 11030
rect 19440 10960 19540 10990
rect 19570 11030 19670 11060
rect 19570 10990 19600 11030
rect 19640 10990 19670 11030
rect 19570 10960 19670 10990
rect 19700 11030 19800 11060
rect 19700 10990 19730 11030
rect 19770 10990 19800 11030
rect 19700 10960 19800 10990
rect 19830 11030 19930 11060
rect 19830 10990 19860 11030
rect 19900 10990 19930 11030
rect 19830 10960 19930 10990
rect 19960 11030 20060 11060
rect 19960 10990 19990 11030
rect 20030 10990 20060 11030
rect 19960 10960 20060 10990
rect 20090 11030 20190 11060
rect 20090 10990 20120 11030
rect 20160 10990 20190 11030
rect 20090 10960 20190 10990
rect 20220 11030 20320 11060
rect 20220 10990 20250 11030
rect 20290 10990 20320 11030
rect 20220 10960 20320 10990
rect 20580 11030 20680 11060
rect 20580 10990 20610 11030
rect 20650 10990 20680 11030
rect 20580 10960 20680 10990
rect 20710 11030 20810 11060
rect 20710 10990 20740 11030
rect 20780 10990 20810 11030
rect 20710 10960 20810 10990
rect 20840 11030 20940 11060
rect 20840 10990 20870 11030
rect 20910 10990 20940 11030
rect 20840 10960 20940 10990
rect 20970 11030 21070 11060
rect 20970 10990 21000 11030
rect 21040 10990 21070 11030
rect 20970 10960 21070 10990
rect 21100 11030 21200 11060
rect 21100 10990 21130 11030
rect 21170 10990 21200 11030
rect 21100 10960 21200 10990
rect 21230 11030 21330 11060
rect 21230 10990 21260 11030
rect 21300 10990 21330 11030
rect 21230 10960 21330 10990
rect 21360 11030 21460 11060
rect 21360 10990 21390 11030
rect 21430 10990 21460 11030
rect 21360 10960 21460 10990
rect 21720 11030 21820 11060
rect 21720 10990 21750 11030
rect 21790 10990 21820 11030
rect 21720 10960 21820 10990
rect 21850 11030 21950 11060
rect 21850 10990 21880 11030
rect 21920 10990 21950 11030
rect 21850 10960 21950 10990
rect 21980 11030 22080 11060
rect 21980 10990 22010 11030
rect 22050 10990 22080 11030
rect 21980 10960 22080 10990
rect 22110 11030 22210 11060
rect 22110 10990 22140 11030
rect 22180 10990 22210 11030
rect 22110 10960 22210 10990
rect 22240 11030 22340 11060
rect 22240 10990 22270 11030
rect 22310 10990 22340 11030
rect 22240 10960 22340 10990
rect 22370 11030 22470 11060
rect 22370 10990 22400 11030
rect 22440 10990 22470 11030
rect 22370 10960 22470 10990
rect 22500 11030 22600 11060
rect 22500 10990 22530 11030
rect 22570 10990 22600 11030
rect 22500 10960 22600 10990
rect 19390 10490 19490 10520
rect 19390 10440 19420 10490
rect 19460 10440 19490 10490
rect 19390 10350 19490 10440
rect 19390 10300 19420 10350
rect 19460 10300 19490 10350
rect 19390 10270 19490 10300
rect 19590 10490 19690 10520
rect 19590 10440 19620 10490
rect 19660 10440 19690 10490
rect 19590 10350 19690 10440
rect 19590 10300 19620 10350
rect 19660 10300 19690 10350
rect 19590 10270 19690 10300
rect 19790 10490 19890 10520
rect 19790 10440 19820 10490
rect 19860 10440 19890 10490
rect 19790 10350 19890 10440
rect 19790 10300 19820 10350
rect 19860 10300 19890 10350
rect 19790 10270 19890 10300
rect 19990 10490 20090 10520
rect 19990 10440 20020 10490
rect 20060 10440 20090 10490
rect 19990 10350 20090 10440
rect 19990 10300 20020 10350
rect 20060 10300 20090 10350
rect 19990 10270 20090 10300
rect 20190 10490 20290 10520
rect 20190 10440 20220 10490
rect 20260 10440 20290 10490
rect 20190 10350 20290 10440
rect 20190 10300 20220 10350
rect 20260 10300 20290 10350
rect 20190 10270 20290 10300
rect 20390 10490 20490 10520
rect 20390 10440 20420 10490
rect 20460 10440 20490 10490
rect 20390 10350 20490 10440
rect 20390 10300 20420 10350
rect 20460 10300 20490 10350
rect 20390 10270 20490 10300
rect 20590 10490 20690 10520
rect 20590 10440 20620 10490
rect 20660 10440 20690 10490
rect 20590 10350 20690 10440
rect 20590 10300 20620 10350
rect 20660 10300 20690 10350
rect 20590 10270 20690 10300
rect 20790 10490 20890 10520
rect 20790 10440 20820 10490
rect 20860 10440 20890 10490
rect 20790 10350 20890 10440
rect 20790 10300 20820 10350
rect 20860 10300 20890 10350
rect 20790 10270 20890 10300
rect 20990 10490 21090 10520
rect 20990 10440 21020 10490
rect 21060 10440 21090 10490
rect 20990 10350 21090 10440
rect 20990 10300 21020 10350
rect 21060 10300 21090 10350
rect 20990 10270 21090 10300
rect 21190 10490 21290 10520
rect 21190 10440 21220 10490
rect 21260 10440 21290 10490
rect 21190 10350 21290 10440
rect 21190 10300 21220 10350
rect 21260 10300 21290 10350
rect 21190 10270 21290 10300
rect 21390 10490 21490 10520
rect 21390 10440 21420 10490
rect 21460 10440 21490 10490
rect 21390 10350 21490 10440
rect 21390 10300 21420 10350
rect 21460 10300 21490 10350
rect 21390 10270 21490 10300
<< pdiff >>
rect 19510 12660 19610 12690
rect 19510 12620 19540 12660
rect 19580 12620 19610 12660
rect 19510 12560 19610 12620
rect 19510 12520 19540 12560
rect 19580 12520 19610 12560
rect 19510 12460 19610 12520
rect 19510 12420 19540 12460
rect 19580 12420 19610 12460
rect 19510 12360 19610 12420
rect 19510 12320 19540 12360
rect 19580 12320 19610 12360
rect 19510 12260 19610 12320
rect 19510 12220 19540 12260
rect 19580 12220 19610 12260
rect 19510 12190 19610 12220
rect 19710 12660 19810 12690
rect 19710 12620 19740 12660
rect 19780 12620 19810 12660
rect 19710 12560 19810 12620
rect 19710 12520 19740 12560
rect 19780 12520 19810 12560
rect 19710 12460 19810 12520
rect 19710 12420 19740 12460
rect 19780 12420 19810 12460
rect 19710 12360 19810 12420
rect 19710 12320 19740 12360
rect 19780 12320 19810 12360
rect 19710 12260 19810 12320
rect 19710 12220 19740 12260
rect 19780 12220 19810 12260
rect 19710 12190 19810 12220
rect 19910 12660 20010 12690
rect 19910 12620 19940 12660
rect 19980 12620 20010 12660
rect 19910 12560 20010 12620
rect 19910 12520 19940 12560
rect 19980 12520 20010 12560
rect 19910 12460 20010 12520
rect 19910 12420 19940 12460
rect 19980 12420 20010 12460
rect 19910 12360 20010 12420
rect 19910 12320 19940 12360
rect 19980 12320 20010 12360
rect 19910 12260 20010 12320
rect 19910 12220 19940 12260
rect 19980 12220 20010 12260
rect 19910 12190 20010 12220
rect 20110 12660 20210 12690
rect 20110 12620 20140 12660
rect 20180 12620 20210 12660
rect 20110 12560 20210 12620
rect 20110 12520 20140 12560
rect 20180 12520 20210 12560
rect 20110 12460 20210 12520
rect 20110 12420 20140 12460
rect 20180 12420 20210 12460
rect 20110 12360 20210 12420
rect 20110 12320 20140 12360
rect 20180 12320 20210 12360
rect 20110 12260 20210 12320
rect 20110 12220 20140 12260
rect 20180 12220 20210 12260
rect 20110 12190 20210 12220
rect 20310 12660 20410 12690
rect 20310 12620 20340 12660
rect 20380 12620 20410 12660
rect 20310 12560 20410 12620
rect 20310 12520 20340 12560
rect 20380 12520 20410 12560
rect 20310 12460 20410 12520
rect 20310 12420 20340 12460
rect 20380 12420 20410 12460
rect 20310 12360 20410 12420
rect 20310 12320 20340 12360
rect 20380 12320 20410 12360
rect 20310 12260 20410 12320
rect 20310 12220 20340 12260
rect 20380 12220 20410 12260
rect 20310 12190 20410 12220
rect 20510 12660 20610 12690
rect 20510 12620 20540 12660
rect 20580 12620 20610 12660
rect 20510 12560 20610 12620
rect 20510 12520 20540 12560
rect 20580 12520 20610 12560
rect 20510 12460 20610 12520
rect 20510 12420 20540 12460
rect 20580 12420 20610 12460
rect 20510 12360 20610 12420
rect 20510 12320 20540 12360
rect 20580 12320 20610 12360
rect 20510 12260 20610 12320
rect 20510 12220 20540 12260
rect 20580 12220 20610 12260
rect 20510 12190 20610 12220
rect 20710 12660 20810 12690
rect 20710 12620 20740 12660
rect 20780 12620 20810 12660
rect 20710 12560 20810 12620
rect 20710 12520 20740 12560
rect 20780 12520 20810 12560
rect 20710 12460 20810 12520
rect 20710 12420 20740 12460
rect 20780 12420 20810 12460
rect 20710 12360 20810 12420
rect 20710 12320 20740 12360
rect 20780 12320 20810 12360
rect 20710 12260 20810 12320
rect 20710 12220 20740 12260
rect 20780 12220 20810 12260
rect 20710 12190 20810 12220
rect 20910 12660 21010 12690
rect 20910 12620 20940 12660
rect 20980 12620 21010 12660
rect 20910 12560 21010 12620
rect 20910 12520 20940 12560
rect 20980 12520 21010 12560
rect 20910 12460 21010 12520
rect 20910 12420 20940 12460
rect 20980 12420 21010 12460
rect 20910 12360 21010 12420
rect 20910 12320 20940 12360
rect 20980 12320 21010 12360
rect 20910 12260 21010 12320
rect 20910 12220 20940 12260
rect 20980 12220 21010 12260
rect 20910 12190 21010 12220
rect 21110 12660 21210 12690
rect 21110 12620 21140 12660
rect 21180 12620 21210 12660
rect 21110 12560 21210 12620
rect 21110 12520 21140 12560
rect 21180 12520 21210 12560
rect 21110 12460 21210 12520
rect 21110 12420 21140 12460
rect 21180 12420 21210 12460
rect 21110 12360 21210 12420
rect 21110 12320 21140 12360
rect 21180 12320 21210 12360
rect 21110 12260 21210 12320
rect 21110 12220 21140 12260
rect 21180 12220 21210 12260
rect 21110 12190 21210 12220
rect 21310 12660 21410 12690
rect 21310 12620 21340 12660
rect 21380 12620 21410 12660
rect 21310 12560 21410 12620
rect 21310 12520 21340 12560
rect 21380 12520 21410 12560
rect 21310 12460 21410 12520
rect 21310 12420 21340 12460
rect 21380 12420 21410 12460
rect 21310 12360 21410 12420
rect 21310 12320 21340 12360
rect 21380 12320 21410 12360
rect 21310 12260 21410 12320
rect 21310 12220 21340 12260
rect 21380 12220 21410 12260
rect 21310 12190 21410 12220
rect 21510 12660 21610 12690
rect 21510 12620 21540 12660
rect 21580 12620 21610 12660
rect 21510 12560 21610 12620
rect 21510 12520 21540 12560
rect 21580 12520 21610 12560
rect 21510 12460 21610 12520
rect 21510 12420 21540 12460
rect 21580 12420 21610 12460
rect 21510 12360 21610 12420
rect 21510 12320 21540 12360
rect 21580 12320 21610 12360
rect 21510 12260 21610 12320
rect 21510 12220 21540 12260
rect 21580 12220 21610 12260
rect 21510 12190 21610 12220
rect 19440 11710 19540 11740
rect 19440 11670 19470 11710
rect 19510 11670 19540 11710
rect 19440 11610 19540 11670
rect 19440 11570 19470 11610
rect 19510 11570 19540 11610
rect 19440 11540 19540 11570
rect 19570 11710 19670 11740
rect 19570 11670 19600 11710
rect 19640 11670 19670 11710
rect 19570 11610 19670 11670
rect 19570 11570 19600 11610
rect 19640 11570 19670 11610
rect 19570 11540 19670 11570
rect 19700 11710 19800 11740
rect 19700 11670 19730 11710
rect 19770 11670 19800 11710
rect 19700 11610 19800 11670
rect 19700 11570 19730 11610
rect 19770 11570 19800 11610
rect 19700 11540 19800 11570
rect 19830 11710 19930 11740
rect 19830 11670 19860 11710
rect 19900 11670 19930 11710
rect 19830 11610 19930 11670
rect 19830 11570 19860 11610
rect 19900 11570 19930 11610
rect 19830 11540 19930 11570
rect 19960 11710 20060 11740
rect 19960 11670 19990 11710
rect 20030 11670 20060 11710
rect 19960 11610 20060 11670
rect 19960 11570 19990 11610
rect 20030 11570 20060 11610
rect 19960 11540 20060 11570
rect 20090 11710 20190 11740
rect 20090 11670 20120 11710
rect 20160 11670 20190 11710
rect 20090 11610 20190 11670
rect 20090 11570 20120 11610
rect 20160 11570 20190 11610
rect 20090 11540 20190 11570
rect 20220 11710 20320 11740
rect 20220 11670 20250 11710
rect 20290 11670 20320 11710
rect 20220 11610 20320 11670
rect 20220 11570 20250 11610
rect 20290 11570 20320 11610
rect 20220 11540 20320 11570
rect 20580 11710 20680 11740
rect 20580 11670 20610 11710
rect 20650 11670 20680 11710
rect 20580 11610 20680 11670
rect 20580 11570 20610 11610
rect 20650 11570 20680 11610
rect 20580 11540 20680 11570
rect 20710 11710 20810 11740
rect 20710 11670 20740 11710
rect 20780 11670 20810 11710
rect 20710 11610 20810 11670
rect 20710 11570 20740 11610
rect 20780 11570 20810 11610
rect 20710 11540 20810 11570
rect 20840 11710 20940 11740
rect 20840 11670 20870 11710
rect 20910 11670 20940 11710
rect 20840 11610 20940 11670
rect 20840 11570 20870 11610
rect 20910 11570 20940 11610
rect 20840 11540 20940 11570
rect 20970 11710 21070 11740
rect 20970 11670 21000 11710
rect 21040 11670 21070 11710
rect 20970 11610 21070 11670
rect 20970 11570 21000 11610
rect 21040 11570 21070 11610
rect 20970 11540 21070 11570
rect 21100 11710 21200 11740
rect 21100 11670 21130 11710
rect 21170 11670 21200 11710
rect 21100 11610 21200 11670
rect 21100 11570 21130 11610
rect 21170 11570 21200 11610
rect 21100 11540 21200 11570
rect 21230 11710 21330 11740
rect 21230 11670 21260 11710
rect 21300 11670 21330 11710
rect 21230 11610 21330 11670
rect 21230 11570 21260 11610
rect 21300 11570 21330 11610
rect 21230 11540 21330 11570
rect 21360 11710 21460 11740
rect 21360 11670 21390 11710
rect 21430 11670 21460 11710
rect 21360 11610 21460 11670
rect 21360 11570 21390 11610
rect 21430 11570 21460 11610
rect 21360 11540 21460 11570
rect 21720 11710 21820 11740
rect 21720 11670 21750 11710
rect 21790 11670 21820 11710
rect 21720 11610 21820 11670
rect 21720 11570 21750 11610
rect 21790 11570 21820 11610
rect 21720 11540 21820 11570
rect 21850 11710 21950 11740
rect 21850 11670 21880 11710
rect 21920 11670 21950 11710
rect 21850 11610 21950 11670
rect 21850 11570 21880 11610
rect 21920 11570 21950 11610
rect 21850 11540 21950 11570
rect 21980 11710 22080 11740
rect 21980 11670 22010 11710
rect 22050 11670 22080 11710
rect 21980 11610 22080 11670
rect 21980 11570 22010 11610
rect 22050 11570 22080 11610
rect 21980 11540 22080 11570
rect 22110 11710 22210 11740
rect 22110 11670 22140 11710
rect 22180 11670 22210 11710
rect 22110 11610 22210 11670
rect 22110 11570 22140 11610
rect 22180 11570 22210 11610
rect 22110 11540 22210 11570
rect 22240 11710 22340 11740
rect 22240 11670 22270 11710
rect 22310 11670 22340 11710
rect 22240 11610 22340 11670
rect 22240 11570 22270 11610
rect 22310 11570 22340 11610
rect 22240 11540 22340 11570
rect 22370 11710 22470 11740
rect 22370 11670 22400 11710
rect 22440 11670 22470 11710
rect 22370 11610 22470 11670
rect 22370 11570 22400 11610
rect 22440 11570 22470 11610
rect 22370 11540 22470 11570
rect 22500 11710 22600 11740
rect 22500 11670 22530 11710
rect 22570 11670 22600 11710
rect 22500 11610 22600 11670
rect 22500 11570 22530 11610
rect 22570 11570 22600 11610
rect 22500 11540 22600 11570
<< ndiffc >>
rect 19470 10990 19510 11030
rect 19600 10990 19640 11030
rect 19730 10990 19770 11030
rect 19860 10990 19900 11030
rect 19990 10990 20030 11030
rect 20120 10990 20160 11030
rect 20250 10990 20290 11030
rect 20610 10990 20650 11030
rect 20740 10990 20780 11030
rect 20870 10990 20910 11030
rect 21000 10990 21040 11030
rect 21130 10990 21170 11030
rect 21260 10990 21300 11030
rect 21390 10990 21430 11030
rect 21750 10990 21790 11030
rect 21880 10990 21920 11030
rect 22010 10990 22050 11030
rect 22140 10990 22180 11030
rect 22270 10990 22310 11030
rect 22400 10990 22440 11030
rect 22530 10990 22570 11030
rect 19420 10440 19460 10490
rect 19420 10300 19460 10350
rect 19620 10440 19660 10490
rect 19620 10300 19660 10350
rect 19820 10440 19860 10490
rect 19820 10300 19860 10350
rect 20020 10440 20060 10490
rect 20020 10300 20060 10350
rect 20220 10440 20260 10490
rect 20220 10300 20260 10350
rect 20420 10440 20460 10490
rect 20420 10300 20460 10350
rect 20620 10440 20660 10490
rect 20620 10300 20660 10350
rect 20820 10440 20860 10490
rect 20820 10300 20860 10350
rect 21020 10440 21060 10490
rect 21020 10300 21060 10350
rect 21220 10440 21260 10490
rect 21220 10300 21260 10350
rect 21420 10440 21460 10490
rect 21420 10300 21460 10350
<< pdiffc >>
rect 19540 12620 19580 12660
rect 19540 12520 19580 12560
rect 19540 12420 19580 12460
rect 19540 12320 19580 12360
rect 19540 12220 19580 12260
rect 19740 12620 19780 12660
rect 19740 12520 19780 12560
rect 19740 12420 19780 12460
rect 19740 12320 19780 12360
rect 19740 12220 19780 12260
rect 19940 12620 19980 12660
rect 19940 12520 19980 12560
rect 19940 12420 19980 12460
rect 19940 12320 19980 12360
rect 19940 12220 19980 12260
rect 20140 12620 20180 12660
rect 20140 12520 20180 12560
rect 20140 12420 20180 12460
rect 20140 12320 20180 12360
rect 20140 12220 20180 12260
rect 20340 12620 20380 12660
rect 20340 12520 20380 12560
rect 20340 12420 20380 12460
rect 20340 12320 20380 12360
rect 20340 12220 20380 12260
rect 20540 12620 20580 12660
rect 20540 12520 20580 12560
rect 20540 12420 20580 12460
rect 20540 12320 20580 12360
rect 20540 12220 20580 12260
rect 20740 12620 20780 12660
rect 20740 12520 20780 12560
rect 20740 12420 20780 12460
rect 20740 12320 20780 12360
rect 20740 12220 20780 12260
rect 20940 12620 20980 12660
rect 20940 12520 20980 12560
rect 20940 12420 20980 12460
rect 20940 12320 20980 12360
rect 20940 12220 20980 12260
rect 21140 12620 21180 12660
rect 21140 12520 21180 12560
rect 21140 12420 21180 12460
rect 21140 12320 21180 12360
rect 21140 12220 21180 12260
rect 21340 12620 21380 12660
rect 21340 12520 21380 12560
rect 21340 12420 21380 12460
rect 21340 12320 21380 12360
rect 21340 12220 21380 12260
rect 21540 12620 21580 12660
rect 21540 12520 21580 12560
rect 21540 12420 21580 12460
rect 21540 12320 21580 12360
rect 21540 12220 21580 12260
rect 19470 11670 19510 11710
rect 19470 11570 19510 11610
rect 19600 11670 19640 11710
rect 19600 11570 19640 11610
rect 19730 11670 19770 11710
rect 19730 11570 19770 11610
rect 19860 11670 19900 11710
rect 19860 11570 19900 11610
rect 19990 11670 20030 11710
rect 19990 11570 20030 11610
rect 20120 11670 20160 11710
rect 20120 11570 20160 11610
rect 20250 11670 20290 11710
rect 20250 11570 20290 11610
rect 20610 11670 20650 11710
rect 20610 11570 20650 11610
rect 20740 11670 20780 11710
rect 20740 11570 20780 11610
rect 20870 11670 20910 11710
rect 20870 11570 20910 11610
rect 21000 11670 21040 11710
rect 21000 11570 21040 11610
rect 21130 11670 21170 11710
rect 21130 11570 21170 11610
rect 21260 11670 21300 11710
rect 21260 11570 21300 11610
rect 21390 11670 21430 11710
rect 21390 11570 21430 11610
rect 21750 11670 21790 11710
rect 21750 11570 21790 11610
rect 21880 11670 21920 11710
rect 21880 11570 21920 11610
rect 22010 11670 22050 11710
rect 22010 11570 22050 11610
rect 22140 11670 22180 11710
rect 22140 11570 22180 11610
rect 22270 11670 22310 11710
rect 22270 11570 22310 11610
rect 22400 11670 22440 11710
rect 22400 11570 22440 11610
rect 22530 11670 22570 11710
rect 22530 11570 22570 11610
<< psubdiff >>
rect 19340 11030 19440 11060
rect 19340 10990 19370 11030
rect 19410 10990 19440 11030
rect 19340 10960 19440 10990
rect 20320 11030 20420 11060
rect 20320 10990 20350 11030
rect 20390 10990 20420 11030
rect 20320 10960 20420 10990
rect 21620 11030 21720 11060
rect 21620 10990 21650 11030
rect 21690 10990 21720 11030
rect 21620 10960 21720 10990
rect 22600 11030 22700 11060
rect 22600 10990 22630 11030
rect 22670 10990 22700 11030
rect 22600 10960 22700 10990
rect 19290 10490 19390 10520
rect 19290 10440 19320 10490
rect 19360 10440 19390 10490
rect 19290 10350 19390 10440
rect 19290 10300 19320 10350
rect 19360 10300 19390 10350
rect 19290 10270 19390 10300
rect 21490 10490 21590 10520
rect 21490 10440 21520 10490
rect 21560 10440 21590 10490
rect 21490 10350 21590 10440
rect 21490 10300 21520 10350
rect 21560 10300 21590 10350
rect 21490 10270 21590 10300
<< nsubdiff >>
rect 23033 13697 23129 13731
rect 23857 13697 23953 13731
rect 23033 13635 23067 13697
rect 19410 12660 19510 12690
rect 19410 12620 19440 12660
rect 19480 12620 19510 12660
rect 19410 12560 19510 12620
rect 19410 12520 19440 12560
rect 19480 12520 19510 12560
rect 19410 12460 19510 12520
rect 19410 12420 19440 12460
rect 19480 12420 19510 12460
rect 19410 12360 19510 12420
rect 19410 12320 19440 12360
rect 19480 12320 19510 12360
rect 19410 12260 19510 12320
rect 19410 12220 19440 12260
rect 19480 12220 19510 12260
rect 19410 12190 19510 12220
rect 21610 12660 21710 12690
rect 21610 12620 21640 12660
rect 21680 12620 21710 12660
rect 21610 12560 21710 12620
rect 21610 12520 21640 12560
rect 21680 12520 21710 12560
rect 21610 12460 21710 12520
rect 21610 12420 21640 12460
rect 21680 12420 21710 12460
rect 21610 12360 21710 12420
rect 21610 12320 21640 12360
rect 21680 12320 21710 12360
rect 21610 12260 21710 12320
rect 21610 12220 21640 12260
rect 21680 12220 21710 12260
rect 21610 12190 21710 12220
rect 20480 11710 20580 11740
rect 20480 11670 20510 11710
rect 20550 11670 20580 11710
rect 20480 11610 20580 11670
rect 20480 11570 20510 11610
rect 20550 11570 20580 11610
rect 20480 11540 20580 11570
rect 21460 11710 21560 11740
rect 21460 11670 21490 11710
rect 21530 11670 21560 11710
rect 21460 11610 21560 11670
rect 21460 11570 21490 11610
rect 21530 11570 21560 11610
rect 21460 11540 21560 11570
rect 21620 11710 21720 11740
rect 21620 11670 21650 11710
rect 21690 11670 21720 11710
rect 21620 11610 21720 11670
rect 21620 11570 21650 11610
rect 21690 11570 21720 11610
rect 21620 11540 21720 11570
rect 22600 11710 22700 11740
rect 22600 11670 22630 11710
rect 22670 11670 22700 11710
rect 22600 11610 22700 11670
rect 22600 11570 22630 11610
rect 22670 11570 22700 11610
rect 22600 11540 22700 11570
rect 23919 13635 23953 13697
rect 23033 11497 23067 11559
rect 23919 11497 23953 11559
rect 23033 11463 23129 11497
rect 23857 11463 23953 11497
rect 23033 11097 23129 11131
rect 23857 11097 23953 11131
rect 23033 11035 23067 11097
rect 23919 11035 23953 11097
rect 23033 9127 23067 9189
rect 23919 9127 23953 9189
rect 23033 9093 23129 9127
rect 23857 9093 23953 9127
<< psubdiffcont >>
rect 19370 10990 19410 11030
rect 20350 10990 20390 11030
rect 21650 10990 21690 11030
rect 22630 10990 22670 11030
rect 19320 10440 19360 10490
rect 19320 10300 19360 10350
rect 21520 10440 21560 10490
rect 21520 10300 21560 10350
<< nsubdiffcont >>
rect 23129 13697 23857 13731
rect 19440 12620 19480 12660
rect 19440 12520 19480 12560
rect 19440 12420 19480 12460
rect 19440 12320 19480 12360
rect 19440 12220 19480 12260
rect 21640 12620 21680 12660
rect 21640 12520 21680 12560
rect 21640 12420 21680 12460
rect 21640 12320 21680 12360
rect 21640 12220 21680 12260
rect 20510 11670 20550 11710
rect 20510 11570 20550 11610
rect 21490 11670 21530 11710
rect 21490 11570 21530 11610
rect 21650 11670 21690 11710
rect 21650 11570 21690 11610
rect 22630 11670 22670 11710
rect 22630 11570 22670 11610
rect 23033 11559 23067 13635
rect 23919 11559 23953 13635
rect 23129 11463 23857 11497
rect 23129 11097 23857 11131
rect 23033 9189 23067 11035
rect 23919 9189 23953 11035
rect 23129 9093 23857 9127
<< poly >>
rect 20320 12780 20400 12800
rect 20320 12740 20340 12780
rect 20380 12740 20400 12780
rect 20720 12780 20800 12800
rect 20720 12740 20740 12780
rect 20780 12740 20800 12780
rect 19610 12690 19710 12720
rect 19810 12710 21310 12740
rect 19810 12690 19910 12710
rect 20010 12690 20110 12710
rect 20210 12690 20310 12710
rect 20410 12690 20510 12710
rect 20610 12690 20710 12710
rect 20810 12690 20910 12710
rect 21010 12690 21110 12710
rect 21210 12690 21310 12710
rect 21410 12690 21510 12720
rect 19610 12160 19710 12190
rect 19810 12160 19910 12190
rect 20010 12160 20110 12190
rect 20210 12160 20310 12190
rect 20410 12160 20510 12190
rect 20610 12160 20710 12190
rect 20810 12160 20910 12190
rect 21010 12160 21110 12190
rect 21210 12160 21310 12190
rect 21410 12160 21510 12190
rect 19520 12140 19710 12160
rect 19520 12100 19540 12140
rect 19580 12130 19710 12140
rect 21410 12140 21600 12160
rect 21410 12130 21540 12140
rect 19580 12100 19600 12130
rect 19520 12080 19600 12100
rect 21520 12100 21540 12130
rect 21580 12100 21600 12140
rect 21520 12080 21600 12100
rect 19510 11830 19590 11850
rect 19510 11790 19530 11830
rect 19570 11790 19590 11830
rect 19510 11770 19590 11790
rect 20170 11830 20250 11850
rect 20170 11790 20190 11830
rect 20230 11790 20250 11830
rect 20170 11770 20250 11790
rect 20650 11830 20730 11850
rect 20650 11790 20670 11830
rect 20710 11790 20730 11830
rect 20650 11770 20730 11790
rect 21310 11830 21390 11850
rect 21310 11790 21330 11830
rect 21370 11790 21390 11830
rect 21310 11770 21390 11790
rect 21790 11830 21870 11850
rect 21790 11790 21810 11830
rect 21850 11790 21870 11830
rect 21790 11770 21870 11790
rect 22450 11830 22530 11850
rect 22450 11790 22470 11830
rect 22510 11790 22530 11830
rect 22450 11770 22530 11790
rect 19540 11740 19570 11770
rect 19670 11740 19700 11770
rect 19800 11740 19830 11770
rect 19930 11740 19960 11770
rect 20060 11740 20090 11770
rect 20190 11740 20220 11770
rect 20680 11740 20710 11770
rect 20810 11740 20840 11770
rect 20940 11740 20970 11770
rect 21070 11740 21100 11770
rect 21200 11740 21230 11770
rect 21330 11740 21360 11770
rect 21820 11740 21850 11770
rect 21950 11740 21980 11770
rect 22080 11740 22110 11770
rect 22210 11740 22240 11770
rect 22340 11740 22370 11770
rect 22470 11740 22500 11770
rect 19540 11510 19570 11540
rect 19670 11520 19700 11540
rect 19800 11520 19830 11540
rect 19670 11510 19830 11520
rect 19620 11490 19830 11510
rect 19930 11520 19960 11540
rect 20060 11520 20090 11540
rect 19930 11510 20090 11520
rect 20190 11510 20220 11540
rect 20680 11510 20710 11540
rect 20810 11520 20840 11540
rect 20940 11520 20970 11540
rect 21070 11520 21100 11540
rect 21200 11520 21230 11540
rect 19930 11490 20140 11510
rect 20810 11490 21230 11520
rect 21330 11510 21360 11540
rect 21820 11510 21850 11540
rect 21950 11510 21980 11540
rect 21900 11490 21980 11510
rect 19620 11450 19640 11490
rect 19680 11450 19700 11490
rect 19620 11430 19700 11450
rect 20060 11450 20080 11490
rect 20120 11450 20140 11490
rect 20060 11430 20140 11450
rect 20850 11480 20930 11490
rect 20850 11440 20870 11480
rect 20910 11440 20930 11480
rect 20850 11420 20930 11440
rect 21900 11450 21920 11490
rect 21960 11460 21980 11490
rect 22080 11460 22110 11540
rect 22210 11460 22240 11540
rect 22340 11460 22370 11540
rect 22470 11510 22500 11540
rect 22740 11490 22820 11510
rect 22740 11460 22760 11490
rect 21960 11450 22760 11460
rect 22800 11450 22820 11490
rect 21900 11430 22820 11450
rect 21900 11270 21980 11290
rect 21900 11230 21920 11270
rect 21960 11230 21980 11270
rect 21900 11210 21980 11230
rect 21950 11170 21980 11210
rect 19710 11150 19790 11170
rect 19710 11110 19730 11150
rect 19770 11110 19790 11150
rect 20760 11150 20840 11170
rect 20760 11110 20780 11150
rect 20820 11110 20840 11150
rect 21200 11150 21280 11170
rect 21200 11110 21220 11150
rect 21260 11110 21280 11150
rect 19540 11060 19570 11090
rect 19670 11080 20090 11110
rect 20760 11090 20970 11110
rect 19670 11060 19700 11080
rect 19800 11060 19830 11080
rect 19930 11060 19960 11080
rect 20060 11060 20090 11080
rect 20190 11060 20220 11090
rect 20680 11060 20710 11090
rect 20810 11080 20970 11090
rect 20810 11060 20840 11080
rect 20940 11060 20970 11080
rect 21070 11090 21280 11110
rect 21950 11150 22820 11170
rect 21950 11140 22760 11150
rect 21070 11080 21230 11090
rect 21070 11060 21100 11080
rect 21200 11060 21230 11080
rect 21330 11060 21360 11090
rect 21820 11060 21850 11090
rect 21950 11060 21980 11140
rect 22080 11060 22110 11140
rect 22210 11060 22240 11140
rect 22340 11060 22370 11140
rect 22740 11110 22760 11140
rect 22800 11110 22820 11150
rect 22740 11090 22820 11110
rect 22470 11060 22500 11090
rect 19540 10930 19570 10960
rect 19670 10930 19700 10960
rect 19800 10930 19830 10960
rect 19930 10930 19960 10960
rect 20060 10930 20090 10960
rect 20190 10930 20220 10960
rect 20680 10930 20710 10960
rect 20810 10930 20840 10960
rect 20940 10930 20970 10960
rect 21070 10930 21100 10960
rect 21200 10930 21230 10960
rect 21330 10930 21360 10960
rect 21820 10930 21850 10960
rect 21950 10930 21980 10960
rect 22080 10930 22110 10960
rect 22210 10930 22240 10960
rect 22340 10930 22370 10960
rect 22470 10930 22500 10960
rect 19510 10910 19600 10930
rect 19510 10860 19530 10910
rect 19580 10860 19600 10910
rect 19510 10840 19600 10860
rect 20160 10910 20250 10930
rect 20160 10860 20180 10910
rect 20230 10860 20250 10910
rect 20160 10840 20250 10860
rect 20650 10910 20730 10930
rect 20650 10870 20670 10910
rect 20710 10870 20730 10910
rect 20650 10850 20730 10870
rect 21310 10910 21390 10930
rect 21310 10870 21330 10910
rect 21370 10870 21390 10910
rect 21310 10850 21390 10870
rect 21790 10910 21870 10930
rect 21790 10870 21810 10910
rect 21850 10870 21870 10910
rect 21790 10850 21870 10870
rect 22450 10910 22530 10930
rect 22450 10870 22470 10910
rect 22510 10870 22530 10910
rect 22450 10850 22530 10870
rect 19400 10610 19480 10630
rect 19400 10570 19420 10610
rect 19460 10580 19480 10610
rect 21400 10610 21480 10630
rect 21400 10580 21420 10610
rect 19460 10570 19590 10580
rect 19400 10550 19590 10570
rect 21290 10570 21420 10580
rect 21460 10570 21480 10610
rect 21290 10550 21480 10570
rect 19490 10520 19590 10550
rect 19690 10520 19790 10550
rect 19890 10520 19990 10550
rect 20090 10520 20190 10550
rect 20290 10520 20390 10550
rect 20490 10520 20590 10550
rect 20690 10520 20790 10550
rect 20890 10520 20990 10550
rect 21090 10520 21190 10550
rect 21290 10520 21390 10550
rect 19490 10240 19590 10270
rect 19690 10250 19790 10270
rect 19890 10250 19990 10270
rect 20090 10250 20190 10270
rect 20290 10250 20390 10270
rect 20490 10250 20590 10270
rect 20690 10250 20790 10270
rect 20890 10250 20990 10270
rect 21090 10250 21190 10270
rect 19690 10220 21190 10250
rect 21290 10240 21390 10270
rect 20200 10180 20220 10220
rect 20260 10180 20280 10220
rect 20200 10160 20280 10180
rect 20600 10180 20620 10220
rect 20660 10180 20680 10220
rect 20600 10160 20680 10180
rect 19244 10024 19674 10040
rect 19244 9990 19260 10024
rect 19294 9990 19674 10024
rect 19244 9974 19674 9990
rect 20154 10024 20584 10040
rect 20154 9990 20534 10024
rect 20568 9990 20584 10024
rect 20154 9974 20584 9990
<< polycont >>
rect 20340 12740 20380 12780
rect 20740 12740 20780 12780
rect 19540 12100 19580 12140
rect 21540 12100 21580 12140
rect 19530 11790 19570 11830
rect 20190 11790 20230 11830
rect 20670 11790 20710 11830
rect 21330 11790 21370 11830
rect 21810 11790 21850 11830
rect 22470 11790 22510 11830
rect 19640 11450 19680 11490
rect 20080 11450 20120 11490
rect 20870 11440 20910 11480
rect 21920 11450 21960 11490
rect 22760 11450 22800 11490
rect 21920 11230 21960 11270
rect 19730 11110 19770 11150
rect 20780 11110 20820 11150
rect 21220 11110 21260 11150
rect 22760 11110 22800 11150
rect 19530 10860 19580 10910
rect 20180 10860 20230 10910
rect 20670 10870 20710 10910
rect 21330 10870 21370 10910
rect 21810 10870 21850 10910
rect 22470 10870 22510 10910
rect 19420 10570 19460 10610
rect 21420 10570 21460 10610
rect 20220 10180 20260 10220
rect 20620 10180 20660 10220
rect 19260 9990 19294 10024
rect 20534 9990 20568 10024
<< xpolycontact >>
rect 23658 13160 23796 13592
rect 23190 11602 23328 12034
rect 23190 10560 23328 10992
rect 23658 9232 23796 9664
<< npolyres >>
rect 19674 9974 20154 10040
<< ppolyres >>
rect 23190 12918 23562 13056
rect 23190 12034 23328 12918
rect 23424 12276 23562 12918
rect 23658 12276 23796 13160
rect 23424 12138 23796 12276
rect 23190 9906 23328 10560
rect 23424 10318 23796 10456
rect 23424 9906 23562 10318
rect 23190 9768 23562 9906
rect 23658 9664 23796 10318
<< locali >>
rect 23033 13697 23129 13731
rect 23857 13697 23953 13731
rect 23033 13635 23067 13697
rect 23010 13170 23033 13190
rect 23919 13635 23953 13697
rect 23067 13170 23090 13190
rect 23010 13130 23030 13170
rect 23070 13130 23090 13170
rect 23010 13110 23033 13130
rect 20320 12780 20400 12800
rect 20320 12740 20340 12780
rect 20380 12740 20400 12780
rect 20320 12720 20400 12740
rect 20720 12780 20800 12800
rect 20720 12740 20740 12780
rect 20780 12740 20800 12780
rect 20720 12720 20800 12740
rect 19420 12660 19600 12680
rect 19420 12620 19440 12660
rect 19480 12620 19540 12660
rect 19580 12620 19600 12660
rect 19420 12560 19600 12620
rect 19420 12520 19440 12560
rect 19480 12520 19540 12560
rect 19580 12520 19600 12560
rect 19420 12460 19600 12520
rect 19420 12420 19440 12460
rect 19480 12420 19540 12460
rect 19580 12420 19600 12460
rect 19420 12360 19600 12420
rect 19420 12320 19440 12360
rect 19480 12320 19540 12360
rect 19580 12320 19600 12360
rect 19420 12260 19600 12320
rect 19420 12220 19440 12260
rect 19480 12220 19540 12260
rect 19580 12220 19600 12260
rect 19420 12200 19600 12220
rect 19720 12660 19800 12680
rect 19720 12620 19740 12660
rect 19780 12620 19800 12660
rect 19720 12560 19800 12620
rect 19720 12520 19740 12560
rect 19780 12520 19800 12560
rect 19720 12460 19800 12520
rect 19720 12420 19740 12460
rect 19780 12420 19800 12460
rect 19720 12360 19800 12420
rect 19720 12320 19740 12360
rect 19780 12320 19800 12360
rect 19720 12260 19800 12320
rect 19720 12220 19740 12260
rect 19780 12220 19800 12260
rect 19720 12200 19800 12220
rect 19920 12660 20000 12680
rect 19920 12620 19940 12660
rect 19980 12620 20000 12660
rect 19920 12560 20000 12620
rect 19920 12520 19940 12560
rect 19980 12520 20000 12560
rect 19920 12460 20000 12520
rect 19920 12420 19940 12460
rect 19980 12420 20000 12460
rect 19920 12360 20000 12420
rect 19920 12320 19940 12360
rect 19980 12320 20000 12360
rect 19920 12260 20000 12320
rect 19920 12220 19940 12260
rect 19980 12220 20000 12260
rect 19920 12200 20000 12220
rect 20120 12660 20200 12680
rect 20120 12620 20140 12660
rect 20180 12620 20200 12660
rect 20120 12560 20200 12620
rect 20120 12520 20140 12560
rect 20180 12520 20200 12560
rect 20120 12460 20200 12520
rect 20120 12420 20140 12460
rect 20180 12420 20200 12460
rect 20120 12360 20200 12420
rect 20120 12320 20140 12360
rect 20180 12320 20200 12360
rect 20120 12260 20200 12320
rect 20120 12220 20140 12260
rect 20180 12220 20200 12260
rect 20120 12200 20200 12220
rect 20320 12660 20400 12680
rect 20320 12620 20340 12660
rect 20380 12620 20400 12660
rect 20320 12560 20400 12620
rect 20320 12520 20340 12560
rect 20380 12520 20400 12560
rect 20320 12460 20400 12520
rect 20320 12420 20340 12460
rect 20380 12420 20400 12460
rect 20320 12360 20400 12420
rect 20320 12320 20340 12360
rect 20380 12320 20400 12360
rect 20320 12260 20400 12320
rect 20320 12220 20340 12260
rect 20380 12220 20400 12260
rect 20320 12200 20400 12220
rect 20520 12660 20600 12680
rect 20520 12620 20540 12660
rect 20580 12620 20600 12660
rect 20520 12560 20600 12620
rect 20520 12520 20540 12560
rect 20580 12520 20600 12560
rect 20520 12460 20600 12520
rect 20520 12420 20540 12460
rect 20580 12420 20600 12460
rect 20520 12360 20600 12420
rect 20520 12320 20540 12360
rect 20580 12320 20600 12360
rect 20520 12260 20600 12320
rect 20520 12220 20540 12260
rect 20580 12220 20600 12260
rect 20520 12200 20600 12220
rect 20720 12660 20800 12680
rect 20720 12620 20740 12660
rect 20780 12620 20800 12660
rect 20720 12560 20800 12620
rect 20720 12520 20740 12560
rect 20780 12520 20800 12560
rect 20720 12460 20800 12520
rect 20720 12420 20740 12460
rect 20780 12420 20800 12460
rect 20720 12360 20800 12420
rect 20720 12320 20740 12360
rect 20780 12320 20800 12360
rect 20720 12260 20800 12320
rect 20720 12220 20740 12260
rect 20780 12220 20800 12260
rect 20720 12200 20800 12220
rect 20920 12660 21000 12680
rect 20920 12620 20940 12660
rect 20980 12620 21000 12660
rect 20920 12560 21000 12620
rect 20920 12520 20940 12560
rect 20980 12520 21000 12560
rect 20920 12460 21000 12520
rect 20920 12420 20940 12460
rect 20980 12420 21000 12460
rect 20920 12360 21000 12420
rect 20920 12320 20940 12360
rect 20980 12320 21000 12360
rect 20920 12260 21000 12320
rect 20920 12220 20940 12260
rect 20980 12220 21000 12260
rect 20920 12200 21000 12220
rect 21120 12660 21200 12680
rect 21120 12620 21140 12660
rect 21180 12620 21200 12660
rect 21120 12560 21200 12620
rect 21120 12520 21140 12560
rect 21180 12520 21200 12560
rect 21120 12460 21200 12520
rect 21120 12420 21140 12460
rect 21180 12420 21200 12460
rect 21120 12360 21200 12420
rect 21120 12320 21140 12360
rect 21180 12320 21200 12360
rect 21120 12260 21200 12320
rect 21120 12220 21140 12260
rect 21180 12220 21200 12260
rect 21120 12200 21200 12220
rect 21320 12660 21400 12680
rect 21320 12620 21340 12660
rect 21380 12620 21400 12660
rect 21320 12560 21400 12620
rect 21320 12520 21340 12560
rect 21380 12520 21400 12560
rect 21320 12460 21400 12520
rect 21320 12420 21340 12460
rect 21380 12420 21400 12460
rect 21320 12360 21400 12420
rect 21320 12320 21340 12360
rect 21380 12320 21400 12360
rect 21320 12260 21400 12320
rect 21320 12220 21340 12260
rect 21380 12220 21400 12260
rect 21320 12200 21400 12220
rect 21520 12660 21700 12680
rect 21520 12620 21540 12660
rect 21580 12620 21640 12660
rect 21680 12620 21700 12660
rect 21520 12560 21700 12620
rect 21520 12520 21540 12560
rect 21580 12520 21640 12560
rect 21680 12520 21700 12560
rect 21520 12460 21700 12520
rect 21520 12420 21540 12460
rect 21580 12420 21640 12460
rect 21680 12420 21700 12460
rect 21520 12360 21700 12420
rect 21520 12320 21540 12360
rect 21580 12320 21640 12360
rect 21680 12320 21700 12360
rect 21520 12260 21700 12320
rect 21520 12220 21540 12260
rect 21580 12220 21640 12260
rect 21680 12220 21700 12260
rect 21520 12200 21700 12220
rect 19520 12140 19600 12200
rect 19520 12100 19540 12140
rect 19580 12100 19600 12140
rect 19520 12080 19600 12100
rect 21520 12140 21600 12160
rect 21520 12100 21540 12140
rect 21580 12100 21600 12140
rect 21520 12080 21600 12100
rect 21000 11980 21080 12000
rect 21000 11940 21020 11980
rect 21060 11940 21080 11980
rect 21000 11920 21080 11940
rect 22120 11980 22200 12000
rect 22120 11940 22140 11980
rect 22180 11940 22200 11980
rect 22120 11920 22200 11940
rect 19920 11870 20000 11890
rect 19510 11830 19590 11850
rect 19510 11810 19530 11830
rect 19470 11790 19530 11810
rect 19570 11810 19590 11830
rect 19920 11830 19940 11870
rect 19980 11830 20000 11870
rect 19920 11810 20000 11830
rect 20170 11830 20250 11850
rect 20170 11810 20190 11830
rect 19570 11790 20190 11810
rect 20230 11810 20250 11830
rect 20650 11830 20730 11850
rect 20650 11810 20670 11830
rect 20230 11790 20290 11810
rect 19470 11770 20290 11790
rect 19470 11730 19510 11770
rect 19600 11730 19640 11770
rect 19860 11730 19900 11770
rect 20120 11730 20160 11770
rect 20250 11730 20290 11770
rect 20610 11790 20670 11810
rect 20710 11810 20730 11830
rect 21000 11810 21040 11920
rect 21310 11830 21390 11850
rect 21310 11810 21330 11830
rect 20710 11790 21330 11810
rect 21370 11810 21390 11830
rect 21790 11830 21870 11850
rect 21790 11810 21810 11830
rect 21370 11790 21430 11810
rect 20610 11770 21430 11790
rect 20610 11730 20650 11770
rect 20740 11730 20780 11770
rect 21000 11730 21040 11770
rect 21260 11730 21300 11770
rect 21390 11730 21430 11770
rect 21750 11790 21810 11810
rect 21850 11810 21870 11830
rect 22140 11810 22180 11920
rect 22450 11830 22530 11850
rect 22450 11810 22470 11830
rect 21850 11790 22470 11810
rect 22510 11810 22530 11830
rect 22510 11790 22570 11810
rect 21750 11770 22570 11790
rect 21750 11730 21790 11770
rect 21880 11730 21920 11770
rect 22140 11730 22180 11770
rect 22400 11730 22440 11770
rect 22530 11730 22570 11770
rect 19450 11710 19530 11730
rect 19450 11670 19470 11710
rect 19510 11670 19530 11710
rect 19450 11610 19530 11670
rect 19450 11570 19470 11610
rect 19510 11570 19530 11610
rect 19450 11550 19530 11570
rect 19580 11710 19660 11730
rect 19580 11670 19600 11710
rect 19640 11670 19660 11710
rect 19580 11610 19660 11670
rect 19580 11570 19600 11610
rect 19640 11570 19660 11610
rect 19580 11550 19660 11570
rect 19710 11710 19790 11730
rect 19710 11670 19730 11710
rect 19770 11670 19790 11710
rect 19710 11610 19790 11670
rect 19710 11570 19730 11610
rect 19770 11570 19790 11610
rect 19710 11550 19790 11570
rect 19840 11710 19920 11730
rect 19840 11670 19860 11710
rect 19900 11670 19920 11710
rect 19840 11610 19920 11670
rect 19840 11570 19860 11610
rect 19900 11570 19920 11610
rect 19840 11550 19920 11570
rect 19970 11710 20050 11730
rect 19970 11670 19990 11710
rect 20030 11670 20050 11710
rect 19970 11610 20050 11670
rect 19970 11570 19990 11610
rect 20030 11570 20050 11610
rect 19970 11550 20050 11570
rect 20100 11710 20190 11730
rect 20100 11670 20120 11710
rect 20160 11670 20190 11710
rect 20100 11610 20190 11670
rect 20100 11570 20120 11610
rect 20160 11570 20190 11610
rect 20100 11550 20190 11570
rect 20230 11710 20310 11730
rect 20230 11670 20250 11710
rect 20290 11670 20310 11710
rect 20230 11610 20310 11670
rect 20230 11570 20250 11610
rect 20290 11570 20310 11610
rect 20230 11550 20310 11570
rect 20490 11710 20670 11730
rect 20490 11670 20510 11710
rect 20550 11670 20610 11710
rect 20650 11670 20670 11710
rect 20490 11610 20670 11670
rect 20490 11570 20510 11610
rect 20550 11570 20610 11610
rect 20650 11570 20670 11610
rect 20490 11550 20670 11570
rect 20720 11710 20800 11730
rect 20720 11670 20740 11710
rect 20780 11670 20800 11710
rect 20720 11610 20800 11670
rect 20720 11570 20740 11610
rect 20780 11570 20800 11610
rect 20720 11550 20800 11570
rect 20850 11710 20930 11730
rect 20850 11670 20870 11710
rect 20910 11670 20930 11710
rect 20850 11610 20930 11670
rect 20850 11570 20870 11610
rect 20910 11570 20930 11610
rect 20850 11550 20930 11570
rect 20980 11710 21060 11730
rect 20980 11670 21000 11710
rect 21040 11670 21060 11710
rect 20980 11610 21060 11670
rect 20980 11570 21000 11610
rect 21040 11570 21060 11610
rect 20980 11550 21060 11570
rect 21110 11710 21190 11730
rect 21110 11670 21130 11710
rect 21170 11670 21190 11710
rect 21110 11610 21190 11670
rect 21110 11570 21130 11610
rect 21170 11570 21190 11610
rect 21110 11550 21190 11570
rect 21240 11710 21320 11730
rect 21240 11670 21260 11710
rect 21300 11670 21320 11710
rect 21240 11610 21320 11670
rect 21240 11570 21260 11610
rect 21300 11570 21320 11610
rect 21240 11550 21320 11570
rect 21370 11710 21550 11730
rect 21370 11670 21390 11710
rect 21430 11670 21490 11710
rect 21530 11670 21550 11710
rect 21370 11610 21550 11670
rect 21370 11570 21390 11610
rect 21430 11570 21490 11610
rect 21530 11570 21550 11610
rect 21370 11550 21550 11570
rect 21630 11710 21810 11730
rect 21630 11670 21650 11710
rect 21690 11670 21750 11710
rect 21790 11670 21810 11710
rect 21630 11610 21810 11670
rect 21630 11570 21650 11610
rect 21690 11570 21750 11610
rect 21790 11570 21810 11610
rect 21630 11550 21810 11570
rect 21860 11710 21940 11730
rect 21860 11670 21880 11710
rect 21920 11670 21940 11710
rect 21860 11610 21940 11670
rect 21860 11570 21880 11610
rect 21920 11570 21940 11610
rect 21860 11550 21940 11570
rect 21990 11710 22070 11730
rect 21990 11670 22010 11710
rect 22050 11670 22070 11710
rect 21990 11610 22070 11670
rect 21990 11570 22010 11610
rect 22050 11570 22070 11610
rect 21990 11550 22070 11570
rect 22120 11710 22200 11730
rect 22120 11670 22140 11710
rect 22180 11670 22200 11710
rect 22120 11610 22200 11670
rect 22120 11570 22140 11610
rect 22180 11570 22200 11610
rect 22120 11550 22200 11570
rect 22250 11710 22330 11730
rect 22250 11670 22270 11710
rect 22310 11670 22330 11710
rect 22250 11610 22330 11670
rect 22250 11570 22270 11610
rect 22310 11570 22330 11610
rect 22250 11550 22330 11570
rect 22380 11710 22460 11730
rect 22380 11670 22400 11710
rect 22440 11670 22460 11710
rect 22380 11610 22460 11670
rect 22380 11570 22400 11610
rect 22440 11570 22460 11610
rect 22380 11550 22460 11570
rect 22510 11710 22690 11730
rect 22510 11670 22530 11710
rect 22570 11670 22630 11710
rect 22670 11670 22690 11710
rect 22510 11610 22690 11670
rect 22510 11570 22530 11610
rect 22570 11570 22630 11610
rect 22670 11570 22690 11610
rect 22510 11550 22690 11570
rect 23067 13110 23090 13130
rect 19620 11490 19700 11510
rect 19620 11450 19640 11490
rect 19680 11450 19700 11490
rect 19620 11430 19700 11450
rect 20060 11490 20140 11510
rect 20060 11450 20080 11490
rect 20120 11450 20140 11490
rect 20060 11430 20140 11450
rect 20850 11480 20930 11500
rect 20850 11440 20870 11480
rect 20910 11440 20930 11480
rect 20850 11420 20930 11440
rect 21900 11490 21980 11510
rect 21900 11450 21920 11490
rect 21960 11450 21980 11490
rect 21900 11430 21980 11450
rect 22030 11340 22070 11550
rect 22250 11340 22290 11550
rect 22740 11490 22820 11510
rect 22740 11450 22760 11490
rect 22800 11450 22820 11490
rect 23033 11497 23067 11559
rect 23919 11497 23953 11559
rect 23033 11463 23129 11497
rect 23857 11463 23953 11497
rect 22740 11430 22820 11450
rect 22030 11320 22110 11340
rect 21900 11270 21980 11290
rect 21900 11230 21920 11270
rect 21960 11230 21980 11270
rect 21900 11210 21980 11230
rect 22030 11280 22050 11320
rect 22090 11280 22110 11320
rect 22030 11260 22110 11280
rect 22230 11320 22310 11340
rect 22230 11280 22250 11320
rect 22290 11280 22310 11320
rect 22230 11260 22310 11280
rect 24060 11320 24140 11340
rect 24060 11280 24080 11320
rect 24120 11280 24140 11320
rect 24060 11260 24140 11280
rect 19710 11150 19790 11170
rect 19710 11110 19730 11150
rect 19770 11110 19790 11150
rect 19710 11090 19790 11110
rect 20760 11150 20840 11170
rect 20760 11110 20780 11150
rect 20820 11110 20840 11150
rect 20760 11090 20840 11110
rect 21200 11150 21280 11170
rect 21200 11110 21220 11150
rect 21260 11110 21280 11150
rect 21200 11090 21280 11110
rect 22030 11050 22070 11260
rect 22250 11050 22290 11260
rect 22740 11150 22820 11170
rect 22740 11110 22760 11150
rect 22800 11110 22820 11150
rect 22740 11090 22820 11110
rect 23033 11097 23129 11131
rect 23857 11097 23953 11131
rect 19350 11030 19530 11050
rect 19350 10990 19370 11030
rect 19410 10990 19470 11030
rect 19510 10990 19530 11030
rect 19350 10970 19530 10990
rect 19580 11030 19660 11050
rect 19580 10990 19600 11030
rect 19640 10990 19660 11030
rect 19580 10970 19660 10990
rect 19710 11030 19790 11050
rect 19710 10990 19730 11030
rect 19770 10990 19790 11030
rect 19710 10970 19790 10990
rect 19840 11030 19920 11050
rect 19840 10990 19860 11030
rect 19900 10990 19920 11030
rect 19840 10970 19920 10990
rect 19970 11030 20050 11050
rect 19970 10990 19990 11030
rect 20030 10990 20050 11030
rect 19970 10970 20050 10990
rect 20100 11030 20180 11050
rect 20100 10990 20120 11030
rect 20160 10990 20180 11030
rect 20100 10970 20180 10990
rect 20230 11030 20410 11050
rect 20230 10990 20250 11030
rect 20290 10990 20350 11030
rect 20390 10990 20410 11030
rect 20230 10970 20410 10990
rect 20590 11030 20670 11050
rect 20590 10990 20610 11030
rect 20650 10990 20670 11030
rect 20590 10970 20670 10990
rect 20720 11030 20800 11050
rect 20720 10990 20740 11030
rect 20780 10990 20800 11030
rect 20720 10970 20800 10990
rect 20850 11030 20930 11050
rect 20850 10990 20870 11030
rect 20910 10990 20930 11030
rect 20850 10970 20930 10990
rect 20980 11030 21060 11050
rect 20980 10990 21000 11030
rect 21040 10990 21060 11030
rect 20980 10970 21060 10990
rect 21110 11030 21190 11050
rect 21110 10990 21130 11030
rect 21170 10990 21190 11030
rect 21110 10970 21190 10990
rect 21240 11030 21320 11050
rect 21240 10990 21260 11030
rect 21300 10990 21320 11030
rect 21240 10970 21320 10990
rect 21370 11030 21450 11050
rect 21370 10990 21390 11030
rect 21430 10990 21450 11030
rect 21370 10970 21450 10990
rect 21630 11030 21810 11050
rect 21630 10990 21650 11030
rect 21690 10990 21750 11030
rect 21790 10990 21810 11030
rect 21630 10970 21810 10990
rect 21860 11030 21940 11050
rect 21860 10990 21880 11030
rect 21920 10990 21940 11030
rect 21860 10970 21940 10990
rect 21990 11030 22070 11050
rect 21990 10990 22010 11030
rect 22050 10990 22070 11030
rect 21990 10970 22070 10990
rect 22120 11030 22200 11050
rect 22120 10990 22140 11030
rect 22180 10990 22200 11030
rect 22120 10970 22200 10990
rect 22250 11030 22330 11050
rect 22250 10990 22270 11030
rect 22310 10990 22330 11030
rect 22250 10970 22330 10990
rect 22380 11030 22460 11050
rect 22380 10990 22400 11030
rect 22440 10990 22460 11030
rect 22380 10970 22460 10990
rect 22510 11030 22690 11050
rect 22510 10990 22530 11030
rect 22570 10990 22630 11030
rect 22670 10990 22690 11030
rect 22510 10970 22690 10990
rect 23033 11035 23067 11097
rect 19470 10930 19510 10970
rect 19600 10930 19640 10970
rect 19860 10930 19900 10970
rect 20120 10930 20160 10970
rect 20250 10930 20290 10970
rect 19470 10910 20290 10930
rect 19470 10890 19530 10910
rect 19510 10860 19530 10890
rect 19580 10890 20180 10910
rect 19580 10860 19600 10890
rect 19510 10840 19600 10860
rect 19860 10780 19900 10890
rect 20160 10860 20180 10890
rect 20230 10890 20290 10910
rect 20610 10930 20650 10970
rect 20740 10930 20780 10970
rect 21000 10930 21040 10970
rect 21260 10930 21300 10970
rect 21390 10930 21430 10970
rect 20610 10910 21430 10930
rect 20610 10890 20670 10910
rect 20230 10860 20250 10890
rect 20160 10840 20250 10860
rect 20650 10870 20670 10890
rect 20710 10890 21330 10910
rect 20710 10870 20730 10890
rect 20650 10850 20730 10870
rect 20980 10870 21060 10890
rect 20980 10830 21000 10870
rect 21040 10830 21060 10870
rect 21310 10870 21330 10890
rect 21370 10890 21430 10910
rect 21750 10930 21790 10970
rect 21880 10930 21920 10970
rect 22140 10930 22180 10970
rect 22400 10930 22440 10970
rect 22530 10930 22570 10970
rect 21750 10910 22570 10930
rect 21370 10870 21390 10890
rect 21750 10880 21810 10910
rect 21310 10850 21390 10870
rect 21790 10870 21810 10880
rect 21850 10880 22470 10910
rect 21850 10870 21870 10880
rect 21790 10850 21870 10870
rect 20980 10810 21060 10830
rect 22140 10780 22180 10880
rect 22450 10870 22470 10880
rect 22510 10880 22570 10910
rect 22510 10870 22530 10880
rect 22450 10850 22530 10870
rect 19840 10760 19920 10780
rect 19840 10720 19860 10760
rect 19900 10720 19920 10760
rect 19840 10700 19920 10720
rect 22120 10760 22200 10780
rect 22120 10720 22140 10760
rect 22180 10720 22200 10760
rect 22120 10700 22200 10720
rect 20980 10650 21060 10670
rect 19400 10610 19480 10630
rect 19400 10570 19420 10610
rect 19460 10570 19480 10610
rect 20980 10610 21000 10650
rect 21040 10610 21060 10650
rect 20980 10590 21060 10610
rect 19400 10550 19480 10570
rect 19820 10550 21060 10590
rect 21400 10610 21480 10630
rect 21400 10570 21420 10610
rect 21460 10570 21480 10610
rect 21400 10550 21480 10570
rect 19420 10510 19460 10550
rect 19820 10510 19860 10550
rect 21020 10510 21060 10550
rect 21420 10510 21460 10550
rect 19300 10490 19480 10510
rect 19300 10440 19320 10490
rect 19360 10440 19420 10490
rect 19460 10440 19480 10490
rect 19300 10350 19480 10440
rect 19300 10300 19320 10350
rect 19360 10300 19420 10350
rect 19460 10300 19480 10350
rect 19300 10280 19480 10300
rect 19600 10490 19680 10510
rect 19600 10440 19620 10490
rect 19660 10440 19680 10490
rect 19600 10350 19680 10440
rect 19600 10300 19620 10350
rect 19660 10300 19680 10350
rect 19600 10280 19680 10300
rect 19800 10490 19880 10510
rect 19800 10440 19820 10490
rect 19860 10440 19880 10490
rect 19800 10350 19880 10440
rect 19800 10300 19820 10350
rect 19860 10300 19880 10350
rect 19800 10280 19880 10300
rect 20000 10490 20080 10510
rect 20000 10440 20020 10490
rect 20060 10440 20080 10490
rect 20000 10350 20080 10440
rect 20000 10300 20020 10350
rect 20060 10300 20080 10350
rect 20000 10280 20080 10300
rect 20200 10490 20280 10510
rect 20200 10440 20220 10490
rect 20260 10440 20280 10490
rect 20200 10350 20280 10440
rect 20200 10300 20220 10350
rect 20260 10300 20280 10350
rect 20200 10280 20280 10300
rect 20400 10490 20480 10510
rect 20400 10440 20420 10490
rect 20460 10440 20480 10490
rect 20400 10350 20480 10440
rect 20400 10300 20420 10350
rect 20460 10300 20480 10350
rect 20400 10280 20480 10300
rect 20600 10490 20680 10510
rect 20600 10440 20620 10490
rect 20660 10440 20680 10490
rect 20600 10350 20680 10440
rect 20600 10300 20620 10350
rect 20660 10300 20680 10350
rect 20600 10280 20680 10300
rect 20800 10490 20880 10510
rect 20800 10440 20820 10490
rect 20860 10440 20880 10490
rect 20800 10350 20880 10440
rect 20800 10300 20820 10350
rect 20860 10300 20880 10350
rect 20800 10280 20880 10300
rect 21000 10490 21080 10510
rect 21000 10440 21020 10490
rect 21060 10440 21080 10490
rect 21000 10350 21080 10440
rect 21000 10300 21020 10350
rect 21060 10300 21080 10350
rect 21000 10280 21080 10300
rect 21200 10490 21280 10510
rect 21200 10440 21220 10490
rect 21260 10440 21280 10490
rect 21200 10350 21280 10440
rect 21200 10300 21220 10350
rect 21260 10300 21280 10350
rect 21200 10280 21280 10300
rect 21400 10490 21580 10510
rect 21400 10440 21420 10490
rect 21460 10440 21520 10490
rect 21560 10440 21580 10490
rect 21400 10350 21580 10440
rect 21400 10300 21420 10350
rect 21460 10300 21520 10350
rect 21560 10300 21580 10350
rect 21400 10280 21580 10300
rect 20220 10240 20260 10280
rect 20620 10240 20660 10280
rect 20200 10220 20680 10240
rect 20200 10180 20220 10220
rect 20260 10180 20620 10220
rect 20660 10180 20680 10220
rect 20200 10160 20680 10180
rect 19140 10040 19260 10050
rect 20590 10040 20680 10160
rect 19140 10030 19294 10040
rect 19140 9990 19160 10030
rect 19200 10024 19294 10030
rect 19200 9990 19260 10024
rect 19140 9974 19294 9990
rect 20534 10024 20680 10040
rect 20568 9990 20680 10024
rect 20534 9974 20680 9990
rect 19140 9970 19260 9974
rect 20560 9970 20680 9974
rect 23010 9640 23033 9660
rect 23919 11035 23953 11097
rect 23067 9640 23090 9660
rect 23010 9600 23030 9640
rect 23070 9600 23090 9640
rect 23010 9580 23033 9600
rect 23067 9580 23090 9600
rect 23033 9127 23067 9189
rect 23680 9130 23780 9150
rect 23680 9127 23700 9130
rect 23760 9127 23780 9130
rect 23919 9127 23953 9189
rect 23033 9093 23129 9127
rect 23857 9093 23953 9127
rect 23680 9070 23700 9093
rect 23760 9070 23780 9093
rect 23680 9050 23780 9070
<< viali >>
rect 23700 13450 23760 13510
rect 23690 13200 23770 13410
rect 23030 13130 23033 13170
rect 23033 13130 23067 13170
rect 23067 13130 23070 13170
rect 20340 12740 20380 12780
rect 20740 12740 20780 12780
rect 19540 12620 19580 12660
rect 19540 12520 19580 12560
rect 19540 12420 19580 12460
rect 19540 12320 19580 12360
rect 19540 12220 19580 12260
rect 19740 12620 19780 12660
rect 19740 12520 19780 12560
rect 19740 12420 19780 12460
rect 19740 12320 19780 12360
rect 19740 12220 19780 12260
rect 19940 12620 19980 12660
rect 19940 12520 19980 12560
rect 19940 12420 19980 12460
rect 19940 12320 19980 12360
rect 19940 12220 19980 12260
rect 20140 12620 20180 12660
rect 20140 12520 20180 12560
rect 20140 12420 20180 12460
rect 20140 12320 20180 12360
rect 20140 12220 20180 12260
rect 20340 12620 20380 12660
rect 20340 12520 20380 12560
rect 20340 12420 20380 12460
rect 20340 12320 20380 12360
rect 20340 12220 20380 12260
rect 20540 12620 20580 12660
rect 20540 12520 20580 12560
rect 20540 12420 20580 12460
rect 20540 12320 20580 12360
rect 20540 12220 20580 12260
rect 20740 12620 20780 12660
rect 20740 12520 20780 12560
rect 20740 12420 20780 12460
rect 20740 12320 20780 12360
rect 20740 12220 20780 12260
rect 20940 12620 20980 12660
rect 20940 12520 20980 12560
rect 20940 12420 20980 12460
rect 20940 12320 20980 12360
rect 20940 12220 20980 12260
rect 21140 12620 21180 12660
rect 21140 12520 21180 12560
rect 21140 12420 21180 12460
rect 21140 12320 21180 12360
rect 21140 12220 21180 12260
rect 21340 12620 21380 12660
rect 21340 12520 21380 12560
rect 21340 12420 21380 12460
rect 21340 12320 21380 12360
rect 21340 12220 21380 12260
rect 21540 12620 21580 12660
rect 21540 12520 21580 12560
rect 21540 12420 21580 12460
rect 21540 12320 21580 12360
rect 21540 12220 21580 12260
rect 19540 12100 19580 12140
rect 21540 12100 21580 12140
rect 21020 11940 21060 11980
rect 22140 11940 22180 11980
rect 19940 11830 19980 11870
rect 19470 11670 19510 11710
rect 19470 11570 19510 11610
rect 19600 11670 19640 11710
rect 19600 11570 19640 11610
rect 19730 11670 19770 11710
rect 19730 11570 19770 11610
rect 19860 11670 19900 11710
rect 19860 11570 19900 11610
rect 19990 11670 20030 11710
rect 19990 11570 20030 11610
rect 20120 11670 20160 11710
rect 20120 11570 20160 11610
rect 20250 11670 20290 11710
rect 20250 11570 20290 11610
rect 20610 11670 20650 11710
rect 20610 11570 20650 11610
rect 20740 11670 20780 11710
rect 20740 11570 20780 11610
rect 20870 11670 20910 11710
rect 20870 11570 20910 11610
rect 21000 11670 21040 11710
rect 21000 11570 21040 11610
rect 21130 11670 21170 11710
rect 21130 11570 21170 11610
rect 21260 11670 21300 11710
rect 21260 11570 21300 11610
rect 21390 11670 21430 11710
rect 21390 11570 21430 11610
rect 23230 11620 23290 12010
rect 19640 11450 19680 11490
rect 20080 11450 20120 11490
rect 20870 11440 20910 11480
rect 21920 11450 21960 11490
rect 22760 11450 22800 11490
rect 21920 11230 21960 11270
rect 22050 11280 22090 11320
rect 22250 11280 22290 11320
rect 24080 11280 24120 11320
rect 19730 11110 19770 11150
rect 20780 11110 20820 11150
rect 21220 11110 21260 11150
rect 22760 11110 22800 11150
rect 19470 10990 19510 11030
rect 19600 10990 19640 11030
rect 19730 10990 19770 11030
rect 19860 10990 19900 11030
rect 19990 10990 20030 11030
rect 20120 10990 20160 11030
rect 20250 10990 20290 11030
rect 20610 10990 20650 11030
rect 20740 10990 20780 11030
rect 20870 10990 20910 11030
rect 21000 10990 21040 11030
rect 21130 10990 21170 11030
rect 21260 10990 21300 11030
rect 21390 10990 21430 11030
rect 21000 10830 21040 10870
rect 19860 10720 19900 10760
rect 22140 10720 22180 10760
rect 19420 10570 19460 10610
rect 21000 10610 21040 10650
rect 21420 10570 21460 10610
rect 19620 10440 19660 10490
rect 19620 10300 19660 10350
rect 20020 10440 20060 10490
rect 20020 10300 20060 10350
rect 20420 10440 20460 10490
rect 20420 10300 20460 10350
rect 20820 10440 20860 10490
rect 20820 10300 20860 10350
rect 21220 10440 21260 10490
rect 21220 10300 21260 10350
rect 19160 9990 19200 10030
rect 23230 10590 23290 10980
rect 23030 9600 23033 9640
rect 23033 9600 23067 9640
rect 23067 9600 23070 9640
rect 23700 9250 23760 9640
rect 23700 9127 23760 9130
rect 23700 9093 23760 9127
rect 23700 9070 23760 9093
<< metal1 >>
rect 23680 13510 23780 13530
rect 23680 13450 23700 13510
rect 23760 13450 23780 13510
rect 23680 13410 23780 13450
rect 23680 13200 23690 13410
rect 23770 13200 23780 13410
rect 23010 13170 23090 13190
rect 23680 13180 23780 13200
rect 23010 13130 23030 13170
rect 23070 13130 23090 13170
rect 23010 13110 23090 13130
rect 19140 12790 19220 12800
rect 19140 12730 19150 12790
rect 19210 12730 19220 12790
rect 19030 11410 19110 11420
rect 19030 11350 19040 11410
rect 19100 11350 19110 11410
rect 19030 11340 19110 11350
rect 18920 11250 19000 11260
rect 18920 11190 18930 11250
rect 18990 11190 19000 11250
rect 18920 11180 19000 11190
rect 19140 10030 19220 12730
rect 20320 12790 20400 12800
rect 20320 12730 20330 12790
rect 20390 12730 20400 12790
rect 19520 12660 19600 12680
rect 19520 12620 19540 12660
rect 19580 12620 19600 12660
rect 19520 12560 19600 12620
rect 19520 12520 19540 12560
rect 19580 12520 19600 12560
rect 19520 12460 19600 12520
rect 19520 12420 19540 12460
rect 19580 12420 19600 12460
rect 19520 12360 19600 12420
rect 19520 12320 19540 12360
rect 19580 12320 19600 12360
rect 19520 12260 19600 12320
rect 19520 12220 19540 12260
rect 19580 12220 19600 12260
rect 19520 12200 19600 12220
rect 19720 12660 19800 12680
rect 19720 12620 19740 12660
rect 19780 12620 19800 12660
rect 19720 12560 19800 12620
rect 19720 12520 19740 12560
rect 19780 12520 19800 12560
rect 19720 12460 19800 12520
rect 19720 12420 19740 12460
rect 19780 12420 19800 12460
rect 19720 12360 19800 12420
rect 19720 12320 19740 12360
rect 19780 12320 19800 12360
rect 19720 12260 19800 12320
rect 19720 12220 19740 12260
rect 19780 12220 19800 12260
rect 19520 12140 19600 12160
rect 19520 12100 19540 12140
rect 19580 12100 19600 12140
rect 19520 11990 19600 12100
rect 19520 11930 19530 11990
rect 19590 11930 19600 11990
rect 19520 11920 19600 11930
rect 19720 11990 19800 12220
rect 19720 11930 19730 11990
rect 19790 11930 19800 11990
rect 19720 11920 19800 11930
rect 19920 12660 20000 12680
rect 19920 12620 19940 12660
rect 19980 12620 20000 12660
rect 19920 12560 20000 12620
rect 19920 12520 19940 12560
rect 19980 12520 20000 12560
rect 19920 12460 20000 12520
rect 19920 12420 19940 12460
rect 19980 12420 20000 12460
rect 19920 12360 20000 12420
rect 19920 12320 19940 12360
rect 19980 12320 20000 12360
rect 19920 12260 20000 12320
rect 19920 12220 19940 12260
rect 19980 12220 20000 12260
rect 19920 12130 20000 12220
rect 19920 12070 19930 12130
rect 19990 12070 20000 12130
rect 19920 11880 20000 12070
rect 20120 12660 20200 12680
rect 20120 12620 20140 12660
rect 20180 12620 20200 12660
rect 20120 12560 20200 12620
rect 20120 12520 20140 12560
rect 20180 12520 20200 12560
rect 20120 12460 20200 12520
rect 20120 12420 20140 12460
rect 20180 12420 20200 12460
rect 20120 12360 20200 12420
rect 20120 12320 20140 12360
rect 20180 12320 20200 12360
rect 20120 12260 20200 12320
rect 20120 12220 20140 12260
rect 20180 12220 20200 12260
rect 20120 11990 20200 12220
rect 20320 12660 20400 12730
rect 20720 12790 20800 12800
rect 20720 12730 20730 12790
rect 20790 12730 20800 12790
rect 20320 12620 20340 12660
rect 20380 12620 20400 12660
rect 20320 12560 20400 12620
rect 20320 12520 20340 12560
rect 20380 12520 20400 12560
rect 20320 12460 20400 12520
rect 20320 12420 20340 12460
rect 20380 12420 20400 12460
rect 20320 12360 20400 12420
rect 20320 12320 20340 12360
rect 20380 12320 20400 12360
rect 20320 12260 20400 12320
rect 20320 12220 20340 12260
rect 20380 12220 20400 12260
rect 20320 12200 20400 12220
rect 20520 12660 20600 12680
rect 20520 12620 20540 12660
rect 20580 12620 20600 12660
rect 20520 12560 20600 12620
rect 20520 12520 20540 12560
rect 20580 12520 20600 12560
rect 20520 12460 20600 12520
rect 20520 12420 20540 12460
rect 20580 12420 20600 12460
rect 20520 12360 20600 12420
rect 20520 12320 20540 12360
rect 20580 12320 20600 12360
rect 20520 12260 20600 12320
rect 20520 12220 20540 12260
rect 20580 12220 20600 12260
rect 20120 11930 20130 11990
rect 20190 11930 20200 11990
rect 20120 11920 20200 11930
rect 20520 11990 20600 12220
rect 20720 12660 20800 12730
rect 20720 12620 20740 12660
rect 20780 12620 20800 12660
rect 20720 12560 20800 12620
rect 20720 12520 20740 12560
rect 20780 12520 20800 12560
rect 20720 12460 20800 12520
rect 20720 12420 20740 12460
rect 20780 12420 20800 12460
rect 20720 12360 20800 12420
rect 20720 12320 20740 12360
rect 20780 12320 20800 12360
rect 20720 12260 20800 12320
rect 20720 12220 20740 12260
rect 20780 12220 20800 12260
rect 20720 12200 20800 12220
rect 20920 12660 21000 12680
rect 20920 12620 20940 12660
rect 20980 12620 21000 12660
rect 20920 12560 21000 12620
rect 20920 12520 20940 12560
rect 20980 12520 21000 12560
rect 20920 12460 21000 12520
rect 20920 12420 20940 12460
rect 20980 12420 21000 12460
rect 20920 12360 21000 12420
rect 20920 12320 20940 12360
rect 20980 12320 21000 12360
rect 20920 12260 21000 12320
rect 20920 12220 20940 12260
rect 20980 12220 21000 12260
rect 20520 11930 20530 11990
rect 20590 11930 20600 11990
rect 20520 11920 20600 11930
rect 20920 12000 21000 12220
rect 21120 12660 21200 12680
rect 21120 12620 21140 12660
rect 21180 12620 21200 12660
rect 21120 12560 21200 12620
rect 21120 12520 21140 12560
rect 21180 12520 21200 12560
rect 21120 12460 21200 12520
rect 21120 12420 21140 12460
rect 21180 12420 21200 12460
rect 21120 12360 21200 12420
rect 21120 12320 21140 12360
rect 21180 12320 21200 12360
rect 21120 12260 21200 12320
rect 21120 12220 21140 12260
rect 21180 12220 21200 12260
rect 21120 12130 21200 12220
rect 21120 12070 21130 12130
rect 21190 12070 21200 12130
rect 21120 12060 21200 12070
rect 21320 12660 21400 12680
rect 21320 12620 21340 12660
rect 21380 12620 21400 12660
rect 21320 12560 21400 12620
rect 21320 12520 21340 12560
rect 21380 12520 21400 12560
rect 21320 12460 21400 12520
rect 21320 12420 21340 12460
rect 21380 12420 21400 12460
rect 21320 12360 21400 12420
rect 21320 12320 21340 12360
rect 21380 12320 21400 12360
rect 21320 12260 21400 12320
rect 21320 12220 21340 12260
rect 21380 12220 21400 12260
rect 20920 11990 21080 12000
rect 20920 11930 20930 11990
rect 20990 11930 21010 11990
rect 21070 11930 21080 11990
rect 20920 11920 21080 11930
rect 21320 11990 21400 12220
rect 21320 11930 21330 11990
rect 21390 11930 21400 11990
rect 21320 11920 21400 11930
rect 21520 12660 21600 12680
rect 21520 12620 21540 12660
rect 21580 12620 21600 12660
rect 21520 12560 21600 12620
rect 21520 12520 21540 12560
rect 21580 12520 21600 12560
rect 21520 12460 21600 12520
rect 21520 12420 21540 12460
rect 21580 12420 21600 12460
rect 21520 12360 21600 12420
rect 21520 12320 21540 12360
rect 21580 12320 21600 12360
rect 21520 12260 21600 12320
rect 21520 12220 21540 12260
rect 21580 12220 21600 12260
rect 21520 12140 21600 12220
rect 21520 12100 21540 12140
rect 21580 12100 21600 12140
rect 21520 11990 21600 12100
rect 23220 12010 23300 12030
rect 21520 11930 21530 11990
rect 21590 11930 21600 11990
rect 21520 11920 21600 11930
rect 22120 11990 22200 12000
rect 22120 11930 22130 11990
rect 22190 11930 22200 11990
rect 22120 11920 22200 11930
rect 19920 11820 19930 11880
rect 19990 11820 20000 11880
rect 19920 11810 20000 11820
rect 19450 11710 19530 11730
rect 19450 11670 19470 11710
rect 19510 11670 19530 11710
rect 19450 11610 19530 11670
rect 19450 11570 19470 11610
rect 19510 11570 19530 11610
rect 19450 11550 19530 11570
rect 19580 11710 19660 11730
rect 19580 11670 19600 11710
rect 19640 11670 19660 11710
rect 19580 11610 19660 11670
rect 19580 11570 19600 11610
rect 19640 11570 19660 11610
rect 19580 11550 19660 11570
rect 19710 11710 19790 11730
rect 19710 11670 19730 11710
rect 19770 11670 19790 11710
rect 19710 11610 19790 11670
rect 19710 11570 19730 11610
rect 19770 11570 19790 11610
rect 19710 11550 19790 11570
rect 19840 11710 19920 11730
rect 19840 11670 19860 11710
rect 19900 11670 19920 11710
rect 19840 11610 19920 11670
rect 19840 11570 19860 11610
rect 19900 11570 19920 11610
rect 19840 11550 19920 11570
rect 19970 11710 20050 11730
rect 19970 11670 19990 11710
rect 20030 11670 20050 11710
rect 19970 11610 20050 11670
rect 19970 11570 19990 11610
rect 20030 11570 20050 11610
rect 19970 11550 20050 11570
rect 20100 11710 20180 11730
rect 20100 11670 20120 11710
rect 20160 11670 20180 11710
rect 20100 11610 20180 11670
rect 20100 11570 20120 11610
rect 20160 11570 20180 11610
rect 20100 11550 20180 11570
rect 20230 11710 20310 11730
rect 20230 11670 20250 11710
rect 20290 11670 20310 11710
rect 20230 11610 20310 11670
rect 20230 11570 20250 11610
rect 20290 11570 20310 11610
rect 20230 11550 20310 11570
rect 20590 11710 20670 11730
rect 20590 11670 20610 11710
rect 20650 11670 20670 11710
rect 20590 11610 20670 11670
rect 20590 11570 20610 11610
rect 20650 11570 20670 11610
rect 20590 11550 20670 11570
rect 20720 11710 20800 11730
rect 20720 11670 20740 11710
rect 20780 11670 20800 11710
rect 20720 11610 20800 11670
rect 20720 11570 20740 11610
rect 20780 11570 20800 11610
rect 20720 11550 20800 11570
rect 20850 11710 20930 11730
rect 20850 11670 20870 11710
rect 20910 11670 20930 11710
rect 20850 11610 20930 11670
rect 20850 11570 20870 11610
rect 20910 11570 20930 11610
rect 19620 11500 19700 11510
rect 19620 11440 19630 11500
rect 19690 11440 19700 11500
rect 19620 11430 19700 11440
rect 19730 11170 19770 11550
rect 19990 11330 20030 11550
rect 20060 11500 20140 11510
rect 20060 11440 20070 11500
rect 20130 11440 20140 11500
rect 20060 11430 20140 11440
rect 20850 11480 20930 11570
rect 20980 11710 21060 11730
rect 20980 11670 21000 11710
rect 21040 11670 21060 11710
rect 20980 11610 21060 11670
rect 20980 11570 21000 11610
rect 21040 11570 21060 11610
rect 20980 11550 21060 11570
rect 21110 11710 21190 11730
rect 21110 11670 21130 11710
rect 21170 11670 21190 11710
rect 21110 11610 21190 11670
rect 21110 11570 21130 11610
rect 21170 11570 21190 11610
rect 21110 11550 21190 11570
rect 21240 11710 21320 11730
rect 21240 11670 21260 11710
rect 21300 11670 21320 11710
rect 21240 11610 21320 11670
rect 21240 11570 21260 11610
rect 21300 11570 21320 11610
rect 21240 11550 21320 11570
rect 21370 11710 21450 11730
rect 21370 11670 21390 11710
rect 21430 11670 21450 11710
rect 21370 11610 21450 11670
rect 21370 11570 21390 11610
rect 21430 11570 21450 11610
rect 21370 11550 21450 11570
rect 23220 11620 23230 12010
rect 23290 11620 23300 12010
rect 20850 11440 20870 11480
rect 20910 11440 20930 11480
rect 19970 11270 19980 11330
rect 20040 11270 20050 11330
rect 19710 11150 19790 11170
rect 19710 11110 19730 11150
rect 19770 11110 19790 11150
rect 19450 11030 19530 11050
rect 19450 10990 19470 11030
rect 19510 10990 19530 11030
rect 19450 10970 19530 10990
rect 19580 11030 19660 11050
rect 19580 10990 19600 11030
rect 19640 10990 19660 11030
rect 19580 10970 19660 10990
rect 19710 11030 19790 11110
rect 19990 11090 20030 11270
rect 20080 11240 20120 11430
rect 20850 11420 20930 11440
rect 21130 11490 21170 11550
rect 21900 11500 21980 11510
rect 21130 11480 21210 11490
rect 21130 11420 21140 11480
rect 21200 11420 21210 11480
rect 21900 11440 21910 11500
rect 21970 11440 21980 11500
rect 21900 11430 21980 11440
rect 22740 11500 22820 11510
rect 22740 11440 22750 11500
rect 22810 11440 22820 11500
rect 22740 11430 22820 11440
rect 23220 11500 23300 11620
rect 23220 11440 23230 11500
rect 23290 11440 23300 11500
rect 23220 11430 23300 11440
rect 24040 11580 24150 11600
rect 24040 11510 24060 11580
rect 24130 11510 24150 11580
rect 20720 11350 20730 11410
rect 20790 11350 20800 11410
rect 20060 11230 20140 11240
rect 20060 11170 20070 11230
rect 20130 11170 20140 11230
rect 20060 11160 20140 11170
rect 20760 11170 20800 11350
rect 20760 11160 20840 11170
rect 20760 11100 20770 11160
rect 20830 11100 20840 11160
rect 20760 11090 20840 11100
rect 19710 10990 19730 11030
rect 19770 10990 19790 11030
rect 19710 10970 19790 10990
rect 19840 11030 19920 11050
rect 19840 10990 19860 11030
rect 19900 10990 19920 11030
rect 19840 10970 19920 10990
rect 19970 11030 20050 11090
rect 20870 11050 20910 11420
rect 21130 11410 21210 11420
rect 21130 11050 21170 11410
rect 22030 11330 22110 11340
rect 21900 11280 21980 11290
rect 21900 11220 21910 11280
rect 21970 11220 21980 11280
rect 22030 11270 22040 11330
rect 22100 11270 22110 11330
rect 22030 11260 22110 11270
rect 22230 11330 22310 11340
rect 22230 11270 22240 11330
rect 22300 11270 22310 11330
rect 22230 11260 22310 11270
rect 24040 11330 24150 11510
rect 24040 11270 24070 11330
rect 24130 11270 24150 11330
rect 21900 11210 21980 11220
rect 21200 11160 21280 11170
rect 21200 11100 21210 11160
rect 21270 11100 21280 11160
rect 21200 11090 21280 11100
rect 22740 11160 22820 11170
rect 22740 11100 22750 11160
rect 22810 11100 22820 11160
rect 22740 11090 22820 11100
rect 23220 11160 23300 11170
rect 23220 11100 23230 11160
rect 23290 11100 23300 11160
rect 19970 10990 19990 11030
rect 20030 10990 20050 11030
rect 19970 10970 20050 10990
rect 20100 11030 20180 11050
rect 20100 10990 20120 11030
rect 20160 10990 20180 11030
rect 20100 10970 20180 10990
rect 20230 11030 20310 11050
rect 20230 10990 20250 11030
rect 20290 10990 20310 11030
rect 20230 10970 20310 10990
rect 20590 11030 20670 11050
rect 20590 10990 20610 11030
rect 20650 10990 20670 11030
rect 20590 10970 20670 10990
rect 20720 11030 20800 11050
rect 20720 10990 20740 11030
rect 20780 10990 20800 11030
rect 20720 10970 20800 10990
rect 20850 11030 20930 11050
rect 20850 10990 20870 11030
rect 20910 10990 20930 11030
rect 20850 10970 20930 10990
rect 20980 11030 21060 11050
rect 20980 10990 21000 11030
rect 21040 10990 21060 11030
rect 20980 10970 21060 10990
rect 21110 11030 21190 11050
rect 21110 10990 21130 11030
rect 21170 10990 21190 11030
rect 21110 10970 21190 10990
rect 21240 11030 21320 11050
rect 21240 10990 21260 11030
rect 21300 10990 21320 11030
rect 21240 10970 21320 10990
rect 21370 11030 21450 11050
rect 21370 10990 21390 11030
rect 21430 10990 21450 11030
rect 21370 10970 21450 10990
rect 23220 10980 23300 11100
rect 24040 11070 24150 11270
rect 24040 11000 24060 11070
rect 24130 11000 24150 11070
rect 24040 10980 24150 11000
rect 20980 10880 21060 10890
rect 20980 10820 20990 10880
rect 21050 10820 21060 10880
rect 19400 10770 19480 10780
rect 19400 10710 19410 10770
rect 19470 10710 19480 10770
rect 19400 10610 19480 10710
rect 19400 10570 19420 10610
rect 19460 10570 19480 10610
rect 19400 10550 19480 10570
rect 19600 10770 19680 10780
rect 19600 10710 19610 10770
rect 19670 10710 19680 10770
rect 19600 10490 19680 10710
rect 19840 10770 19920 10780
rect 19840 10710 19850 10770
rect 19910 10710 19920 10770
rect 19840 10700 19920 10710
rect 20000 10770 20080 10780
rect 20000 10710 20010 10770
rect 20070 10710 20080 10770
rect 19600 10440 19620 10490
rect 19660 10440 19680 10490
rect 19600 10350 19680 10440
rect 19600 10300 19620 10350
rect 19660 10300 19680 10350
rect 19600 10280 19680 10300
rect 20000 10490 20080 10710
rect 20000 10440 20020 10490
rect 20060 10440 20080 10490
rect 20000 10350 20080 10440
rect 20000 10300 20020 10350
rect 20060 10300 20080 10350
rect 20000 10280 20080 10300
rect 20400 10770 20480 10780
rect 20400 10710 20410 10770
rect 20470 10710 20480 10770
rect 20400 10490 20480 10710
rect 20400 10440 20420 10490
rect 20460 10440 20480 10490
rect 20400 10350 20480 10440
rect 20400 10300 20420 10350
rect 20460 10300 20480 10350
rect 20400 10280 20480 10300
rect 20800 10770 20880 10780
rect 20800 10710 20810 10770
rect 20870 10710 20880 10770
rect 20800 10490 20880 10710
rect 20980 10660 21060 10820
rect 20980 10600 20990 10660
rect 21050 10600 21060 10660
rect 20980 10590 21060 10600
rect 21200 10770 21280 10780
rect 21200 10710 21210 10770
rect 21270 10710 21280 10770
rect 20800 10440 20820 10490
rect 20860 10440 20880 10490
rect 20800 10350 20880 10440
rect 20800 10300 20820 10350
rect 20860 10300 20880 10350
rect 20800 10280 20880 10300
rect 21200 10490 21280 10710
rect 21400 10770 21480 10780
rect 21400 10710 21410 10770
rect 21470 10710 21480 10770
rect 21400 10610 21480 10710
rect 22120 10770 22200 10780
rect 22120 10710 22130 10770
rect 22190 10710 22200 10770
rect 22120 10700 22200 10710
rect 21400 10570 21420 10610
rect 21460 10570 21480 10610
rect 23220 10590 23230 10980
rect 23290 10590 23300 10980
rect 23220 10570 23300 10590
rect 21400 10550 21480 10570
rect 21200 10440 21220 10490
rect 21260 10440 21280 10490
rect 21200 10350 21280 10440
rect 21200 10300 21220 10350
rect 21260 10300 21280 10350
rect 21200 10280 21280 10300
rect 19140 9990 19160 10030
rect 19200 9990 19220 10030
rect 19140 9970 19220 9990
rect 23010 9650 23090 9660
rect 23010 9590 23020 9650
rect 23080 9590 23090 9650
rect 23010 9580 23090 9590
rect 23680 9640 23780 9660
rect 23680 9250 23700 9640
rect 23760 9250 23780 9640
rect 23680 9130 23780 9250
rect 23680 9070 23700 9130
rect 23760 9070 23780 9130
rect 23680 9050 23780 9070
<< via1 >>
rect 23700 13450 23760 13510
rect 19150 12730 19210 12790
rect 19040 11350 19100 11410
rect 18930 11190 18990 11250
rect 20330 12780 20390 12790
rect 20330 12740 20340 12780
rect 20340 12740 20380 12780
rect 20380 12740 20390 12780
rect 20330 12730 20390 12740
rect 19530 11930 19590 11990
rect 19730 11930 19790 11990
rect 19930 12070 19990 12130
rect 20730 12780 20790 12790
rect 20730 12740 20740 12780
rect 20740 12740 20780 12780
rect 20780 12740 20790 12780
rect 20730 12730 20790 12740
rect 20130 11930 20190 11990
rect 20530 11930 20590 11990
rect 21130 12070 21190 12130
rect 20930 11930 20990 11990
rect 21010 11980 21070 11990
rect 21010 11940 21020 11980
rect 21020 11940 21060 11980
rect 21060 11940 21070 11980
rect 21010 11930 21070 11940
rect 21330 11930 21390 11990
rect 21530 11930 21590 11990
rect 22130 11980 22190 11990
rect 22130 11940 22140 11980
rect 22140 11940 22180 11980
rect 22180 11940 22190 11980
rect 22130 11930 22190 11940
rect 19930 11870 19990 11880
rect 19930 11830 19940 11870
rect 19940 11830 19980 11870
rect 19980 11830 19990 11870
rect 19930 11820 19990 11830
rect 19630 11490 19690 11500
rect 19630 11450 19640 11490
rect 19640 11450 19680 11490
rect 19680 11450 19690 11490
rect 19630 11440 19690 11450
rect 20070 11490 20130 11500
rect 20070 11450 20080 11490
rect 20080 11450 20120 11490
rect 20120 11450 20130 11490
rect 20070 11440 20130 11450
rect 19980 11270 20040 11330
rect 21140 11420 21200 11480
rect 21910 11490 21970 11500
rect 21910 11450 21920 11490
rect 21920 11450 21960 11490
rect 21960 11450 21970 11490
rect 21910 11440 21970 11450
rect 22750 11490 22810 11500
rect 22750 11450 22760 11490
rect 22760 11450 22800 11490
rect 22800 11450 22810 11490
rect 22750 11440 22810 11450
rect 23230 11440 23290 11500
rect 24060 11510 24130 11580
rect 20730 11350 20790 11410
rect 20070 11170 20130 11230
rect 20770 11150 20830 11160
rect 20770 11110 20780 11150
rect 20780 11110 20820 11150
rect 20820 11110 20830 11150
rect 20770 11100 20830 11110
rect 21910 11270 21970 11280
rect 21910 11230 21920 11270
rect 21920 11230 21960 11270
rect 21960 11230 21970 11270
rect 21910 11220 21970 11230
rect 22040 11320 22100 11330
rect 22040 11280 22050 11320
rect 22050 11280 22090 11320
rect 22090 11280 22100 11320
rect 22040 11270 22100 11280
rect 22240 11320 22300 11330
rect 22240 11280 22250 11320
rect 22250 11280 22290 11320
rect 22290 11280 22300 11320
rect 22240 11270 22300 11280
rect 24070 11320 24130 11330
rect 24070 11280 24080 11320
rect 24080 11280 24120 11320
rect 24120 11280 24130 11320
rect 24070 11270 24130 11280
rect 21210 11150 21270 11160
rect 21210 11110 21220 11150
rect 21220 11110 21260 11150
rect 21260 11110 21270 11150
rect 21210 11100 21270 11110
rect 22750 11150 22810 11160
rect 22750 11110 22760 11150
rect 22760 11110 22800 11150
rect 22800 11110 22810 11150
rect 22750 11100 22810 11110
rect 23230 11100 23290 11160
rect 24060 11000 24130 11070
rect 20990 10870 21050 10880
rect 20990 10830 21000 10870
rect 21000 10830 21040 10870
rect 21040 10830 21050 10870
rect 20990 10820 21050 10830
rect 19410 10710 19470 10770
rect 19610 10710 19670 10770
rect 19850 10760 19910 10770
rect 19850 10720 19860 10760
rect 19860 10720 19900 10760
rect 19900 10720 19910 10760
rect 19850 10710 19910 10720
rect 20010 10710 20070 10770
rect 20410 10710 20470 10770
rect 20810 10710 20870 10770
rect 20990 10650 21050 10660
rect 20990 10610 21000 10650
rect 21000 10610 21040 10650
rect 21040 10610 21050 10650
rect 20990 10600 21050 10610
rect 21210 10710 21270 10770
rect 21410 10710 21470 10770
rect 22130 10760 22190 10770
rect 22130 10720 22140 10760
rect 22140 10720 22180 10760
rect 22180 10720 22190 10760
rect 22130 10710 22190 10720
rect 23020 9640 23080 9650
rect 23020 9600 23030 9640
rect 23030 9600 23070 9640
rect 23070 9600 23080 9640
rect 23020 9590 23080 9600
rect 23700 9070 23760 9130
<< metal2 >>
rect 23680 13510 23780 13530
rect 23680 13450 23700 13510
rect 23760 13450 23780 13510
rect 23680 13430 23780 13450
rect 18790 13110 23010 13190
rect 19140 12790 20800 12800
rect 19140 12730 19150 12790
rect 19210 12730 20330 12790
rect 20390 12730 20730 12790
rect 20790 12730 20800 12790
rect 19140 12720 20800 12730
rect 19920 12130 21200 12140
rect 19920 12070 19930 12130
rect 19990 12070 21130 12130
rect 21190 12070 21200 12130
rect 19920 12060 21200 12070
rect 18790 11990 22200 12000
rect 18790 11930 19530 11990
rect 19590 11930 19730 11990
rect 19790 11930 20130 11990
rect 20190 11930 20530 11990
rect 20590 11930 20930 11990
rect 20990 11930 21010 11990
rect 21070 11930 21330 11990
rect 21390 11930 21530 11990
rect 21590 11930 22130 11990
rect 22190 11930 22200 11990
rect 18790 11920 22200 11930
rect 19920 11880 20000 11890
rect 19920 11820 19930 11880
rect 19990 11820 20000 11880
rect 19920 11810 20000 11820
rect 24040 11580 24150 11600
rect 24040 11510 24060 11580
rect 24130 11510 24150 11580
rect 19620 11500 19700 11510
rect 19620 11440 19630 11500
rect 19690 11440 19700 11500
rect 19030 11410 19110 11420
rect 19030 11350 19040 11410
rect 19100 11400 19110 11410
rect 19620 11400 19700 11440
rect 20060 11500 20140 11510
rect 20060 11440 20070 11500
rect 20130 11440 20140 11500
rect 21900 11500 21980 11510
rect 20060 11430 20140 11440
rect 21130 11480 21210 11490
rect 21130 11420 21140 11480
rect 21200 11470 21210 11480
rect 21900 11470 21910 11500
rect 21200 11440 21910 11470
rect 21970 11440 21980 11500
rect 21200 11430 21980 11440
rect 22740 11500 23300 11510
rect 22740 11440 22750 11500
rect 22810 11440 23230 11500
rect 23290 11440 23300 11500
rect 24040 11490 24150 11510
rect 22740 11430 23300 11440
rect 21200 11420 21210 11430
rect 21130 11410 21210 11420
rect 20720 11400 20730 11410
rect 19100 11360 20730 11400
rect 19100 11350 19110 11360
rect 20720 11350 20730 11360
rect 20790 11350 20800 11410
rect 19030 11340 19110 11350
rect 22030 11330 26450 11340
rect 19970 11270 19980 11330
rect 20040 11320 20050 11330
rect 20040 11280 21980 11320
rect 20040 11270 20050 11280
rect 18920 11250 19000 11260
rect 18920 11190 18930 11250
rect 18990 11240 19000 11250
rect 18990 11230 21280 11240
rect 18990 11200 20070 11230
rect 18990 11190 19000 11200
rect 18920 11180 19000 11190
rect 20060 11170 20070 11200
rect 20130 11200 21280 11230
rect 21900 11220 21910 11280
rect 21970 11220 21980 11280
rect 22030 11270 22040 11330
rect 22100 11270 22240 11330
rect 22300 11270 24070 11330
rect 24130 11270 26450 11330
rect 22030 11260 26450 11270
rect 21900 11210 21980 11220
rect 20130 11170 20140 11200
rect 20060 11160 20140 11170
rect 20760 11160 20840 11170
rect 20760 11100 20770 11160
rect 20830 11100 20840 11160
rect 20760 11090 20840 11100
rect 21200 11160 21280 11200
rect 21200 11100 21210 11160
rect 21270 11100 21280 11160
rect 21200 11090 21280 11100
rect 22740 11160 23300 11170
rect 22740 11100 22750 11160
rect 22810 11100 23230 11160
rect 23290 11100 23300 11160
rect 22740 11090 23300 11100
rect 24040 11070 24150 11090
rect 24040 11000 24060 11070
rect 24130 11000 24150 11070
rect 24040 10980 24150 11000
rect 20980 10880 21060 10890
rect 20980 10820 20990 10880
rect 21050 10820 21060 10880
rect 20980 10810 21060 10820
rect 18790 10770 22200 10780
rect 18790 10710 19410 10770
rect 19470 10710 19610 10770
rect 19670 10710 19850 10770
rect 19910 10710 20010 10770
rect 20070 10710 20410 10770
rect 20470 10710 20810 10770
rect 20870 10710 21210 10770
rect 21270 10710 21410 10770
rect 21470 10710 22130 10770
rect 22190 10710 22200 10770
rect 18790 10700 22200 10710
rect 20980 10660 21060 10670
rect 20980 10600 20990 10660
rect 21050 10600 21060 10660
rect 20980 10590 21060 10600
rect 18790 9650 23090 9660
rect 18790 9590 23020 9650
rect 23080 9590 23090 9650
rect 18790 9580 23090 9590
rect 23680 9130 23780 9150
rect 23680 9070 23700 9130
rect 23760 9070 23780 9130
rect 23680 9050 23780 9070
<< via2 >>
rect 23700 13450 23760 13510
rect 24060 11510 24130 11580
rect 24060 11000 24130 11070
rect 23700 9070 23760 9130
<< metal3 >>
rect 23680 13520 23780 13530
rect 23680 13510 26450 13520
rect 23680 13450 23700 13510
rect 23760 13450 26450 13510
rect 23680 13430 26450 13450
rect 24040 11580 24150 11600
rect 24040 11510 24060 11580
rect 24130 11510 24150 11580
rect 24040 11490 24150 11510
rect 24390 11460 26450 13430
rect 24040 11070 24150 11090
rect 24040 11000 24060 11070
rect 24130 11000 24150 11070
rect 24040 10980 24150 11000
rect 24390 9150 26450 11120
rect 23680 9130 26450 9150
rect 23680 9070 23700 9130
rect 23760 9070 26450 9130
rect 23680 9060 26450 9070
rect 23680 9050 23780 9060
<< via3 >>
rect 24060 11510 24130 11580
rect 24060 11000 24130 11070
<< mimcap >>
rect 24420 11580 26420 13490
rect 24420 11510 24440 11580
rect 24510 11510 26420 11580
rect 24420 11490 26420 11510
rect 24420 11070 26420 11090
rect 24420 11000 24440 11070
rect 24510 11000 26420 11070
rect 24420 9090 26420 11000
<< mimcapcontact >>
rect 24440 11510 24510 11580
rect 24440 11000 24510 11070
<< metal4 >>
rect 24040 11580 24520 11600
rect 24040 11510 24060 11580
rect 24130 11510 24440 11580
rect 24510 11510 24520 11580
rect 24040 11490 24520 11510
rect 24040 11070 24520 11090
rect 24040 11000 24060 11070
rect 24130 11000 24440 11070
rect 24510 11000 24520 11070
rect 24040 10980 24520 11000
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
