magic
tech sky130A
magscale 1 2
timestamp 1757089566
<< nwell >>
rect 14817 19209 17503 19733
<< nsubdiff >>
rect 14853 19663 14949 19697
rect 17371 19663 17467 19697
rect 14853 19601 14887 19663
rect 17433 19601 17467 19663
rect 14853 19279 14887 19341
rect 17433 19279 17467 19341
rect 14853 19245 14949 19279
rect 17371 19245 17467 19279
<< nsubdiffcont >>
rect 14949 19663 17371 19697
rect 14853 19341 14887 19601
rect 17433 19341 17467 19601
rect 14949 19245 17371 19279
<< xpolycontact >>
rect 14992 19436 15424 19506
rect 16896 19436 17328 19506
<< xpolyres >>
rect 15424 19436 16896 19506
<< locali >>
rect 16120 19697 16200 19700
rect 14853 19663 14949 19697
rect 17371 19663 17467 19697
rect 14853 19601 14887 19663
rect 16120 19640 16140 19663
rect 16180 19640 16200 19663
rect 16120 19620 16200 19640
rect 17433 19601 17467 19663
rect 14853 19279 14887 19341
rect 17433 19279 17467 19341
rect 14853 19245 14949 19279
rect 17371 19245 17467 19279
<< viali >>
rect 16140 19663 16180 19680
rect 16140 19640 16180 19663
rect 15010 19452 15407 19490
rect 16913 19452 17310 19490
<< metal1 >>
rect 16120 19690 16200 19700
rect 16120 19630 16130 19690
rect 16190 19630 16200 19690
rect 16120 19620 16200 19630
rect 14990 19500 15420 19510
rect 14990 19440 15000 19500
rect 15410 19440 15420 19500
rect 14990 19430 15420 19440
rect 16900 19500 17330 19510
rect 16900 19440 16910 19500
rect 17320 19440 17330 19500
rect 16900 19430 17330 19440
rect 25990 19500 26090 19520
rect 25990 19440 26010 19500
rect 26070 19440 26090 19500
rect 25990 19420 26090 19440
<< via1 >>
rect 16130 19680 16190 19690
rect 16130 19640 16140 19680
rect 16140 19640 16180 19680
rect 16180 19640 16190 19680
rect 16130 19630 16190 19640
rect 15000 19490 15410 19500
rect 15000 19452 15010 19490
rect 15010 19452 15407 19490
rect 15407 19452 15410 19490
rect 15000 19440 15410 19452
rect 16910 19490 17320 19500
rect 16910 19452 16913 19490
rect 16913 19452 17310 19490
rect 17310 19452 17320 19490
rect 16910 19440 17320 19452
rect 26010 19440 26070 19500
<< metal2 >>
rect 7720 19790 23410 19810
rect 7720 19720 22820 19790
rect 22890 19720 23320 19790
rect 23390 19720 23410 19790
rect 7720 19700 23410 19720
rect 16120 19690 16200 19700
rect 16120 19630 16130 19690
rect 16190 19630 16200 19690
rect 16120 19620 16200 19630
rect 8920 19510 9020 19520
rect 25990 19510 26090 19520
rect 8920 19500 15420 19510
rect 8920 19440 8940 19500
rect 9000 19440 15000 19500
rect 15410 19440 15420 19500
rect 8920 19430 15420 19440
rect 16900 19500 26090 19510
rect 16900 19440 16910 19500
rect 17320 19440 26010 19500
rect 26070 19440 26090 19500
rect 16900 19430 26090 19440
rect 8920 19420 9020 19430
rect 25990 19420 26090 19430
<< via2 >>
rect 22820 19720 22890 19790
rect 23320 19720 23390 19790
rect 8940 19440 9000 19500
rect 26010 19440 26070 19500
<< metal3 >>
rect 8920 20050 22940 32110
rect 23270 20050 26090 32110
rect 8920 19500 9020 20050
rect 22800 19790 22910 19810
rect 22800 19720 22820 19790
rect 22890 19720 22910 19790
rect 22800 19700 22910 19720
rect 23300 19790 23410 19810
rect 23300 19720 23320 19790
rect 23390 19720 23410 19790
rect 23300 19700 23410 19720
rect 8920 19440 8940 19500
rect 9000 19440 9020 19500
rect 8920 19420 9020 19440
rect 25990 19500 26090 20050
rect 25990 19440 26010 19500
rect 26070 19440 26090 19500
rect 25990 19420 26090 19440
<< via3 >>
rect 22820 19720 22890 19790
rect 23320 19720 23390 19790
<< mimcap >>
rect 8950 20170 22910 32080
rect 8950 20100 22820 20170
rect 22890 20100 22910 20170
rect 8950 20080 22910 20100
rect 23300 20170 26060 32080
rect 23300 20100 23320 20170
rect 23390 20100 26060 20170
rect 23300 20080 26060 20100
<< mimcapcontact >>
rect 22820 20100 22890 20170
rect 23320 20100 23390 20170
<< metal4 >>
rect 22800 20170 22910 20180
rect 22800 20100 22820 20170
rect 22890 20100 22910 20170
rect 22800 19790 22910 20100
rect 22800 19720 22820 19790
rect 22890 19720 22910 19790
rect 22800 19700 22910 19720
rect 23300 20170 23410 20180
rect 23300 20100 23320 20170
rect 23390 20100 23410 20170
rect 23300 19790 23410 20100
rect 23300 19720 23320 19790
rect 23390 19720 23410 19790
rect 23300 19700 23410 19720
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
