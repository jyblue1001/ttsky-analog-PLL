magic
tech sky130A
magscale 1 2
timestamp 1757102137
<< error_p >>
rect 8564 17176 8668 17420
rect 9683 16777 9787 17567
rect 16897 17383 17001 17940
rect 17684 17176 17788 17940
rect 10210 16782 10314 17036
rect 10464 16246 10568 16782
rect 16116 16246 16220 17036
rect 13240 14650 13320 14754
<< nwell >>
rect 8227 17041 8751 18633
rect 9014 16642 9870 18636
rect 10127 16111 10983 18633
rect 15447 16111 16303 18633
rect 16560 17248 17084 18630
rect 17347 17041 17871 18633
rect 10400 11580 13130 11860
rect 13430 11580 16160 11860
rect 11500 10020 15060 10700
rect 15360 10220 16130 10500
rect 11510 9420 13150 9700
rect 13410 9420 15050 9700
<< pwell >>
rect 13240 18810 13320 19090
rect 11250 18657 12590 18810
rect 11250 17623 11403 18657
rect 12437 17623 12590 18657
rect 11250 17470 12590 17623
rect 12610 18657 13950 18810
rect 12610 17623 12763 18657
rect 13797 17623 13950 18657
rect 12610 17470 13950 17623
rect 13970 18657 15310 18810
rect 13970 17623 14123 18657
rect 15157 17623 15310 18657
rect 13970 17470 15310 17623
rect 11250 17297 12590 17450
rect 11250 16263 11403 17297
rect 12437 16263 12590 17297
rect 11250 16110 12590 16263
rect 12610 17297 13950 17450
rect 12610 16263 12763 17297
rect 13797 16263 13950 17297
rect 12610 16110 13950 16263
rect 13970 17297 15310 17450
rect 13970 16263 14123 17297
rect 15157 16263 15310 17297
rect 13970 16110 15310 16263
rect 11250 15937 12590 16090
rect 11250 14903 11403 15937
rect 12437 14903 12590 15937
rect 11250 14750 12590 14903
rect 12610 15937 13950 16090
rect 12610 14903 12763 15937
rect 13797 14903 13950 15937
rect 12610 14750 13950 14903
rect 13970 15937 15310 16090
rect 13970 14903 14123 15937
rect 15157 14903 15310 15937
rect 13970 14750 15310 14903
<< nbase >>
rect 11403 17623 12437 18657
rect 12763 17623 13797 18657
rect 14123 17623 15157 18657
rect 11403 16263 12437 17297
rect 12763 16263 13797 17297
rect 14123 16263 15157 17297
rect 11403 14903 12437 15937
rect 12763 14903 13797 15937
rect 14123 14903 15157 15937
<< nmos >>
rect 11240 14080 13240 14280
rect 13320 14080 15320 14280
rect 10820 13170 11820 13670
rect 12060 13170 13060 13670
rect 13500 13170 14500 13670
rect 14740 13170 15740 13670
rect 11440 12560 11480 12660
rect 11560 12560 11600 12660
rect 11680 12560 11720 12660
rect 11800 12560 11840 12660
rect 11920 12560 11960 12660
rect 12040 12560 12080 12660
rect 12160 12560 12200 12660
rect 12280 12560 12320 12660
rect 12400 12560 12440 12660
rect 12520 12560 12560 12660
rect 14000 12560 14040 12660
rect 14120 12560 14160 12660
rect 14240 12560 14280 12660
rect 14360 12560 14400 12660
rect 14480 12560 14520 12660
rect 14600 12560 14640 12660
rect 14720 12560 14760 12660
rect 14840 12560 14880 12660
rect 14960 12560 15000 12660
rect 15080 12560 15120 12660
<< pmos >>
rect 10600 11620 10640 11820
rect 10720 11620 10760 11820
rect 10840 11620 10880 11820
rect 10960 11620 11000 11820
rect 11080 11620 11120 11820
rect 11200 11620 11240 11820
rect 11320 11620 11360 11820
rect 11440 11620 11480 11820
rect 11560 11620 11600 11820
rect 11680 11620 11720 11820
rect 11800 11620 11840 11820
rect 11920 11620 11960 11820
rect 12040 11620 12080 11820
rect 12160 11620 12200 11820
rect 12280 11620 12320 11820
rect 12400 11620 12440 11820
rect 12520 11620 12560 11820
rect 12640 11620 12680 11820
rect 12760 11620 12800 11820
rect 12880 11620 12920 11820
rect 13640 11620 13680 11820
rect 13760 11620 13800 11820
rect 13880 11620 13920 11820
rect 14000 11620 14040 11820
rect 14120 11620 14160 11820
rect 14240 11620 14280 11820
rect 14360 11620 14400 11820
rect 14480 11620 14520 11820
rect 14600 11620 14640 11820
rect 14720 11620 14760 11820
rect 14840 11620 14880 11820
rect 14960 11620 15000 11820
rect 15080 11620 15120 11820
rect 15200 11620 15240 11820
rect 15320 11620 15360 11820
rect 15440 11620 15480 11820
rect 15560 11620 15600 11820
rect 15680 11620 15720 11820
rect 15800 11620 15840 11820
rect 15920 11620 15960 11820
rect 11700 10060 11800 10660
rect 11880 10060 11980 10660
rect 12060 10060 12160 10660
rect 12240 10060 12340 10660
rect 12420 10060 12520 10660
rect 12600 10060 12700 10660
rect 12780 10060 12880 10660
rect 12960 10060 13060 10660
rect 13140 10060 13240 10660
rect 13320 10060 13420 10660
rect 13500 10060 13600 10660
rect 13680 10060 13780 10660
rect 13860 10060 13960 10660
rect 14040 10060 14140 10660
rect 14220 10060 14320 10660
rect 14400 10060 14500 10660
rect 14580 10060 14680 10660
rect 14760 10060 14860 10660
rect 15570 10260 15600 10460
rect 15680 10260 15710 10460
rect 15790 10260 15820 10460
rect 15900 10260 15930 10460
rect 11710 9460 11740 9660
rect 11820 9460 11850 9660
rect 11930 9460 11960 9660
rect 12040 9460 12070 9660
rect 12150 9460 12180 9660
rect 12260 9460 12290 9660
rect 12370 9460 12400 9660
rect 12480 9460 12510 9660
rect 12590 9460 12620 9660
rect 12700 9460 12730 9660
rect 12810 9460 12840 9660
rect 12920 9460 12950 9660
rect 13610 9460 13640 9660
rect 13720 9460 13750 9660
rect 13830 9460 13860 9660
rect 13940 9460 13970 9660
rect 14050 9460 14080 9660
rect 14160 9460 14190 9660
rect 14270 9460 14300 9660
rect 14380 9460 14410 9660
rect 14490 9460 14520 9660
rect 14600 9460 14630 9660
rect 14710 9460 14740 9660
rect 14820 9460 14850 9660
<< ndiff >>
rect 11160 14250 11240 14280
rect 11160 14210 11180 14250
rect 11220 14210 11240 14250
rect 11160 14150 11240 14210
rect 11160 14110 11180 14150
rect 11220 14110 11240 14150
rect 11160 14080 11240 14110
rect 13240 14250 13320 14280
rect 13240 14210 13260 14250
rect 13300 14210 13320 14250
rect 13240 14150 13320 14210
rect 13240 14110 13260 14150
rect 13300 14110 13320 14150
rect 13240 14080 13320 14110
rect 15320 14250 15400 14280
rect 15320 14210 15340 14250
rect 15380 14210 15400 14250
rect 15320 14150 15400 14210
rect 15320 14110 15340 14150
rect 15380 14110 15400 14150
rect 15320 14080 15400 14110
rect 10740 13640 10820 13670
rect 10740 13600 10760 13640
rect 10800 13600 10820 13640
rect 10740 13540 10820 13600
rect 10740 13500 10760 13540
rect 10800 13500 10820 13540
rect 10740 13440 10820 13500
rect 10740 13400 10760 13440
rect 10800 13400 10820 13440
rect 10740 13340 10820 13400
rect 10740 13300 10760 13340
rect 10800 13300 10820 13340
rect 10740 13240 10820 13300
rect 10740 13200 10760 13240
rect 10800 13200 10820 13240
rect 10740 13170 10820 13200
rect 11820 13640 11900 13670
rect 11980 13640 12060 13670
rect 11820 13600 11840 13640
rect 11880 13600 11900 13640
rect 11980 13600 12000 13640
rect 12040 13600 12060 13640
rect 11820 13540 11900 13600
rect 11980 13540 12060 13600
rect 11820 13500 11840 13540
rect 11880 13500 11900 13540
rect 11980 13500 12000 13540
rect 12040 13500 12060 13540
rect 11820 13440 11900 13500
rect 11980 13440 12060 13500
rect 11820 13400 11840 13440
rect 11880 13400 11900 13440
rect 11980 13400 12000 13440
rect 12040 13400 12060 13440
rect 11820 13340 11900 13400
rect 11980 13340 12060 13400
rect 11820 13300 11840 13340
rect 11880 13300 11900 13340
rect 11980 13300 12000 13340
rect 12040 13300 12060 13340
rect 11820 13240 11900 13300
rect 11980 13240 12060 13300
rect 11820 13200 11840 13240
rect 11880 13200 11900 13240
rect 11980 13200 12000 13240
rect 12040 13200 12060 13240
rect 11820 13170 11900 13200
rect 11980 13170 12060 13200
rect 13060 13640 13140 13670
rect 13060 13600 13080 13640
rect 13120 13600 13140 13640
rect 13060 13540 13140 13600
rect 13060 13500 13080 13540
rect 13120 13500 13140 13540
rect 13060 13440 13140 13500
rect 13060 13400 13080 13440
rect 13120 13400 13140 13440
rect 13060 13340 13140 13400
rect 13060 13300 13080 13340
rect 13120 13300 13140 13340
rect 13060 13240 13140 13300
rect 13060 13200 13080 13240
rect 13120 13200 13140 13240
rect 13060 13170 13140 13200
rect 13420 13640 13500 13670
rect 13420 13600 13440 13640
rect 13480 13600 13500 13640
rect 13420 13540 13500 13600
rect 13420 13500 13440 13540
rect 13480 13500 13500 13540
rect 13420 13440 13500 13500
rect 13420 13400 13440 13440
rect 13480 13400 13500 13440
rect 13420 13340 13500 13400
rect 13420 13300 13440 13340
rect 13480 13300 13500 13340
rect 13420 13240 13500 13300
rect 13420 13200 13440 13240
rect 13480 13200 13500 13240
rect 13420 13170 13500 13200
rect 14500 13640 14580 13670
rect 14660 13640 14740 13670
rect 14500 13600 14520 13640
rect 14560 13600 14580 13640
rect 14660 13600 14680 13640
rect 14720 13600 14740 13640
rect 14500 13540 14580 13600
rect 14660 13540 14740 13600
rect 14500 13500 14520 13540
rect 14560 13500 14580 13540
rect 14660 13500 14680 13540
rect 14720 13500 14740 13540
rect 14500 13440 14580 13500
rect 14660 13440 14740 13500
rect 14500 13400 14520 13440
rect 14560 13400 14580 13440
rect 14660 13400 14680 13440
rect 14720 13400 14740 13440
rect 14500 13340 14580 13400
rect 14660 13340 14740 13400
rect 14500 13300 14520 13340
rect 14560 13300 14580 13340
rect 14660 13300 14680 13340
rect 14720 13300 14740 13340
rect 14500 13240 14580 13300
rect 14660 13240 14740 13300
rect 14500 13200 14520 13240
rect 14560 13200 14580 13240
rect 14660 13200 14680 13240
rect 14720 13200 14740 13240
rect 14500 13170 14580 13200
rect 14660 13170 14740 13200
rect 15740 13640 15820 13670
rect 15740 13600 15760 13640
rect 15800 13600 15820 13640
rect 15740 13540 15820 13600
rect 15740 13500 15760 13540
rect 15800 13500 15820 13540
rect 15740 13440 15820 13500
rect 15740 13400 15760 13440
rect 15800 13400 15820 13440
rect 15740 13340 15820 13400
rect 15740 13300 15760 13340
rect 15800 13300 15820 13340
rect 15740 13240 15820 13300
rect 15740 13200 15760 13240
rect 15800 13200 15820 13240
rect 15740 13170 15820 13200
rect 11360 12630 11440 12660
rect 11360 12590 11380 12630
rect 11420 12590 11440 12630
rect 11360 12560 11440 12590
rect 11480 12630 11560 12660
rect 11480 12590 11500 12630
rect 11540 12590 11560 12630
rect 11480 12560 11560 12590
rect 11600 12630 11680 12660
rect 11600 12590 11620 12630
rect 11660 12590 11680 12630
rect 11600 12560 11680 12590
rect 11720 12630 11800 12660
rect 11720 12590 11740 12630
rect 11780 12590 11800 12630
rect 11720 12560 11800 12590
rect 11840 12630 11920 12660
rect 11840 12590 11860 12630
rect 11900 12590 11920 12630
rect 11840 12560 11920 12590
rect 11960 12630 12040 12660
rect 11960 12590 11980 12630
rect 12020 12590 12040 12630
rect 11960 12560 12040 12590
rect 12080 12630 12160 12660
rect 12080 12590 12100 12630
rect 12140 12590 12160 12630
rect 12080 12560 12160 12590
rect 12200 12630 12280 12660
rect 12200 12590 12220 12630
rect 12260 12590 12280 12630
rect 12200 12560 12280 12590
rect 12320 12630 12400 12660
rect 12320 12590 12340 12630
rect 12380 12590 12400 12630
rect 12320 12560 12400 12590
rect 12440 12630 12520 12660
rect 12440 12590 12460 12630
rect 12500 12590 12520 12630
rect 12440 12560 12520 12590
rect 12560 12630 12640 12660
rect 12560 12590 12580 12630
rect 12620 12590 12640 12630
rect 12560 12560 12640 12590
rect 13920 12630 14000 12660
rect 13920 12590 13940 12630
rect 13980 12590 14000 12630
rect 13920 12560 14000 12590
rect 14040 12630 14120 12660
rect 14040 12590 14060 12630
rect 14100 12590 14120 12630
rect 14040 12560 14120 12590
rect 14160 12630 14240 12660
rect 14160 12590 14180 12630
rect 14220 12590 14240 12630
rect 14160 12560 14240 12590
rect 14280 12630 14360 12660
rect 14280 12590 14300 12630
rect 14340 12590 14360 12630
rect 14280 12560 14360 12590
rect 14400 12630 14480 12660
rect 14400 12590 14420 12630
rect 14460 12590 14480 12630
rect 14400 12560 14480 12590
rect 14520 12630 14600 12660
rect 14520 12590 14540 12630
rect 14580 12590 14600 12630
rect 14520 12560 14600 12590
rect 14640 12630 14720 12660
rect 14640 12590 14660 12630
rect 14700 12590 14720 12630
rect 14640 12560 14720 12590
rect 14760 12630 14840 12660
rect 14760 12590 14780 12630
rect 14820 12590 14840 12630
rect 14760 12560 14840 12590
rect 14880 12630 14960 12660
rect 14880 12590 14900 12630
rect 14940 12590 14960 12630
rect 14880 12560 14960 12590
rect 15000 12630 15080 12660
rect 15000 12590 15020 12630
rect 15060 12590 15080 12630
rect 15000 12560 15080 12590
rect 15120 12630 15200 12660
rect 15120 12590 15140 12630
rect 15180 12590 15200 12630
rect 15120 12560 15200 12590
<< pdiff >>
rect 11580 18426 12260 18480
rect 11580 18392 11632 18426
rect 11666 18392 11722 18426
rect 11756 18392 11812 18426
rect 11846 18392 11902 18426
rect 11936 18392 11992 18426
rect 12026 18392 12082 18426
rect 12116 18392 12172 18426
rect 12206 18392 12260 18426
rect 11580 18336 12260 18392
rect 11580 18302 11632 18336
rect 11666 18302 11722 18336
rect 11756 18302 11812 18336
rect 11846 18302 11902 18336
rect 11936 18302 11992 18336
rect 12026 18302 12082 18336
rect 12116 18302 12172 18336
rect 12206 18302 12260 18336
rect 11580 18246 12260 18302
rect 11580 18212 11632 18246
rect 11666 18212 11722 18246
rect 11756 18212 11812 18246
rect 11846 18212 11902 18246
rect 11936 18212 11992 18246
rect 12026 18212 12082 18246
rect 12116 18212 12172 18246
rect 12206 18212 12260 18246
rect 11580 18156 12260 18212
rect 11580 18122 11632 18156
rect 11666 18122 11722 18156
rect 11756 18122 11812 18156
rect 11846 18122 11902 18156
rect 11936 18122 11992 18156
rect 12026 18122 12082 18156
rect 12116 18122 12172 18156
rect 12206 18122 12260 18156
rect 11580 18066 12260 18122
rect 11580 18032 11632 18066
rect 11666 18032 11722 18066
rect 11756 18032 11812 18066
rect 11846 18032 11902 18066
rect 11936 18032 11992 18066
rect 12026 18032 12082 18066
rect 12116 18032 12172 18066
rect 12206 18032 12260 18066
rect 11580 17976 12260 18032
rect 11580 17942 11632 17976
rect 11666 17942 11722 17976
rect 11756 17942 11812 17976
rect 11846 17942 11902 17976
rect 11936 17942 11992 17976
rect 12026 17942 12082 17976
rect 12116 17942 12172 17976
rect 12206 17942 12260 17976
rect 11580 17886 12260 17942
rect 11580 17852 11632 17886
rect 11666 17852 11722 17886
rect 11756 17852 11812 17886
rect 11846 17852 11902 17886
rect 11936 17852 11992 17886
rect 12026 17852 12082 17886
rect 12116 17852 12172 17886
rect 12206 17852 12260 17886
rect 11580 17800 12260 17852
rect 12940 18426 13620 18480
rect 12940 18392 12992 18426
rect 13026 18392 13082 18426
rect 13116 18392 13172 18426
rect 13206 18392 13262 18426
rect 13296 18392 13352 18426
rect 13386 18392 13442 18426
rect 13476 18392 13532 18426
rect 13566 18392 13620 18426
rect 12940 18336 13620 18392
rect 12940 18302 12992 18336
rect 13026 18302 13082 18336
rect 13116 18302 13172 18336
rect 13206 18302 13262 18336
rect 13296 18302 13352 18336
rect 13386 18302 13442 18336
rect 13476 18302 13532 18336
rect 13566 18302 13620 18336
rect 12940 18246 13620 18302
rect 12940 18212 12992 18246
rect 13026 18212 13082 18246
rect 13116 18212 13172 18246
rect 13206 18212 13262 18246
rect 13296 18212 13352 18246
rect 13386 18212 13442 18246
rect 13476 18212 13532 18246
rect 13566 18212 13620 18246
rect 12940 18156 13620 18212
rect 12940 18122 12992 18156
rect 13026 18122 13082 18156
rect 13116 18122 13172 18156
rect 13206 18122 13262 18156
rect 13296 18122 13352 18156
rect 13386 18122 13442 18156
rect 13476 18122 13532 18156
rect 13566 18122 13620 18156
rect 12940 18066 13620 18122
rect 12940 18032 12992 18066
rect 13026 18032 13082 18066
rect 13116 18032 13172 18066
rect 13206 18032 13262 18066
rect 13296 18032 13352 18066
rect 13386 18032 13442 18066
rect 13476 18032 13532 18066
rect 13566 18032 13620 18066
rect 12940 17976 13620 18032
rect 12940 17942 12992 17976
rect 13026 17942 13082 17976
rect 13116 17942 13172 17976
rect 13206 17942 13262 17976
rect 13296 17942 13352 17976
rect 13386 17942 13442 17976
rect 13476 17942 13532 17976
rect 13566 17942 13620 17976
rect 12940 17886 13620 17942
rect 12940 17852 12992 17886
rect 13026 17852 13082 17886
rect 13116 17852 13172 17886
rect 13206 17852 13262 17886
rect 13296 17852 13352 17886
rect 13386 17852 13442 17886
rect 13476 17852 13532 17886
rect 13566 17852 13620 17886
rect 12940 17800 13620 17852
rect 14300 18426 14980 18480
rect 14300 18392 14352 18426
rect 14386 18392 14442 18426
rect 14476 18392 14532 18426
rect 14566 18392 14622 18426
rect 14656 18392 14712 18426
rect 14746 18392 14802 18426
rect 14836 18392 14892 18426
rect 14926 18392 14980 18426
rect 14300 18336 14980 18392
rect 14300 18302 14352 18336
rect 14386 18302 14442 18336
rect 14476 18302 14532 18336
rect 14566 18302 14622 18336
rect 14656 18302 14712 18336
rect 14746 18302 14802 18336
rect 14836 18302 14892 18336
rect 14926 18302 14980 18336
rect 14300 18246 14980 18302
rect 14300 18212 14352 18246
rect 14386 18212 14442 18246
rect 14476 18212 14532 18246
rect 14566 18212 14622 18246
rect 14656 18212 14712 18246
rect 14746 18212 14802 18246
rect 14836 18212 14892 18246
rect 14926 18212 14980 18246
rect 14300 18156 14980 18212
rect 14300 18122 14352 18156
rect 14386 18122 14442 18156
rect 14476 18122 14532 18156
rect 14566 18122 14622 18156
rect 14656 18122 14712 18156
rect 14746 18122 14802 18156
rect 14836 18122 14892 18156
rect 14926 18122 14980 18156
rect 14300 18066 14980 18122
rect 14300 18032 14352 18066
rect 14386 18032 14442 18066
rect 14476 18032 14532 18066
rect 14566 18032 14622 18066
rect 14656 18032 14712 18066
rect 14746 18032 14802 18066
rect 14836 18032 14892 18066
rect 14926 18032 14980 18066
rect 14300 17976 14980 18032
rect 14300 17942 14352 17976
rect 14386 17942 14442 17976
rect 14476 17942 14532 17976
rect 14566 17942 14622 17976
rect 14656 17942 14712 17976
rect 14746 17942 14802 17976
rect 14836 17942 14892 17976
rect 14926 17942 14980 17976
rect 14300 17886 14980 17942
rect 14300 17852 14352 17886
rect 14386 17852 14442 17886
rect 14476 17852 14532 17886
rect 14566 17852 14622 17886
rect 14656 17852 14712 17886
rect 14746 17852 14802 17886
rect 14836 17852 14892 17886
rect 14926 17852 14980 17886
rect 14300 17800 14980 17852
rect 11580 17066 12260 17120
rect 11580 17032 11632 17066
rect 11666 17032 11722 17066
rect 11756 17032 11812 17066
rect 11846 17032 11902 17066
rect 11936 17032 11992 17066
rect 12026 17032 12082 17066
rect 12116 17032 12172 17066
rect 12206 17032 12260 17066
rect 11580 16976 12260 17032
rect 11580 16942 11632 16976
rect 11666 16942 11722 16976
rect 11756 16942 11812 16976
rect 11846 16942 11902 16976
rect 11936 16942 11992 16976
rect 12026 16942 12082 16976
rect 12116 16942 12172 16976
rect 12206 16942 12260 16976
rect 11580 16886 12260 16942
rect 11580 16852 11632 16886
rect 11666 16852 11722 16886
rect 11756 16852 11812 16886
rect 11846 16852 11902 16886
rect 11936 16852 11992 16886
rect 12026 16852 12082 16886
rect 12116 16852 12172 16886
rect 12206 16852 12260 16886
rect 11580 16796 12260 16852
rect 11580 16762 11632 16796
rect 11666 16762 11722 16796
rect 11756 16762 11812 16796
rect 11846 16762 11902 16796
rect 11936 16762 11992 16796
rect 12026 16762 12082 16796
rect 12116 16762 12172 16796
rect 12206 16762 12260 16796
rect 11580 16706 12260 16762
rect 11580 16672 11632 16706
rect 11666 16672 11722 16706
rect 11756 16672 11812 16706
rect 11846 16672 11902 16706
rect 11936 16672 11992 16706
rect 12026 16672 12082 16706
rect 12116 16672 12172 16706
rect 12206 16672 12260 16706
rect 11580 16616 12260 16672
rect 11580 16582 11632 16616
rect 11666 16582 11722 16616
rect 11756 16582 11812 16616
rect 11846 16582 11902 16616
rect 11936 16582 11992 16616
rect 12026 16582 12082 16616
rect 12116 16582 12172 16616
rect 12206 16582 12260 16616
rect 11580 16526 12260 16582
rect 11580 16492 11632 16526
rect 11666 16492 11722 16526
rect 11756 16492 11812 16526
rect 11846 16492 11902 16526
rect 11936 16492 11992 16526
rect 12026 16492 12082 16526
rect 12116 16492 12172 16526
rect 12206 16492 12260 16526
rect 11580 16440 12260 16492
rect 12940 17066 13620 17120
rect 12940 17032 12992 17066
rect 13026 17032 13082 17066
rect 13116 17032 13172 17066
rect 13206 17032 13262 17066
rect 13296 17032 13352 17066
rect 13386 17032 13442 17066
rect 13476 17032 13532 17066
rect 13566 17032 13620 17066
rect 12940 16976 13620 17032
rect 12940 16942 12992 16976
rect 13026 16942 13082 16976
rect 13116 16942 13172 16976
rect 13206 16942 13262 16976
rect 13296 16942 13352 16976
rect 13386 16942 13442 16976
rect 13476 16942 13532 16976
rect 13566 16942 13620 16976
rect 12940 16886 13620 16942
rect 12940 16852 12992 16886
rect 13026 16852 13082 16886
rect 13116 16852 13172 16886
rect 13206 16852 13262 16886
rect 13296 16852 13352 16886
rect 13386 16852 13442 16886
rect 13476 16852 13532 16886
rect 13566 16852 13620 16886
rect 12940 16796 13620 16852
rect 12940 16762 12992 16796
rect 13026 16762 13082 16796
rect 13116 16762 13172 16796
rect 13206 16762 13262 16796
rect 13296 16762 13352 16796
rect 13386 16762 13442 16796
rect 13476 16762 13532 16796
rect 13566 16762 13620 16796
rect 12940 16706 13620 16762
rect 12940 16672 12992 16706
rect 13026 16672 13082 16706
rect 13116 16672 13172 16706
rect 13206 16672 13262 16706
rect 13296 16672 13352 16706
rect 13386 16672 13442 16706
rect 13476 16672 13532 16706
rect 13566 16672 13620 16706
rect 12940 16616 13620 16672
rect 12940 16582 12992 16616
rect 13026 16582 13082 16616
rect 13116 16582 13172 16616
rect 13206 16582 13262 16616
rect 13296 16582 13352 16616
rect 13386 16582 13442 16616
rect 13476 16582 13532 16616
rect 13566 16582 13620 16616
rect 12940 16526 13620 16582
rect 12940 16492 12992 16526
rect 13026 16492 13082 16526
rect 13116 16492 13172 16526
rect 13206 16492 13262 16526
rect 13296 16492 13352 16526
rect 13386 16492 13442 16526
rect 13476 16492 13532 16526
rect 13566 16492 13620 16526
rect 12940 16440 13620 16492
rect 14300 17066 14980 17120
rect 14300 17032 14352 17066
rect 14386 17032 14442 17066
rect 14476 17032 14532 17066
rect 14566 17032 14622 17066
rect 14656 17032 14712 17066
rect 14746 17032 14802 17066
rect 14836 17032 14892 17066
rect 14926 17032 14980 17066
rect 14300 16976 14980 17032
rect 14300 16942 14352 16976
rect 14386 16942 14442 16976
rect 14476 16942 14532 16976
rect 14566 16942 14622 16976
rect 14656 16942 14712 16976
rect 14746 16942 14802 16976
rect 14836 16942 14892 16976
rect 14926 16942 14980 16976
rect 14300 16886 14980 16942
rect 14300 16852 14352 16886
rect 14386 16852 14442 16886
rect 14476 16852 14532 16886
rect 14566 16852 14622 16886
rect 14656 16852 14712 16886
rect 14746 16852 14802 16886
rect 14836 16852 14892 16886
rect 14926 16852 14980 16886
rect 14300 16796 14980 16852
rect 14300 16762 14352 16796
rect 14386 16762 14442 16796
rect 14476 16762 14532 16796
rect 14566 16762 14622 16796
rect 14656 16762 14712 16796
rect 14746 16762 14802 16796
rect 14836 16762 14892 16796
rect 14926 16762 14980 16796
rect 14300 16706 14980 16762
rect 14300 16672 14352 16706
rect 14386 16672 14442 16706
rect 14476 16672 14532 16706
rect 14566 16672 14622 16706
rect 14656 16672 14712 16706
rect 14746 16672 14802 16706
rect 14836 16672 14892 16706
rect 14926 16672 14980 16706
rect 14300 16616 14980 16672
rect 14300 16582 14352 16616
rect 14386 16582 14442 16616
rect 14476 16582 14532 16616
rect 14566 16582 14622 16616
rect 14656 16582 14712 16616
rect 14746 16582 14802 16616
rect 14836 16582 14892 16616
rect 14926 16582 14980 16616
rect 14300 16526 14980 16582
rect 14300 16492 14352 16526
rect 14386 16492 14442 16526
rect 14476 16492 14532 16526
rect 14566 16492 14622 16526
rect 14656 16492 14712 16526
rect 14746 16492 14802 16526
rect 14836 16492 14892 16526
rect 14926 16492 14980 16526
rect 14300 16440 14980 16492
rect 11580 15706 12260 15760
rect 11580 15672 11632 15706
rect 11666 15672 11722 15706
rect 11756 15672 11812 15706
rect 11846 15672 11902 15706
rect 11936 15672 11992 15706
rect 12026 15672 12082 15706
rect 12116 15672 12172 15706
rect 12206 15672 12260 15706
rect 11580 15616 12260 15672
rect 11580 15582 11632 15616
rect 11666 15582 11722 15616
rect 11756 15582 11812 15616
rect 11846 15582 11902 15616
rect 11936 15582 11992 15616
rect 12026 15582 12082 15616
rect 12116 15582 12172 15616
rect 12206 15582 12260 15616
rect 11580 15526 12260 15582
rect 11580 15492 11632 15526
rect 11666 15492 11722 15526
rect 11756 15492 11812 15526
rect 11846 15492 11902 15526
rect 11936 15492 11992 15526
rect 12026 15492 12082 15526
rect 12116 15492 12172 15526
rect 12206 15492 12260 15526
rect 11580 15436 12260 15492
rect 11580 15402 11632 15436
rect 11666 15402 11722 15436
rect 11756 15402 11812 15436
rect 11846 15402 11902 15436
rect 11936 15402 11992 15436
rect 12026 15402 12082 15436
rect 12116 15402 12172 15436
rect 12206 15402 12260 15436
rect 11580 15346 12260 15402
rect 11580 15312 11632 15346
rect 11666 15312 11722 15346
rect 11756 15312 11812 15346
rect 11846 15312 11902 15346
rect 11936 15312 11992 15346
rect 12026 15312 12082 15346
rect 12116 15312 12172 15346
rect 12206 15312 12260 15346
rect 11580 15256 12260 15312
rect 11580 15222 11632 15256
rect 11666 15222 11722 15256
rect 11756 15222 11812 15256
rect 11846 15222 11902 15256
rect 11936 15222 11992 15256
rect 12026 15222 12082 15256
rect 12116 15222 12172 15256
rect 12206 15222 12260 15256
rect 11580 15166 12260 15222
rect 11580 15132 11632 15166
rect 11666 15132 11722 15166
rect 11756 15132 11812 15166
rect 11846 15132 11902 15166
rect 11936 15132 11992 15166
rect 12026 15132 12082 15166
rect 12116 15132 12172 15166
rect 12206 15132 12260 15166
rect 11580 15080 12260 15132
rect 12940 15706 13620 15760
rect 12940 15672 12992 15706
rect 13026 15672 13082 15706
rect 13116 15672 13172 15706
rect 13206 15672 13262 15706
rect 13296 15672 13352 15706
rect 13386 15672 13442 15706
rect 13476 15672 13532 15706
rect 13566 15672 13620 15706
rect 12940 15616 13620 15672
rect 12940 15582 12992 15616
rect 13026 15582 13082 15616
rect 13116 15582 13172 15616
rect 13206 15582 13262 15616
rect 13296 15582 13352 15616
rect 13386 15582 13442 15616
rect 13476 15582 13532 15616
rect 13566 15582 13620 15616
rect 12940 15526 13620 15582
rect 12940 15492 12992 15526
rect 13026 15492 13082 15526
rect 13116 15492 13172 15526
rect 13206 15492 13262 15526
rect 13296 15492 13352 15526
rect 13386 15492 13442 15526
rect 13476 15492 13532 15526
rect 13566 15492 13620 15526
rect 12940 15436 13620 15492
rect 12940 15402 12992 15436
rect 13026 15402 13082 15436
rect 13116 15402 13172 15436
rect 13206 15402 13262 15436
rect 13296 15402 13352 15436
rect 13386 15402 13442 15436
rect 13476 15402 13532 15436
rect 13566 15402 13620 15436
rect 12940 15346 13620 15402
rect 12940 15312 12992 15346
rect 13026 15312 13082 15346
rect 13116 15312 13172 15346
rect 13206 15312 13262 15346
rect 13296 15312 13352 15346
rect 13386 15312 13442 15346
rect 13476 15312 13532 15346
rect 13566 15312 13620 15346
rect 12940 15256 13620 15312
rect 12940 15222 12992 15256
rect 13026 15222 13082 15256
rect 13116 15222 13172 15256
rect 13206 15222 13262 15256
rect 13296 15222 13352 15256
rect 13386 15222 13442 15256
rect 13476 15222 13532 15256
rect 13566 15222 13620 15256
rect 12940 15166 13620 15222
rect 12940 15132 12992 15166
rect 13026 15132 13082 15166
rect 13116 15132 13172 15166
rect 13206 15132 13262 15166
rect 13296 15132 13352 15166
rect 13386 15132 13442 15166
rect 13476 15132 13532 15166
rect 13566 15132 13620 15166
rect 12940 15080 13620 15132
rect 14300 15706 14980 15760
rect 14300 15672 14352 15706
rect 14386 15672 14442 15706
rect 14476 15672 14532 15706
rect 14566 15672 14622 15706
rect 14656 15672 14712 15706
rect 14746 15672 14802 15706
rect 14836 15672 14892 15706
rect 14926 15672 14980 15706
rect 14300 15616 14980 15672
rect 14300 15582 14352 15616
rect 14386 15582 14442 15616
rect 14476 15582 14532 15616
rect 14566 15582 14622 15616
rect 14656 15582 14712 15616
rect 14746 15582 14802 15616
rect 14836 15582 14892 15616
rect 14926 15582 14980 15616
rect 14300 15526 14980 15582
rect 14300 15492 14352 15526
rect 14386 15492 14442 15526
rect 14476 15492 14532 15526
rect 14566 15492 14622 15526
rect 14656 15492 14712 15526
rect 14746 15492 14802 15526
rect 14836 15492 14892 15526
rect 14926 15492 14980 15526
rect 14300 15436 14980 15492
rect 14300 15402 14352 15436
rect 14386 15402 14442 15436
rect 14476 15402 14532 15436
rect 14566 15402 14622 15436
rect 14656 15402 14712 15436
rect 14746 15402 14802 15436
rect 14836 15402 14892 15436
rect 14926 15402 14980 15436
rect 14300 15346 14980 15402
rect 14300 15312 14352 15346
rect 14386 15312 14442 15346
rect 14476 15312 14532 15346
rect 14566 15312 14622 15346
rect 14656 15312 14712 15346
rect 14746 15312 14802 15346
rect 14836 15312 14892 15346
rect 14926 15312 14980 15346
rect 14300 15256 14980 15312
rect 14300 15222 14352 15256
rect 14386 15222 14442 15256
rect 14476 15222 14532 15256
rect 14566 15222 14622 15256
rect 14656 15222 14712 15256
rect 14746 15222 14802 15256
rect 14836 15222 14892 15256
rect 14926 15222 14980 15256
rect 14300 15166 14980 15222
rect 14300 15132 14352 15166
rect 14386 15132 14442 15166
rect 14476 15132 14532 15166
rect 14566 15132 14622 15166
rect 14656 15132 14712 15166
rect 14746 15132 14802 15166
rect 14836 15132 14892 15166
rect 14926 15132 14980 15166
rect 14300 15080 14980 15132
rect 10520 11790 10600 11820
rect 10520 11750 10540 11790
rect 10580 11750 10600 11790
rect 10520 11690 10600 11750
rect 10520 11650 10540 11690
rect 10580 11650 10600 11690
rect 10520 11620 10600 11650
rect 10640 11790 10720 11820
rect 10640 11750 10660 11790
rect 10700 11750 10720 11790
rect 10640 11690 10720 11750
rect 10640 11650 10660 11690
rect 10700 11650 10720 11690
rect 10640 11620 10720 11650
rect 10760 11790 10840 11820
rect 10760 11750 10780 11790
rect 10820 11750 10840 11790
rect 10760 11690 10840 11750
rect 10760 11650 10780 11690
rect 10820 11650 10840 11690
rect 10760 11620 10840 11650
rect 10880 11790 10960 11820
rect 10880 11750 10900 11790
rect 10940 11750 10960 11790
rect 10880 11690 10960 11750
rect 10880 11650 10900 11690
rect 10940 11650 10960 11690
rect 10880 11620 10960 11650
rect 11000 11790 11080 11820
rect 11000 11750 11020 11790
rect 11060 11750 11080 11790
rect 11000 11690 11080 11750
rect 11000 11650 11020 11690
rect 11060 11650 11080 11690
rect 11000 11620 11080 11650
rect 11120 11790 11200 11820
rect 11120 11750 11140 11790
rect 11180 11750 11200 11790
rect 11120 11690 11200 11750
rect 11120 11650 11140 11690
rect 11180 11650 11200 11690
rect 11120 11620 11200 11650
rect 11240 11790 11320 11820
rect 11240 11750 11260 11790
rect 11300 11750 11320 11790
rect 11240 11690 11320 11750
rect 11240 11650 11260 11690
rect 11300 11650 11320 11690
rect 11240 11620 11320 11650
rect 11360 11790 11440 11820
rect 11360 11750 11380 11790
rect 11420 11750 11440 11790
rect 11360 11690 11440 11750
rect 11360 11650 11380 11690
rect 11420 11650 11440 11690
rect 11360 11620 11440 11650
rect 11480 11790 11560 11820
rect 11480 11750 11500 11790
rect 11540 11750 11560 11790
rect 11480 11690 11560 11750
rect 11480 11650 11500 11690
rect 11540 11650 11560 11690
rect 11480 11620 11560 11650
rect 11600 11790 11680 11820
rect 11600 11750 11620 11790
rect 11660 11750 11680 11790
rect 11600 11690 11680 11750
rect 11600 11650 11620 11690
rect 11660 11650 11680 11690
rect 11600 11620 11680 11650
rect 11720 11790 11800 11820
rect 11720 11750 11740 11790
rect 11780 11750 11800 11790
rect 11720 11690 11800 11750
rect 11720 11650 11740 11690
rect 11780 11650 11800 11690
rect 11720 11620 11800 11650
rect 11840 11790 11920 11820
rect 11840 11750 11860 11790
rect 11900 11750 11920 11790
rect 11840 11690 11920 11750
rect 11840 11650 11860 11690
rect 11900 11650 11920 11690
rect 11840 11620 11920 11650
rect 11960 11790 12040 11820
rect 11960 11750 11980 11790
rect 12020 11750 12040 11790
rect 11960 11690 12040 11750
rect 11960 11650 11980 11690
rect 12020 11650 12040 11690
rect 11960 11620 12040 11650
rect 12080 11790 12160 11820
rect 12080 11750 12100 11790
rect 12140 11750 12160 11790
rect 12080 11690 12160 11750
rect 12080 11650 12100 11690
rect 12140 11650 12160 11690
rect 12080 11620 12160 11650
rect 12200 11790 12280 11820
rect 12200 11750 12220 11790
rect 12260 11750 12280 11790
rect 12200 11690 12280 11750
rect 12200 11650 12220 11690
rect 12260 11650 12280 11690
rect 12200 11620 12280 11650
rect 12320 11790 12400 11820
rect 12320 11750 12340 11790
rect 12380 11750 12400 11790
rect 12320 11690 12400 11750
rect 12320 11650 12340 11690
rect 12380 11650 12400 11690
rect 12320 11620 12400 11650
rect 12440 11790 12520 11820
rect 12440 11750 12460 11790
rect 12500 11750 12520 11790
rect 12440 11690 12520 11750
rect 12440 11650 12460 11690
rect 12500 11650 12520 11690
rect 12440 11620 12520 11650
rect 12560 11790 12640 11820
rect 12560 11750 12580 11790
rect 12620 11750 12640 11790
rect 12560 11690 12640 11750
rect 12560 11650 12580 11690
rect 12620 11650 12640 11690
rect 12560 11620 12640 11650
rect 12680 11790 12760 11820
rect 12680 11750 12700 11790
rect 12740 11750 12760 11790
rect 12680 11690 12760 11750
rect 12680 11650 12700 11690
rect 12740 11650 12760 11690
rect 12680 11620 12760 11650
rect 12800 11790 12880 11820
rect 12800 11750 12820 11790
rect 12860 11750 12880 11790
rect 12800 11690 12880 11750
rect 12800 11650 12820 11690
rect 12860 11650 12880 11690
rect 12800 11620 12880 11650
rect 12920 11790 13000 11820
rect 12920 11750 12940 11790
rect 12980 11750 13000 11790
rect 12920 11690 13000 11750
rect 12920 11650 12940 11690
rect 12980 11650 13000 11690
rect 12920 11620 13000 11650
rect 13560 11790 13640 11820
rect 13560 11750 13580 11790
rect 13620 11750 13640 11790
rect 13560 11690 13640 11750
rect 13560 11650 13580 11690
rect 13620 11650 13640 11690
rect 13560 11620 13640 11650
rect 13680 11790 13760 11820
rect 13680 11750 13700 11790
rect 13740 11750 13760 11790
rect 13680 11690 13760 11750
rect 13680 11650 13700 11690
rect 13740 11650 13760 11690
rect 13680 11620 13760 11650
rect 13800 11790 13880 11820
rect 13800 11750 13820 11790
rect 13860 11750 13880 11790
rect 13800 11690 13880 11750
rect 13800 11650 13820 11690
rect 13860 11650 13880 11690
rect 13800 11620 13880 11650
rect 13920 11790 14000 11820
rect 13920 11750 13940 11790
rect 13980 11750 14000 11790
rect 13920 11690 14000 11750
rect 13920 11650 13940 11690
rect 13980 11650 14000 11690
rect 13920 11620 14000 11650
rect 14040 11790 14120 11820
rect 14040 11750 14060 11790
rect 14100 11750 14120 11790
rect 14040 11690 14120 11750
rect 14040 11650 14060 11690
rect 14100 11650 14120 11690
rect 14040 11620 14120 11650
rect 14160 11790 14240 11820
rect 14160 11750 14180 11790
rect 14220 11750 14240 11790
rect 14160 11690 14240 11750
rect 14160 11650 14180 11690
rect 14220 11650 14240 11690
rect 14160 11620 14240 11650
rect 14280 11790 14360 11820
rect 14280 11750 14300 11790
rect 14340 11750 14360 11790
rect 14280 11690 14360 11750
rect 14280 11650 14300 11690
rect 14340 11650 14360 11690
rect 14280 11620 14360 11650
rect 14400 11790 14480 11820
rect 14400 11750 14420 11790
rect 14460 11750 14480 11790
rect 14400 11690 14480 11750
rect 14400 11650 14420 11690
rect 14460 11650 14480 11690
rect 14400 11620 14480 11650
rect 14520 11790 14600 11820
rect 14520 11750 14540 11790
rect 14580 11750 14600 11790
rect 14520 11690 14600 11750
rect 14520 11650 14540 11690
rect 14580 11650 14600 11690
rect 14520 11620 14600 11650
rect 14640 11790 14720 11820
rect 14640 11750 14660 11790
rect 14700 11750 14720 11790
rect 14640 11690 14720 11750
rect 14640 11650 14660 11690
rect 14700 11650 14720 11690
rect 14640 11620 14720 11650
rect 14760 11790 14840 11820
rect 14760 11750 14780 11790
rect 14820 11750 14840 11790
rect 14760 11690 14840 11750
rect 14760 11650 14780 11690
rect 14820 11650 14840 11690
rect 14760 11620 14840 11650
rect 14880 11790 14960 11820
rect 14880 11750 14900 11790
rect 14940 11750 14960 11790
rect 14880 11690 14960 11750
rect 14880 11650 14900 11690
rect 14940 11650 14960 11690
rect 14880 11620 14960 11650
rect 15000 11790 15080 11820
rect 15000 11750 15020 11790
rect 15060 11750 15080 11790
rect 15000 11690 15080 11750
rect 15000 11650 15020 11690
rect 15060 11650 15080 11690
rect 15000 11620 15080 11650
rect 15120 11790 15200 11820
rect 15120 11750 15140 11790
rect 15180 11750 15200 11790
rect 15120 11690 15200 11750
rect 15120 11650 15140 11690
rect 15180 11650 15200 11690
rect 15120 11620 15200 11650
rect 15240 11790 15320 11820
rect 15240 11750 15260 11790
rect 15300 11750 15320 11790
rect 15240 11690 15320 11750
rect 15240 11650 15260 11690
rect 15300 11650 15320 11690
rect 15240 11620 15320 11650
rect 15360 11790 15440 11820
rect 15360 11750 15380 11790
rect 15420 11750 15440 11790
rect 15360 11690 15440 11750
rect 15360 11650 15380 11690
rect 15420 11650 15440 11690
rect 15360 11620 15440 11650
rect 15480 11790 15560 11820
rect 15480 11750 15500 11790
rect 15540 11750 15560 11790
rect 15480 11690 15560 11750
rect 15480 11650 15500 11690
rect 15540 11650 15560 11690
rect 15480 11620 15560 11650
rect 15600 11790 15680 11820
rect 15600 11750 15620 11790
rect 15660 11750 15680 11790
rect 15600 11690 15680 11750
rect 15600 11650 15620 11690
rect 15660 11650 15680 11690
rect 15600 11620 15680 11650
rect 15720 11790 15800 11820
rect 15720 11750 15740 11790
rect 15780 11750 15800 11790
rect 15720 11690 15800 11750
rect 15720 11650 15740 11690
rect 15780 11650 15800 11690
rect 15720 11620 15800 11650
rect 15840 11790 15920 11820
rect 15840 11750 15860 11790
rect 15900 11750 15920 11790
rect 15840 11690 15920 11750
rect 15840 11650 15860 11690
rect 15900 11650 15920 11690
rect 15840 11620 15920 11650
rect 15960 11790 16040 11820
rect 15960 11750 15980 11790
rect 16020 11750 16040 11790
rect 15960 11690 16040 11750
rect 15960 11650 15980 11690
rect 16020 11650 16040 11690
rect 15960 11620 16040 11650
rect 11620 10630 11700 10660
rect 11620 10590 11640 10630
rect 11680 10590 11700 10630
rect 11620 10530 11700 10590
rect 11620 10490 11640 10530
rect 11680 10490 11700 10530
rect 11620 10430 11700 10490
rect 11620 10390 11640 10430
rect 11680 10390 11700 10430
rect 11620 10330 11700 10390
rect 11620 10290 11640 10330
rect 11680 10290 11700 10330
rect 11620 10230 11700 10290
rect 11620 10190 11640 10230
rect 11680 10190 11700 10230
rect 11620 10130 11700 10190
rect 11620 10090 11640 10130
rect 11680 10090 11700 10130
rect 11620 10060 11700 10090
rect 11800 10630 11880 10660
rect 11800 10590 11820 10630
rect 11860 10590 11880 10630
rect 11800 10530 11880 10590
rect 11800 10490 11820 10530
rect 11860 10490 11880 10530
rect 11800 10430 11880 10490
rect 11800 10390 11820 10430
rect 11860 10390 11880 10430
rect 11800 10330 11880 10390
rect 11800 10290 11820 10330
rect 11860 10290 11880 10330
rect 11800 10230 11880 10290
rect 11800 10190 11820 10230
rect 11860 10190 11880 10230
rect 11800 10130 11880 10190
rect 11800 10090 11820 10130
rect 11860 10090 11880 10130
rect 11800 10060 11880 10090
rect 11980 10630 12060 10660
rect 11980 10590 12000 10630
rect 12040 10590 12060 10630
rect 11980 10530 12060 10590
rect 11980 10490 12000 10530
rect 12040 10490 12060 10530
rect 11980 10430 12060 10490
rect 11980 10390 12000 10430
rect 12040 10390 12060 10430
rect 11980 10330 12060 10390
rect 11980 10290 12000 10330
rect 12040 10290 12060 10330
rect 11980 10230 12060 10290
rect 11980 10190 12000 10230
rect 12040 10190 12060 10230
rect 11980 10130 12060 10190
rect 11980 10090 12000 10130
rect 12040 10090 12060 10130
rect 11980 10060 12060 10090
rect 12160 10630 12240 10660
rect 12160 10590 12180 10630
rect 12220 10590 12240 10630
rect 12160 10530 12240 10590
rect 12160 10490 12180 10530
rect 12220 10490 12240 10530
rect 12160 10430 12240 10490
rect 12160 10390 12180 10430
rect 12220 10390 12240 10430
rect 12160 10330 12240 10390
rect 12160 10290 12180 10330
rect 12220 10290 12240 10330
rect 12160 10230 12240 10290
rect 12160 10190 12180 10230
rect 12220 10190 12240 10230
rect 12160 10130 12240 10190
rect 12160 10090 12180 10130
rect 12220 10090 12240 10130
rect 12160 10060 12240 10090
rect 12340 10630 12420 10660
rect 12340 10590 12360 10630
rect 12400 10590 12420 10630
rect 12340 10530 12420 10590
rect 12340 10490 12360 10530
rect 12400 10490 12420 10530
rect 12340 10430 12420 10490
rect 12340 10390 12360 10430
rect 12400 10390 12420 10430
rect 12340 10330 12420 10390
rect 12340 10290 12360 10330
rect 12400 10290 12420 10330
rect 12340 10230 12420 10290
rect 12340 10190 12360 10230
rect 12400 10190 12420 10230
rect 12340 10130 12420 10190
rect 12340 10090 12360 10130
rect 12400 10090 12420 10130
rect 12340 10060 12420 10090
rect 12520 10630 12600 10660
rect 12520 10590 12540 10630
rect 12580 10590 12600 10630
rect 12520 10530 12600 10590
rect 12520 10490 12540 10530
rect 12580 10490 12600 10530
rect 12520 10430 12600 10490
rect 12520 10390 12540 10430
rect 12580 10390 12600 10430
rect 12520 10330 12600 10390
rect 12520 10290 12540 10330
rect 12580 10290 12600 10330
rect 12520 10230 12600 10290
rect 12520 10190 12540 10230
rect 12580 10190 12600 10230
rect 12520 10130 12600 10190
rect 12520 10090 12540 10130
rect 12580 10090 12600 10130
rect 12520 10060 12600 10090
rect 12700 10630 12780 10660
rect 12700 10590 12720 10630
rect 12760 10590 12780 10630
rect 12700 10530 12780 10590
rect 12700 10490 12720 10530
rect 12760 10490 12780 10530
rect 12700 10430 12780 10490
rect 12700 10390 12720 10430
rect 12760 10390 12780 10430
rect 12700 10330 12780 10390
rect 12700 10290 12720 10330
rect 12760 10290 12780 10330
rect 12700 10230 12780 10290
rect 12700 10190 12720 10230
rect 12760 10190 12780 10230
rect 12700 10130 12780 10190
rect 12700 10090 12720 10130
rect 12760 10090 12780 10130
rect 12700 10060 12780 10090
rect 12880 10630 12960 10660
rect 12880 10590 12900 10630
rect 12940 10590 12960 10630
rect 12880 10530 12960 10590
rect 12880 10490 12900 10530
rect 12940 10490 12960 10530
rect 12880 10430 12960 10490
rect 12880 10390 12900 10430
rect 12940 10390 12960 10430
rect 12880 10330 12960 10390
rect 12880 10290 12900 10330
rect 12940 10290 12960 10330
rect 12880 10230 12960 10290
rect 12880 10190 12900 10230
rect 12940 10190 12960 10230
rect 12880 10130 12960 10190
rect 12880 10090 12900 10130
rect 12940 10090 12960 10130
rect 12880 10060 12960 10090
rect 13060 10630 13140 10660
rect 13060 10590 13080 10630
rect 13120 10590 13140 10630
rect 13060 10530 13140 10590
rect 13060 10490 13080 10530
rect 13120 10490 13140 10530
rect 13060 10430 13140 10490
rect 13060 10390 13080 10430
rect 13120 10390 13140 10430
rect 13060 10330 13140 10390
rect 13060 10290 13080 10330
rect 13120 10290 13140 10330
rect 13060 10230 13140 10290
rect 13060 10190 13080 10230
rect 13120 10190 13140 10230
rect 13060 10130 13140 10190
rect 13060 10090 13080 10130
rect 13120 10090 13140 10130
rect 13060 10060 13140 10090
rect 13240 10630 13320 10660
rect 13240 10590 13260 10630
rect 13300 10590 13320 10630
rect 13240 10530 13320 10590
rect 13240 10490 13260 10530
rect 13300 10490 13320 10530
rect 13240 10430 13320 10490
rect 13240 10390 13260 10430
rect 13300 10390 13320 10430
rect 13240 10330 13320 10390
rect 13240 10290 13260 10330
rect 13300 10290 13320 10330
rect 13240 10230 13320 10290
rect 13240 10190 13260 10230
rect 13300 10190 13320 10230
rect 13240 10130 13320 10190
rect 13240 10090 13260 10130
rect 13300 10090 13320 10130
rect 13240 10060 13320 10090
rect 13420 10630 13500 10660
rect 13420 10590 13440 10630
rect 13480 10590 13500 10630
rect 13420 10530 13500 10590
rect 13420 10490 13440 10530
rect 13480 10490 13500 10530
rect 13420 10430 13500 10490
rect 13420 10390 13440 10430
rect 13480 10390 13500 10430
rect 13420 10330 13500 10390
rect 13420 10290 13440 10330
rect 13480 10290 13500 10330
rect 13420 10230 13500 10290
rect 13420 10190 13440 10230
rect 13480 10190 13500 10230
rect 13420 10130 13500 10190
rect 13420 10090 13440 10130
rect 13480 10090 13500 10130
rect 13420 10060 13500 10090
rect 13600 10630 13680 10660
rect 13600 10590 13620 10630
rect 13660 10590 13680 10630
rect 13600 10530 13680 10590
rect 13600 10490 13620 10530
rect 13660 10490 13680 10530
rect 13600 10430 13680 10490
rect 13600 10390 13620 10430
rect 13660 10390 13680 10430
rect 13600 10330 13680 10390
rect 13600 10290 13620 10330
rect 13660 10290 13680 10330
rect 13600 10230 13680 10290
rect 13600 10190 13620 10230
rect 13660 10190 13680 10230
rect 13600 10130 13680 10190
rect 13600 10090 13620 10130
rect 13660 10090 13680 10130
rect 13600 10060 13680 10090
rect 13780 10630 13860 10660
rect 13780 10590 13800 10630
rect 13840 10590 13860 10630
rect 13780 10530 13860 10590
rect 13780 10490 13800 10530
rect 13840 10490 13860 10530
rect 13780 10430 13860 10490
rect 13780 10390 13800 10430
rect 13840 10390 13860 10430
rect 13780 10330 13860 10390
rect 13780 10290 13800 10330
rect 13840 10290 13860 10330
rect 13780 10230 13860 10290
rect 13780 10190 13800 10230
rect 13840 10190 13860 10230
rect 13780 10130 13860 10190
rect 13780 10090 13800 10130
rect 13840 10090 13860 10130
rect 13780 10060 13860 10090
rect 13960 10630 14040 10660
rect 13960 10590 13980 10630
rect 14020 10590 14040 10630
rect 13960 10530 14040 10590
rect 13960 10490 13980 10530
rect 14020 10490 14040 10530
rect 13960 10430 14040 10490
rect 13960 10390 13980 10430
rect 14020 10390 14040 10430
rect 13960 10330 14040 10390
rect 13960 10290 13980 10330
rect 14020 10290 14040 10330
rect 13960 10230 14040 10290
rect 13960 10190 13980 10230
rect 14020 10190 14040 10230
rect 13960 10130 14040 10190
rect 13960 10090 13980 10130
rect 14020 10090 14040 10130
rect 13960 10060 14040 10090
rect 14140 10630 14220 10660
rect 14140 10590 14160 10630
rect 14200 10590 14220 10630
rect 14140 10530 14220 10590
rect 14140 10490 14160 10530
rect 14200 10490 14220 10530
rect 14140 10430 14220 10490
rect 14140 10390 14160 10430
rect 14200 10390 14220 10430
rect 14140 10330 14220 10390
rect 14140 10290 14160 10330
rect 14200 10290 14220 10330
rect 14140 10230 14220 10290
rect 14140 10190 14160 10230
rect 14200 10190 14220 10230
rect 14140 10130 14220 10190
rect 14140 10090 14160 10130
rect 14200 10090 14220 10130
rect 14140 10060 14220 10090
rect 14320 10630 14400 10660
rect 14320 10590 14340 10630
rect 14380 10590 14400 10630
rect 14320 10530 14400 10590
rect 14320 10490 14340 10530
rect 14380 10490 14400 10530
rect 14320 10430 14400 10490
rect 14320 10390 14340 10430
rect 14380 10390 14400 10430
rect 14320 10330 14400 10390
rect 14320 10290 14340 10330
rect 14380 10290 14400 10330
rect 14320 10230 14400 10290
rect 14320 10190 14340 10230
rect 14380 10190 14400 10230
rect 14320 10130 14400 10190
rect 14320 10090 14340 10130
rect 14380 10090 14400 10130
rect 14320 10060 14400 10090
rect 14500 10630 14580 10660
rect 14500 10590 14520 10630
rect 14560 10590 14580 10630
rect 14500 10530 14580 10590
rect 14500 10490 14520 10530
rect 14560 10490 14580 10530
rect 14500 10430 14580 10490
rect 14500 10390 14520 10430
rect 14560 10390 14580 10430
rect 14500 10330 14580 10390
rect 14500 10290 14520 10330
rect 14560 10290 14580 10330
rect 14500 10230 14580 10290
rect 14500 10190 14520 10230
rect 14560 10190 14580 10230
rect 14500 10130 14580 10190
rect 14500 10090 14520 10130
rect 14560 10090 14580 10130
rect 14500 10060 14580 10090
rect 14680 10630 14760 10660
rect 14680 10590 14700 10630
rect 14740 10590 14760 10630
rect 14680 10530 14760 10590
rect 14680 10490 14700 10530
rect 14740 10490 14760 10530
rect 14680 10430 14760 10490
rect 14680 10390 14700 10430
rect 14740 10390 14760 10430
rect 14680 10330 14760 10390
rect 14680 10290 14700 10330
rect 14740 10290 14760 10330
rect 14680 10230 14760 10290
rect 14680 10190 14700 10230
rect 14740 10190 14760 10230
rect 14680 10130 14760 10190
rect 14680 10090 14700 10130
rect 14740 10090 14760 10130
rect 14680 10060 14760 10090
rect 14860 10630 14940 10660
rect 14860 10590 14880 10630
rect 14920 10590 14940 10630
rect 14860 10530 14940 10590
rect 14860 10490 14880 10530
rect 14920 10490 14940 10530
rect 14860 10430 14940 10490
rect 14860 10390 14880 10430
rect 14920 10390 14940 10430
rect 14860 10330 14940 10390
rect 14860 10290 14880 10330
rect 14920 10290 14940 10330
rect 14860 10230 14940 10290
rect 15480 10430 15570 10460
rect 15480 10390 15510 10430
rect 15550 10390 15570 10430
rect 15480 10330 15570 10390
rect 15480 10290 15510 10330
rect 15550 10290 15570 10330
rect 15480 10260 15570 10290
rect 15600 10430 15680 10460
rect 15600 10390 15620 10430
rect 15660 10390 15680 10430
rect 15600 10330 15680 10390
rect 15600 10290 15620 10330
rect 15660 10290 15680 10330
rect 15600 10260 15680 10290
rect 15710 10430 15790 10460
rect 15710 10390 15730 10430
rect 15770 10390 15790 10430
rect 15710 10330 15790 10390
rect 15710 10290 15730 10330
rect 15770 10290 15790 10330
rect 15710 10260 15790 10290
rect 15820 10430 15900 10460
rect 15820 10390 15840 10430
rect 15880 10390 15900 10430
rect 15820 10330 15900 10390
rect 15820 10290 15840 10330
rect 15880 10290 15900 10330
rect 15820 10260 15900 10290
rect 15930 10430 16010 10460
rect 15930 10390 15950 10430
rect 15990 10390 16010 10430
rect 15930 10330 16010 10390
rect 15930 10290 15950 10330
rect 15990 10290 16010 10330
rect 15930 10260 16010 10290
rect 14860 10190 14880 10230
rect 14920 10190 14940 10230
rect 14860 10130 14940 10190
rect 14860 10090 14880 10130
rect 14920 10090 14940 10130
rect 14860 10060 14940 10090
rect 11630 9630 11710 9660
rect 11630 9590 11650 9630
rect 11690 9590 11710 9630
rect 11630 9530 11710 9590
rect 11630 9490 11650 9530
rect 11690 9490 11710 9530
rect 11630 9460 11710 9490
rect 11740 9630 11820 9660
rect 11740 9590 11760 9630
rect 11800 9590 11820 9630
rect 11740 9530 11820 9590
rect 11740 9490 11760 9530
rect 11800 9490 11820 9530
rect 11740 9460 11820 9490
rect 11850 9630 11930 9660
rect 11850 9590 11870 9630
rect 11910 9590 11930 9630
rect 11850 9530 11930 9590
rect 11850 9490 11870 9530
rect 11910 9490 11930 9530
rect 11850 9460 11930 9490
rect 11960 9630 12040 9660
rect 11960 9590 11980 9630
rect 12020 9590 12040 9630
rect 11960 9530 12040 9590
rect 11960 9490 11980 9530
rect 12020 9490 12040 9530
rect 11960 9460 12040 9490
rect 12070 9630 12150 9660
rect 12070 9590 12090 9630
rect 12130 9590 12150 9630
rect 12070 9530 12150 9590
rect 12070 9490 12090 9530
rect 12130 9490 12150 9530
rect 12070 9460 12150 9490
rect 12180 9630 12260 9660
rect 12180 9590 12200 9630
rect 12240 9590 12260 9630
rect 12180 9530 12260 9590
rect 12180 9490 12200 9530
rect 12240 9490 12260 9530
rect 12180 9460 12260 9490
rect 12290 9630 12370 9660
rect 12290 9590 12310 9630
rect 12350 9590 12370 9630
rect 12290 9530 12370 9590
rect 12290 9490 12310 9530
rect 12350 9490 12370 9530
rect 12290 9460 12370 9490
rect 12400 9630 12480 9660
rect 12400 9590 12420 9630
rect 12460 9590 12480 9630
rect 12400 9530 12480 9590
rect 12400 9490 12420 9530
rect 12460 9490 12480 9530
rect 12400 9460 12480 9490
rect 12510 9630 12590 9660
rect 12510 9590 12530 9630
rect 12570 9590 12590 9630
rect 12510 9530 12590 9590
rect 12510 9490 12530 9530
rect 12570 9490 12590 9530
rect 12510 9460 12590 9490
rect 12620 9630 12700 9660
rect 12620 9590 12640 9630
rect 12680 9590 12700 9630
rect 12620 9530 12700 9590
rect 12620 9490 12640 9530
rect 12680 9490 12700 9530
rect 12620 9460 12700 9490
rect 12730 9630 12810 9660
rect 12730 9590 12750 9630
rect 12790 9590 12810 9630
rect 12730 9530 12810 9590
rect 12730 9490 12750 9530
rect 12790 9490 12810 9530
rect 12730 9460 12810 9490
rect 12840 9630 12920 9660
rect 12840 9590 12860 9630
rect 12900 9590 12920 9630
rect 12840 9530 12920 9590
rect 12840 9490 12860 9530
rect 12900 9490 12920 9530
rect 12840 9460 12920 9490
rect 12950 9630 13030 9660
rect 12950 9590 12970 9630
rect 13010 9590 13030 9630
rect 12950 9530 13030 9590
rect 12950 9490 12970 9530
rect 13010 9490 13030 9530
rect 12950 9460 13030 9490
rect 13530 9630 13610 9660
rect 13530 9590 13550 9630
rect 13590 9590 13610 9630
rect 13530 9530 13610 9590
rect 13530 9490 13550 9530
rect 13590 9490 13610 9530
rect 13530 9460 13610 9490
rect 13640 9630 13720 9660
rect 13640 9590 13660 9630
rect 13700 9590 13720 9630
rect 13640 9530 13720 9590
rect 13640 9490 13660 9530
rect 13700 9490 13720 9530
rect 13640 9460 13720 9490
rect 13750 9630 13830 9660
rect 13750 9590 13770 9630
rect 13810 9590 13830 9630
rect 13750 9530 13830 9590
rect 13750 9490 13770 9530
rect 13810 9490 13830 9530
rect 13750 9460 13830 9490
rect 13860 9630 13940 9660
rect 13860 9590 13880 9630
rect 13920 9590 13940 9630
rect 13860 9530 13940 9590
rect 13860 9490 13880 9530
rect 13920 9490 13940 9530
rect 13860 9460 13940 9490
rect 13970 9630 14050 9660
rect 13970 9590 13990 9630
rect 14030 9590 14050 9630
rect 13970 9530 14050 9590
rect 13970 9490 13990 9530
rect 14030 9490 14050 9530
rect 13970 9460 14050 9490
rect 14080 9630 14160 9660
rect 14080 9590 14100 9630
rect 14140 9590 14160 9630
rect 14080 9530 14160 9590
rect 14080 9490 14100 9530
rect 14140 9490 14160 9530
rect 14080 9460 14160 9490
rect 14190 9630 14270 9660
rect 14190 9590 14210 9630
rect 14250 9590 14270 9630
rect 14190 9530 14270 9590
rect 14190 9490 14210 9530
rect 14250 9490 14270 9530
rect 14190 9460 14270 9490
rect 14300 9630 14380 9660
rect 14300 9590 14320 9630
rect 14360 9590 14380 9630
rect 14300 9530 14380 9590
rect 14300 9490 14320 9530
rect 14360 9490 14380 9530
rect 14300 9460 14380 9490
rect 14410 9630 14490 9660
rect 14410 9590 14430 9630
rect 14470 9590 14490 9630
rect 14410 9530 14490 9590
rect 14410 9490 14430 9530
rect 14470 9490 14490 9530
rect 14410 9460 14490 9490
rect 14520 9630 14600 9660
rect 14520 9590 14540 9630
rect 14580 9590 14600 9630
rect 14520 9530 14600 9590
rect 14520 9490 14540 9530
rect 14580 9490 14600 9530
rect 14520 9460 14600 9490
rect 14630 9630 14710 9660
rect 14630 9590 14650 9630
rect 14690 9590 14710 9630
rect 14630 9530 14710 9590
rect 14630 9490 14650 9530
rect 14690 9490 14710 9530
rect 14630 9460 14710 9490
rect 14740 9630 14820 9660
rect 14740 9590 14760 9630
rect 14800 9590 14820 9630
rect 14740 9530 14820 9590
rect 14740 9490 14760 9530
rect 14800 9490 14820 9530
rect 14740 9460 14820 9490
rect 14850 9630 14930 9660
rect 14850 9590 14870 9630
rect 14910 9590 14930 9630
rect 14850 9530 14930 9590
rect 14850 9490 14870 9530
rect 14910 9490 14930 9530
rect 14850 9460 14930 9490
<< ndiffc >>
rect 11180 14210 11220 14250
rect 11180 14110 11220 14150
rect 13260 14210 13300 14250
rect 13260 14110 13300 14150
rect 15340 14210 15380 14250
rect 15340 14110 15380 14150
rect 10760 13600 10800 13640
rect 10760 13500 10800 13540
rect 10760 13400 10800 13440
rect 10760 13300 10800 13340
rect 10760 13200 10800 13240
rect 11840 13600 11880 13640
rect 12000 13600 12040 13640
rect 11840 13500 11880 13540
rect 12000 13500 12040 13540
rect 11840 13400 11880 13440
rect 12000 13400 12040 13440
rect 11840 13300 11880 13340
rect 12000 13300 12040 13340
rect 11840 13200 11880 13240
rect 12000 13200 12040 13240
rect 13080 13600 13120 13640
rect 13080 13500 13120 13540
rect 13080 13400 13120 13440
rect 13080 13300 13120 13340
rect 13080 13200 13120 13240
rect 13440 13600 13480 13640
rect 13440 13500 13480 13540
rect 13440 13400 13480 13440
rect 13440 13300 13480 13340
rect 13440 13200 13480 13240
rect 14520 13600 14560 13640
rect 14680 13600 14720 13640
rect 14520 13500 14560 13540
rect 14680 13500 14720 13540
rect 14520 13400 14560 13440
rect 14680 13400 14720 13440
rect 14520 13300 14560 13340
rect 14680 13300 14720 13340
rect 14520 13200 14560 13240
rect 14680 13200 14720 13240
rect 15760 13600 15800 13640
rect 15760 13500 15800 13540
rect 15760 13400 15800 13440
rect 15760 13300 15800 13340
rect 15760 13200 15800 13240
rect 11380 12590 11420 12630
rect 11500 12590 11540 12630
rect 11620 12590 11660 12630
rect 11740 12590 11780 12630
rect 11860 12590 11900 12630
rect 11980 12590 12020 12630
rect 12100 12590 12140 12630
rect 12220 12590 12260 12630
rect 12340 12590 12380 12630
rect 12460 12590 12500 12630
rect 12580 12590 12620 12630
rect 13940 12590 13980 12630
rect 14060 12590 14100 12630
rect 14180 12590 14220 12630
rect 14300 12590 14340 12630
rect 14420 12590 14460 12630
rect 14540 12590 14580 12630
rect 14660 12590 14700 12630
rect 14780 12590 14820 12630
rect 14900 12590 14940 12630
rect 15020 12590 15060 12630
rect 15140 12590 15180 12630
<< pdiffc >>
rect 11632 18392 11666 18426
rect 11722 18392 11756 18426
rect 11812 18392 11846 18426
rect 11902 18392 11936 18426
rect 11992 18392 12026 18426
rect 12082 18392 12116 18426
rect 12172 18392 12206 18426
rect 11632 18302 11666 18336
rect 11722 18302 11756 18336
rect 11812 18302 11846 18336
rect 11902 18302 11936 18336
rect 11992 18302 12026 18336
rect 12082 18302 12116 18336
rect 12172 18302 12206 18336
rect 11632 18212 11666 18246
rect 11722 18212 11756 18246
rect 11812 18212 11846 18246
rect 11902 18212 11936 18246
rect 11992 18212 12026 18246
rect 12082 18212 12116 18246
rect 12172 18212 12206 18246
rect 11632 18122 11666 18156
rect 11722 18122 11756 18156
rect 11812 18122 11846 18156
rect 11902 18122 11936 18156
rect 11992 18122 12026 18156
rect 12082 18122 12116 18156
rect 12172 18122 12206 18156
rect 11632 18032 11666 18066
rect 11722 18032 11756 18066
rect 11812 18032 11846 18066
rect 11902 18032 11936 18066
rect 11992 18032 12026 18066
rect 12082 18032 12116 18066
rect 12172 18032 12206 18066
rect 11632 17942 11666 17976
rect 11722 17942 11756 17976
rect 11812 17942 11846 17976
rect 11902 17942 11936 17976
rect 11992 17942 12026 17976
rect 12082 17942 12116 17976
rect 12172 17942 12206 17976
rect 11632 17852 11666 17886
rect 11722 17852 11756 17886
rect 11812 17852 11846 17886
rect 11902 17852 11936 17886
rect 11992 17852 12026 17886
rect 12082 17852 12116 17886
rect 12172 17852 12206 17886
rect 12992 18392 13026 18426
rect 13082 18392 13116 18426
rect 13172 18392 13206 18426
rect 13262 18392 13296 18426
rect 13352 18392 13386 18426
rect 13442 18392 13476 18426
rect 13532 18392 13566 18426
rect 12992 18302 13026 18336
rect 13082 18302 13116 18336
rect 13172 18302 13206 18336
rect 13262 18302 13296 18336
rect 13352 18302 13386 18336
rect 13442 18302 13476 18336
rect 13532 18302 13566 18336
rect 12992 18212 13026 18246
rect 13082 18212 13116 18246
rect 13172 18212 13206 18246
rect 13262 18212 13296 18246
rect 13352 18212 13386 18246
rect 13442 18212 13476 18246
rect 13532 18212 13566 18246
rect 12992 18122 13026 18156
rect 13082 18122 13116 18156
rect 13172 18122 13206 18156
rect 13262 18122 13296 18156
rect 13352 18122 13386 18156
rect 13442 18122 13476 18156
rect 13532 18122 13566 18156
rect 12992 18032 13026 18066
rect 13082 18032 13116 18066
rect 13172 18032 13206 18066
rect 13262 18032 13296 18066
rect 13352 18032 13386 18066
rect 13442 18032 13476 18066
rect 13532 18032 13566 18066
rect 12992 17942 13026 17976
rect 13082 17942 13116 17976
rect 13172 17942 13206 17976
rect 13262 17942 13296 17976
rect 13352 17942 13386 17976
rect 13442 17942 13476 17976
rect 13532 17942 13566 17976
rect 12992 17852 13026 17886
rect 13082 17852 13116 17886
rect 13172 17852 13206 17886
rect 13262 17852 13296 17886
rect 13352 17852 13386 17886
rect 13442 17852 13476 17886
rect 13532 17852 13566 17886
rect 14352 18392 14386 18426
rect 14442 18392 14476 18426
rect 14532 18392 14566 18426
rect 14622 18392 14656 18426
rect 14712 18392 14746 18426
rect 14802 18392 14836 18426
rect 14892 18392 14926 18426
rect 14352 18302 14386 18336
rect 14442 18302 14476 18336
rect 14532 18302 14566 18336
rect 14622 18302 14656 18336
rect 14712 18302 14746 18336
rect 14802 18302 14836 18336
rect 14892 18302 14926 18336
rect 14352 18212 14386 18246
rect 14442 18212 14476 18246
rect 14532 18212 14566 18246
rect 14622 18212 14656 18246
rect 14712 18212 14746 18246
rect 14802 18212 14836 18246
rect 14892 18212 14926 18246
rect 14352 18122 14386 18156
rect 14442 18122 14476 18156
rect 14532 18122 14566 18156
rect 14622 18122 14656 18156
rect 14712 18122 14746 18156
rect 14802 18122 14836 18156
rect 14892 18122 14926 18156
rect 14352 18032 14386 18066
rect 14442 18032 14476 18066
rect 14532 18032 14566 18066
rect 14622 18032 14656 18066
rect 14712 18032 14746 18066
rect 14802 18032 14836 18066
rect 14892 18032 14926 18066
rect 14352 17942 14386 17976
rect 14442 17942 14476 17976
rect 14532 17942 14566 17976
rect 14622 17942 14656 17976
rect 14712 17942 14746 17976
rect 14802 17942 14836 17976
rect 14892 17942 14926 17976
rect 14352 17852 14386 17886
rect 14442 17852 14476 17886
rect 14532 17852 14566 17886
rect 14622 17852 14656 17886
rect 14712 17852 14746 17886
rect 14802 17852 14836 17886
rect 14892 17852 14926 17886
rect 11632 17032 11666 17066
rect 11722 17032 11756 17066
rect 11812 17032 11846 17066
rect 11902 17032 11936 17066
rect 11992 17032 12026 17066
rect 12082 17032 12116 17066
rect 12172 17032 12206 17066
rect 11632 16942 11666 16976
rect 11722 16942 11756 16976
rect 11812 16942 11846 16976
rect 11902 16942 11936 16976
rect 11992 16942 12026 16976
rect 12082 16942 12116 16976
rect 12172 16942 12206 16976
rect 11632 16852 11666 16886
rect 11722 16852 11756 16886
rect 11812 16852 11846 16886
rect 11902 16852 11936 16886
rect 11992 16852 12026 16886
rect 12082 16852 12116 16886
rect 12172 16852 12206 16886
rect 11632 16762 11666 16796
rect 11722 16762 11756 16796
rect 11812 16762 11846 16796
rect 11902 16762 11936 16796
rect 11992 16762 12026 16796
rect 12082 16762 12116 16796
rect 12172 16762 12206 16796
rect 11632 16672 11666 16706
rect 11722 16672 11756 16706
rect 11812 16672 11846 16706
rect 11902 16672 11936 16706
rect 11992 16672 12026 16706
rect 12082 16672 12116 16706
rect 12172 16672 12206 16706
rect 11632 16582 11666 16616
rect 11722 16582 11756 16616
rect 11812 16582 11846 16616
rect 11902 16582 11936 16616
rect 11992 16582 12026 16616
rect 12082 16582 12116 16616
rect 12172 16582 12206 16616
rect 11632 16492 11666 16526
rect 11722 16492 11756 16526
rect 11812 16492 11846 16526
rect 11902 16492 11936 16526
rect 11992 16492 12026 16526
rect 12082 16492 12116 16526
rect 12172 16492 12206 16526
rect 12992 17032 13026 17066
rect 13082 17032 13116 17066
rect 13172 17032 13206 17066
rect 13262 17032 13296 17066
rect 13352 17032 13386 17066
rect 13442 17032 13476 17066
rect 13532 17032 13566 17066
rect 12992 16942 13026 16976
rect 13082 16942 13116 16976
rect 13172 16942 13206 16976
rect 13262 16942 13296 16976
rect 13352 16942 13386 16976
rect 13442 16942 13476 16976
rect 13532 16942 13566 16976
rect 12992 16852 13026 16886
rect 13082 16852 13116 16886
rect 13172 16852 13206 16886
rect 13262 16852 13296 16886
rect 13352 16852 13386 16886
rect 13442 16852 13476 16886
rect 13532 16852 13566 16886
rect 12992 16762 13026 16796
rect 13082 16762 13116 16796
rect 13172 16762 13206 16796
rect 13262 16762 13296 16796
rect 13352 16762 13386 16796
rect 13442 16762 13476 16796
rect 13532 16762 13566 16796
rect 12992 16672 13026 16706
rect 13082 16672 13116 16706
rect 13172 16672 13206 16706
rect 13262 16672 13296 16706
rect 13352 16672 13386 16706
rect 13442 16672 13476 16706
rect 13532 16672 13566 16706
rect 12992 16582 13026 16616
rect 13082 16582 13116 16616
rect 13172 16582 13206 16616
rect 13262 16582 13296 16616
rect 13352 16582 13386 16616
rect 13442 16582 13476 16616
rect 13532 16582 13566 16616
rect 12992 16492 13026 16526
rect 13082 16492 13116 16526
rect 13172 16492 13206 16526
rect 13262 16492 13296 16526
rect 13352 16492 13386 16526
rect 13442 16492 13476 16526
rect 13532 16492 13566 16526
rect 14352 17032 14386 17066
rect 14442 17032 14476 17066
rect 14532 17032 14566 17066
rect 14622 17032 14656 17066
rect 14712 17032 14746 17066
rect 14802 17032 14836 17066
rect 14892 17032 14926 17066
rect 14352 16942 14386 16976
rect 14442 16942 14476 16976
rect 14532 16942 14566 16976
rect 14622 16942 14656 16976
rect 14712 16942 14746 16976
rect 14802 16942 14836 16976
rect 14892 16942 14926 16976
rect 14352 16852 14386 16886
rect 14442 16852 14476 16886
rect 14532 16852 14566 16886
rect 14622 16852 14656 16886
rect 14712 16852 14746 16886
rect 14802 16852 14836 16886
rect 14892 16852 14926 16886
rect 14352 16762 14386 16796
rect 14442 16762 14476 16796
rect 14532 16762 14566 16796
rect 14622 16762 14656 16796
rect 14712 16762 14746 16796
rect 14802 16762 14836 16796
rect 14892 16762 14926 16796
rect 14352 16672 14386 16706
rect 14442 16672 14476 16706
rect 14532 16672 14566 16706
rect 14622 16672 14656 16706
rect 14712 16672 14746 16706
rect 14802 16672 14836 16706
rect 14892 16672 14926 16706
rect 14352 16582 14386 16616
rect 14442 16582 14476 16616
rect 14532 16582 14566 16616
rect 14622 16582 14656 16616
rect 14712 16582 14746 16616
rect 14802 16582 14836 16616
rect 14892 16582 14926 16616
rect 14352 16492 14386 16526
rect 14442 16492 14476 16526
rect 14532 16492 14566 16526
rect 14622 16492 14656 16526
rect 14712 16492 14746 16526
rect 14802 16492 14836 16526
rect 14892 16492 14926 16526
rect 11632 15672 11666 15706
rect 11722 15672 11756 15706
rect 11812 15672 11846 15706
rect 11902 15672 11936 15706
rect 11992 15672 12026 15706
rect 12082 15672 12116 15706
rect 12172 15672 12206 15706
rect 11632 15582 11666 15616
rect 11722 15582 11756 15616
rect 11812 15582 11846 15616
rect 11902 15582 11936 15616
rect 11992 15582 12026 15616
rect 12082 15582 12116 15616
rect 12172 15582 12206 15616
rect 11632 15492 11666 15526
rect 11722 15492 11756 15526
rect 11812 15492 11846 15526
rect 11902 15492 11936 15526
rect 11992 15492 12026 15526
rect 12082 15492 12116 15526
rect 12172 15492 12206 15526
rect 11632 15402 11666 15436
rect 11722 15402 11756 15436
rect 11812 15402 11846 15436
rect 11902 15402 11936 15436
rect 11992 15402 12026 15436
rect 12082 15402 12116 15436
rect 12172 15402 12206 15436
rect 11632 15312 11666 15346
rect 11722 15312 11756 15346
rect 11812 15312 11846 15346
rect 11902 15312 11936 15346
rect 11992 15312 12026 15346
rect 12082 15312 12116 15346
rect 12172 15312 12206 15346
rect 11632 15222 11666 15256
rect 11722 15222 11756 15256
rect 11812 15222 11846 15256
rect 11902 15222 11936 15256
rect 11992 15222 12026 15256
rect 12082 15222 12116 15256
rect 12172 15222 12206 15256
rect 11632 15132 11666 15166
rect 11722 15132 11756 15166
rect 11812 15132 11846 15166
rect 11902 15132 11936 15166
rect 11992 15132 12026 15166
rect 12082 15132 12116 15166
rect 12172 15132 12206 15166
rect 12992 15672 13026 15706
rect 13082 15672 13116 15706
rect 13172 15672 13206 15706
rect 13262 15672 13296 15706
rect 13352 15672 13386 15706
rect 13442 15672 13476 15706
rect 13532 15672 13566 15706
rect 12992 15582 13026 15616
rect 13082 15582 13116 15616
rect 13172 15582 13206 15616
rect 13262 15582 13296 15616
rect 13352 15582 13386 15616
rect 13442 15582 13476 15616
rect 13532 15582 13566 15616
rect 12992 15492 13026 15526
rect 13082 15492 13116 15526
rect 13172 15492 13206 15526
rect 13262 15492 13296 15526
rect 13352 15492 13386 15526
rect 13442 15492 13476 15526
rect 13532 15492 13566 15526
rect 12992 15402 13026 15436
rect 13082 15402 13116 15436
rect 13172 15402 13206 15436
rect 13262 15402 13296 15436
rect 13352 15402 13386 15436
rect 13442 15402 13476 15436
rect 13532 15402 13566 15436
rect 12992 15312 13026 15346
rect 13082 15312 13116 15346
rect 13172 15312 13206 15346
rect 13262 15312 13296 15346
rect 13352 15312 13386 15346
rect 13442 15312 13476 15346
rect 13532 15312 13566 15346
rect 12992 15222 13026 15256
rect 13082 15222 13116 15256
rect 13172 15222 13206 15256
rect 13262 15222 13296 15256
rect 13352 15222 13386 15256
rect 13442 15222 13476 15256
rect 13532 15222 13566 15256
rect 12992 15132 13026 15166
rect 13082 15132 13116 15166
rect 13172 15132 13206 15166
rect 13262 15132 13296 15166
rect 13352 15132 13386 15166
rect 13442 15132 13476 15166
rect 13532 15132 13566 15166
rect 14352 15672 14386 15706
rect 14442 15672 14476 15706
rect 14532 15672 14566 15706
rect 14622 15672 14656 15706
rect 14712 15672 14746 15706
rect 14802 15672 14836 15706
rect 14892 15672 14926 15706
rect 14352 15582 14386 15616
rect 14442 15582 14476 15616
rect 14532 15582 14566 15616
rect 14622 15582 14656 15616
rect 14712 15582 14746 15616
rect 14802 15582 14836 15616
rect 14892 15582 14926 15616
rect 14352 15492 14386 15526
rect 14442 15492 14476 15526
rect 14532 15492 14566 15526
rect 14622 15492 14656 15526
rect 14712 15492 14746 15526
rect 14802 15492 14836 15526
rect 14892 15492 14926 15526
rect 14352 15402 14386 15436
rect 14442 15402 14476 15436
rect 14532 15402 14566 15436
rect 14622 15402 14656 15436
rect 14712 15402 14746 15436
rect 14802 15402 14836 15436
rect 14892 15402 14926 15436
rect 14352 15312 14386 15346
rect 14442 15312 14476 15346
rect 14532 15312 14566 15346
rect 14622 15312 14656 15346
rect 14712 15312 14746 15346
rect 14802 15312 14836 15346
rect 14892 15312 14926 15346
rect 14352 15222 14386 15256
rect 14442 15222 14476 15256
rect 14532 15222 14566 15256
rect 14622 15222 14656 15256
rect 14712 15222 14746 15256
rect 14802 15222 14836 15256
rect 14892 15222 14926 15256
rect 14352 15132 14386 15166
rect 14442 15132 14476 15166
rect 14532 15132 14566 15166
rect 14622 15132 14656 15166
rect 14712 15132 14746 15166
rect 14802 15132 14836 15166
rect 14892 15132 14926 15166
rect 10540 11750 10580 11790
rect 10540 11650 10580 11690
rect 10660 11750 10700 11790
rect 10660 11650 10700 11690
rect 10780 11750 10820 11790
rect 10780 11650 10820 11690
rect 10900 11750 10940 11790
rect 10900 11650 10940 11690
rect 11020 11750 11060 11790
rect 11020 11650 11060 11690
rect 11140 11750 11180 11790
rect 11140 11650 11180 11690
rect 11260 11750 11300 11790
rect 11260 11650 11300 11690
rect 11380 11750 11420 11790
rect 11380 11650 11420 11690
rect 11500 11750 11540 11790
rect 11500 11650 11540 11690
rect 11620 11750 11660 11790
rect 11620 11650 11660 11690
rect 11740 11750 11780 11790
rect 11740 11650 11780 11690
rect 11860 11750 11900 11790
rect 11860 11650 11900 11690
rect 11980 11750 12020 11790
rect 11980 11650 12020 11690
rect 12100 11750 12140 11790
rect 12100 11650 12140 11690
rect 12220 11750 12260 11790
rect 12220 11650 12260 11690
rect 12340 11750 12380 11790
rect 12340 11650 12380 11690
rect 12460 11750 12500 11790
rect 12460 11650 12500 11690
rect 12580 11750 12620 11790
rect 12580 11650 12620 11690
rect 12700 11750 12740 11790
rect 12700 11650 12740 11690
rect 12820 11750 12860 11790
rect 12820 11650 12860 11690
rect 12940 11750 12980 11790
rect 12940 11650 12980 11690
rect 13580 11750 13620 11790
rect 13580 11650 13620 11690
rect 13700 11750 13740 11790
rect 13700 11650 13740 11690
rect 13820 11750 13860 11790
rect 13820 11650 13860 11690
rect 13940 11750 13980 11790
rect 13940 11650 13980 11690
rect 14060 11750 14100 11790
rect 14060 11650 14100 11690
rect 14180 11750 14220 11790
rect 14180 11650 14220 11690
rect 14300 11750 14340 11790
rect 14300 11650 14340 11690
rect 14420 11750 14460 11790
rect 14420 11650 14460 11690
rect 14540 11750 14580 11790
rect 14540 11650 14580 11690
rect 14660 11750 14700 11790
rect 14660 11650 14700 11690
rect 14780 11750 14820 11790
rect 14780 11650 14820 11690
rect 14900 11750 14940 11790
rect 14900 11650 14940 11690
rect 15020 11750 15060 11790
rect 15020 11650 15060 11690
rect 15140 11750 15180 11790
rect 15140 11650 15180 11690
rect 15260 11750 15300 11790
rect 15260 11650 15300 11690
rect 15380 11750 15420 11790
rect 15380 11650 15420 11690
rect 15500 11750 15540 11790
rect 15500 11650 15540 11690
rect 15620 11750 15660 11790
rect 15620 11650 15660 11690
rect 15740 11750 15780 11790
rect 15740 11650 15780 11690
rect 15860 11750 15900 11790
rect 15860 11650 15900 11690
rect 15980 11750 16020 11790
rect 15980 11650 16020 11690
rect 11640 10590 11680 10630
rect 11640 10490 11680 10530
rect 11640 10390 11680 10430
rect 11640 10290 11680 10330
rect 11640 10190 11680 10230
rect 11640 10090 11680 10130
rect 11820 10590 11860 10630
rect 11820 10490 11860 10530
rect 11820 10390 11860 10430
rect 11820 10290 11860 10330
rect 11820 10190 11860 10230
rect 11820 10090 11860 10130
rect 12000 10590 12040 10630
rect 12000 10490 12040 10530
rect 12000 10390 12040 10430
rect 12000 10290 12040 10330
rect 12000 10190 12040 10230
rect 12000 10090 12040 10130
rect 12180 10590 12220 10630
rect 12180 10490 12220 10530
rect 12180 10390 12220 10430
rect 12180 10290 12220 10330
rect 12180 10190 12220 10230
rect 12180 10090 12220 10130
rect 12360 10590 12400 10630
rect 12360 10490 12400 10530
rect 12360 10390 12400 10430
rect 12360 10290 12400 10330
rect 12360 10190 12400 10230
rect 12360 10090 12400 10130
rect 12540 10590 12580 10630
rect 12540 10490 12580 10530
rect 12540 10390 12580 10430
rect 12540 10290 12580 10330
rect 12540 10190 12580 10230
rect 12540 10090 12580 10130
rect 12720 10590 12760 10630
rect 12720 10490 12760 10530
rect 12720 10390 12760 10430
rect 12720 10290 12760 10330
rect 12720 10190 12760 10230
rect 12720 10090 12760 10130
rect 12900 10590 12940 10630
rect 12900 10490 12940 10530
rect 12900 10390 12940 10430
rect 12900 10290 12940 10330
rect 12900 10190 12940 10230
rect 12900 10090 12940 10130
rect 13080 10590 13120 10630
rect 13080 10490 13120 10530
rect 13080 10390 13120 10430
rect 13080 10290 13120 10330
rect 13080 10190 13120 10230
rect 13080 10090 13120 10130
rect 13260 10590 13300 10630
rect 13260 10490 13300 10530
rect 13260 10390 13300 10430
rect 13260 10290 13300 10330
rect 13260 10190 13300 10230
rect 13260 10090 13300 10130
rect 13440 10590 13480 10630
rect 13440 10490 13480 10530
rect 13440 10390 13480 10430
rect 13440 10290 13480 10330
rect 13440 10190 13480 10230
rect 13440 10090 13480 10130
rect 13620 10590 13660 10630
rect 13620 10490 13660 10530
rect 13620 10390 13660 10430
rect 13620 10290 13660 10330
rect 13620 10190 13660 10230
rect 13620 10090 13660 10130
rect 13800 10590 13840 10630
rect 13800 10490 13840 10530
rect 13800 10390 13840 10430
rect 13800 10290 13840 10330
rect 13800 10190 13840 10230
rect 13800 10090 13840 10130
rect 13980 10590 14020 10630
rect 13980 10490 14020 10530
rect 13980 10390 14020 10430
rect 13980 10290 14020 10330
rect 13980 10190 14020 10230
rect 13980 10090 14020 10130
rect 14160 10590 14200 10630
rect 14160 10490 14200 10530
rect 14160 10390 14200 10430
rect 14160 10290 14200 10330
rect 14160 10190 14200 10230
rect 14160 10090 14200 10130
rect 14340 10590 14380 10630
rect 14340 10490 14380 10530
rect 14340 10390 14380 10430
rect 14340 10290 14380 10330
rect 14340 10190 14380 10230
rect 14340 10090 14380 10130
rect 14520 10590 14560 10630
rect 14520 10490 14560 10530
rect 14520 10390 14560 10430
rect 14520 10290 14560 10330
rect 14520 10190 14560 10230
rect 14520 10090 14560 10130
rect 14700 10590 14740 10630
rect 14700 10490 14740 10530
rect 14700 10390 14740 10430
rect 14700 10290 14740 10330
rect 14700 10190 14740 10230
rect 14700 10090 14740 10130
rect 14880 10590 14920 10630
rect 14880 10490 14920 10530
rect 14880 10390 14920 10430
rect 14880 10290 14920 10330
rect 15510 10390 15550 10430
rect 15510 10290 15550 10330
rect 15620 10390 15660 10430
rect 15620 10290 15660 10330
rect 15730 10390 15770 10430
rect 15730 10290 15770 10330
rect 15840 10390 15880 10430
rect 15840 10290 15880 10330
rect 15950 10390 15990 10430
rect 15950 10290 15990 10330
rect 14880 10190 14920 10230
rect 14880 10090 14920 10130
rect 11650 9590 11690 9630
rect 11650 9490 11690 9530
rect 11760 9590 11800 9630
rect 11760 9490 11800 9530
rect 11870 9590 11910 9630
rect 11870 9490 11910 9530
rect 11980 9590 12020 9630
rect 11980 9490 12020 9530
rect 12090 9590 12130 9630
rect 12090 9490 12130 9530
rect 12200 9590 12240 9630
rect 12200 9490 12240 9530
rect 12310 9590 12350 9630
rect 12310 9490 12350 9530
rect 12420 9590 12460 9630
rect 12420 9490 12460 9530
rect 12530 9590 12570 9630
rect 12530 9490 12570 9530
rect 12640 9590 12680 9630
rect 12640 9490 12680 9530
rect 12750 9590 12790 9630
rect 12750 9490 12790 9530
rect 12860 9590 12900 9630
rect 12860 9490 12900 9530
rect 12970 9590 13010 9630
rect 12970 9490 13010 9530
rect 13550 9590 13590 9630
rect 13550 9490 13590 9530
rect 13660 9590 13700 9630
rect 13660 9490 13700 9530
rect 13770 9590 13810 9630
rect 13770 9490 13810 9530
rect 13880 9590 13920 9630
rect 13880 9490 13920 9530
rect 13990 9590 14030 9630
rect 13990 9490 14030 9530
rect 14100 9590 14140 9630
rect 14100 9490 14140 9530
rect 14210 9590 14250 9630
rect 14210 9490 14250 9530
rect 14320 9590 14360 9630
rect 14320 9490 14360 9530
rect 14430 9590 14470 9630
rect 14430 9490 14470 9530
rect 14540 9590 14580 9630
rect 14540 9490 14580 9530
rect 14650 9590 14690 9630
rect 14650 9490 14690 9530
rect 14760 9590 14800 9630
rect 14760 9490 14800 9530
rect 14870 9590 14910 9630
rect 14870 9490 14910 9530
<< psubdiff >>
rect 13230 19070 13330 19100
rect 13230 19030 13260 19070
rect 13300 19030 13330 19070
rect 13230 18990 13330 19030
rect 13230 18950 13260 18990
rect 13300 18950 13330 18990
rect 13230 18910 13330 18950
rect 13230 18870 13260 18910
rect 13300 18870 13330 18910
rect 13230 18840 13330 18870
rect 11276 18752 12564 18784
rect 11276 18718 11410 18752
rect 11444 18718 11500 18752
rect 11534 18718 11590 18752
rect 11624 18718 11680 18752
rect 11714 18718 11770 18752
rect 11804 18718 11860 18752
rect 11894 18718 11950 18752
rect 11984 18718 12040 18752
rect 12074 18718 12130 18752
rect 12164 18718 12220 18752
rect 12254 18718 12310 18752
rect 12344 18718 12400 18752
rect 12434 18718 12564 18752
rect 11276 18683 12564 18718
rect 11276 18668 11377 18683
rect 11276 18634 11309 18668
rect 11343 18634 11377 18668
rect 11276 18578 11377 18634
rect 12463 18668 12564 18683
rect 12463 18634 12496 18668
rect 12530 18634 12564 18668
rect 11276 18544 11309 18578
rect 11343 18544 11377 18578
rect 11276 18488 11377 18544
rect 11276 18454 11309 18488
rect 11343 18454 11377 18488
rect 11276 18398 11377 18454
rect 11276 18364 11309 18398
rect 11343 18364 11377 18398
rect 11276 18308 11377 18364
rect 11276 18274 11309 18308
rect 11343 18274 11377 18308
rect 11276 18218 11377 18274
rect 11276 18184 11309 18218
rect 11343 18184 11377 18218
rect 11276 18128 11377 18184
rect 11276 18094 11309 18128
rect 11343 18094 11377 18128
rect 11276 18038 11377 18094
rect 11276 18004 11309 18038
rect 11343 18004 11377 18038
rect 11276 17948 11377 18004
rect 11276 17914 11309 17948
rect 11343 17914 11377 17948
rect 11276 17858 11377 17914
rect 11276 17824 11309 17858
rect 11343 17824 11377 17858
rect 11276 17768 11377 17824
rect 11276 17734 11309 17768
rect 11343 17734 11377 17768
rect 11276 17678 11377 17734
rect 11276 17644 11309 17678
rect 11343 17644 11377 17678
rect 12463 18578 12564 18634
rect 12463 18544 12496 18578
rect 12530 18544 12564 18578
rect 12463 18488 12564 18544
rect 12463 18454 12496 18488
rect 12530 18454 12564 18488
rect 12463 18398 12564 18454
rect 12463 18364 12496 18398
rect 12530 18364 12564 18398
rect 12463 18308 12564 18364
rect 12463 18274 12496 18308
rect 12530 18274 12564 18308
rect 12463 18218 12564 18274
rect 12463 18184 12496 18218
rect 12530 18184 12564 18218
rect 12463 18128 12564 18184
rect 12463 18094 12496 18128
rect 12530 18094 12564 18128
rect 12463 18038 12564 18094
rect 12463 18004 12496 18038
rect 12530 18004 12564 18038
rect 12463 17948 12564 18004
rect 12463 17914 12496 17948
rect 12530 17914 12564 17948
rect 12463 17858 12564 17914
rect 12463 17824 12496 17858
rect 12530 17824 12564 17858
rect 12463 17768 12564 17824
rect 12463 17734 12496 17768
rect 12530 17734 12564 17768
rect 12463 17678 12564 17734
rect 11276 17597 11377 17644
rect 12463 17644 12496 17678
rect 12530 17644 12564 17678
rect 12463 17597 12564 17644
rect 11276 17588 12564 17597
rect 11276 17554 11309 17588
rect 11343 17565 12496 17588
rect 11343 17554 11410 17565
rect 11276 17531 11410 17554
rect 11444 17531 11500 17565
rect 11534 17531 11590 17565
rect 11624 17531 11680 17565
rect 11714 17531 11770 17565
rect 11804 17531 11860 17565
rect 11894 17531 11950 17565
rect 11984 17531 12040 17565
rect 12074 17531 12130 17565
rect 12164 17531 12220 17565
rect 12254 17531 12310 17565
rect 12344 17531 12400 17565
rect 12434 17554 12496 17565
rect 12530 17554 12564 17588
rect 12434 17531 12564 17554
rect 11276 17496 12564 17531
rect 12636 18752 13924 18784
rect 12636 18718 12770 18752
rect 12804 18718 12860 18752
rect 12894 18718 12950 18752
rect 12984 18718 13040 18752
rect 13074 18718 13130 18752
rect 13164 18718 13220 18752
rect 13254 18718 13310 18752
rect 13344 18718 13400 18752
rect 13434 18718 13490 18752
rect 13524 18718 13580 18752
rect 13614 18718 13670 18752
rect 13704 18718 13760 18752
rect 13794 18718 13924 18752
rect 12636 18683 13924 18718
rect 12636 18668 12737 18683
rect 12636 18634 12669 18668
rect 12703 18634 12737 18668
rect 12636 18578 12737 18634
rect 13823 18668 13924 18683
rect 13823 18634 13856 18668
rect 13890 18634 13924 18668
rect 12636 18544 12669 18578
rect 12703 18544 12737 18578
rect 12636 18488 12737 18544
rect 12636 18454 12669 18488
rect 12703 18454 12737 18488
rect 12636 18398 12737 18454
rect 12636 18364 12669 18398
rect 12703 18364 12737 18398
rect 12636 18308 12737 18364
rect 12636 18274 12669 18308
rect 12703 18274 12737 18308
rect 12636 18218 12737 18274
rect 12636 18184 12669 18218
rect 12703 18184 12737 18218
rect 12636 18128 12737 18184
rect 12636 18094 12669 18128
rect 12703 18094 12737 18128
rect 12636 18038 12737 18094
rect 12636 18004 12669 18038
rect 12703 18004 12737 18038
rect 12636 17948 12737 18004
rect 12636 17914 12669 17948
rect 12703 17914 12737 17948
rect 12636 17858 12737 17914
rect 12636 17824 12669 17858
rect 12703 17824 12737 17858
rect 12636 17768 12737 17824
rect 12636 17734 12669 17768
rect 12703 17734 12737 17768
rect 12636 17678 12737 17734
rect 12636 17644 12669 17678
rect 12703 17644 12737 17678
rect 13823 18578 13924 18634
rect 13823 18544 13856 18578
rect 13890 18544 13924 18578
rect 13823 18488 13924 18544
rect 13823 18454 13856 18488
rect 13890 18454 13924 18488
rect 13823 18398 13924 18454
rect 13823 18364 13856 18398
rect 13890 18364 13924 18398
rect 13823 18308 13924 18364
rect 13823 18274 13856 18308
rect 13890 18274 13924 18308
rect 13823 18218 13924 18274
rect 13823 18184 13856 18218
rect 13890 18184 13924 18218
rect 13823 18128 13924 18184
rect 13823 18094 13856 18128
rect 13890 18094 13924 18128
rect 13823 18038 13924 18094
rect 13823 18004 13856 18038
rect 13890 18004 13924 18038
rect 13823 17948 13924 18004
rect 13823 17914 13856 17948
rect 13890 17914 13924 17948
rect 13823 17858 13924 17914
rect 13823 17824 13856 17858
rect 13890 17824 13924 17858
rect 13823 17768 13924 17824
rect 13823 17734 13856 17768
rect 13890 17734 13924 17768
rect 13823 17678 13924 17734
rect 12636 17597 12737 17644
rect 13823 17644 13856 17678
rect 13890 17644 13924 17678
rect 13823 17597 13924 17644
rect 12636 17588 13924 17597
rect 12636 17554 12669 17588
rect 12703 17565 13856 17588
rect 12703 17554 12770 17565
rect 12636 17531 12770 17554
rect 12804 17531 12860 17565
rect 12894 17531 12950 17565
rect 12984 17531 13040 17565
rect 13074 17531 13130 17565
rect 13164 17531 13220 17565
rect 13254 17531 13310 17565
rect 13344 17531 13400 17565
rect 13434 17531 13490 17565
rect 13524 17531 13580 17565
rect 13614 17531 13670 17565
rect 13704 17531 13760 17565
rect 13794 17554 13856 17565
rect 13890 17554 13924 17588
rect 13794 17531 13924 17554
rect 12636 17496 13924 17531
rect 13996 18752 15284 18784
rect 13996 18718 14130 18752
rect 14164 18718 14220 18752
rect 14254 18718 14310 18752
rect 14344 18718 14400 18752
rect 14434 18718 14490 18752
rect 14524 18718 14580 18752
rect 14614 18718 14670 18752
rect 14704 18718 14760 18752
rect 14794 18718 14850 18752
rect 14884 18718 14940 18752
rect 14974 18718 15030 18752
rect 15064 18718 15120 18752
rect 15154 18718 15284 18752
rect 13996 18683 15284 18718
rect 13996 18668 14097 18683
rect 13996 18634 14029 18668
rect 14063 18634 14097 18668
rect 13996 18578 14097 18634
rect 15183 18668 15284 18683
rect 15183 18634 15216 18668
rect 15250 18634 15284 18668
rect 13996 18544 14029 18578
rect 14063 18544 14097 18578
rect 13996 18488 14097 18544
rect 13996 18454 14029 18488
rect 14063 18454 14097 18488
rect 13996 18398 14097 18454
rect 13996 18364 14029 18398
rect 14063 18364 14097 18398
rect 13996 18308 14097 18364
rect 13996 18274 14029 18308
rect 14063 18274 14097 18308
rect 13996 18218 14097 18274
rect 13996 18184 14029 18218
rect 14063 18184 14097 18218
rect 13996 18128 14097 18184
rect 13996 18094 14029 18128
rect 14063 18094 14097 18128
rect 13996 18038 14097 18094
rect 13996 18004 14029 18038
rect 14063 18004 14097 18038
rect 13996 17948 14097 18004
rect 13996 17914 14029 17948
rect 14063 17914 14097 17948
rect 13996 17858 14097 17914
rect 13996 17824 14029 17858
rect 14063 17824 14097 17858
rect 13996 17768 14097 17824
rect 13996 17734 14029 17768
rect 14063 17734 14097 17768
rect 13996 17678 14097 17734
rect 13996 17644 14029 17678
rect 14063 17644 14097 17678
rect 15183 18578 15284 18634
rect 15183 18544 15216 18578
rect 15250 18544 15284 18578
rect 15183 18488 15284 18544
rect 15183 18454 15216 18488
rect 15250 18454 15284 18488
rect 15183 18398 15284 18454
rect 15183 18364 15216 18398
rect 15250 18364 15284 18398
rect 15183 18308 15284 18364
rect 15183 18274 15216 18308
rect 15250 18274 15284 18308
rect 15183 18218 15284 18274
rect 15183 18184 15216 18218
rect 15250 18184 15284 18218
rect 15183 18128 15284 18184
rect 15183 18094 15216 18128
rect 15250 18094 15284 18128
rect 15183 18038 15284 18094
rect 15183 18004 15216 18038
rect 15250 18004 15284 18038
rect 15183 17948 15284 18004
rect 15183 17914 15216 17948
rect 15250 17914 15284 17948
rect 15183 17858 15284 17914
rect 15183 17824 15216 17858
rect 15250 17824 15284 17858
rect 15183 17768 15284 17824
rect 15183 17734 15216 17768
rect 15250 17734 15284 17768
rect 15183 17678 15284 17734
rect 13996 17597 14097 17644
rect 15183 17644 15216 17678
rect 15250 17644 15284 17678
rect 15183 17597 15284 17644
rect 13996 17588 15284 17597
rect 13996 17554 14029 17588
rect 14063 17565 15216 17588
rect 14063 17554 14130 17565
rect 13996 17531 14130 17554
rect 14164 17531 14220 17565
rect 14254 17531 14310 17565
rect 14344 17531 14400 17565
rect 14434 17531 14490 17565
rect 14524 17531 14580 17565
rect 14614 17531 14670 17565
rect 14704 17531 14760 17565
rect 14794 17531 14850 17565
rect 14884 17531 14940 17565
rect 14974 17531 15030 17565
rect 15064 17531 15120 17565
rect 15154 17554 15216 17565
rect 15250 17554 15284 17588
rect 15154 17531 15284 17554
rect 13996 17496 15284 17531
rect 11276 17392 12564 17424
rect 11276 17358 11410 17392
rect 11444 17358 11500 17392
rect 11534 17358 11590 17392
rect 11624 17358 11680 17392
rect 11714 17358 11770 17392
rect 11804 17358 11860 17392
rect 11894 17358 11950 17392
rect 11984 17358 12040 17392
rect 12074 17358 12130 17392
rect 12164 17358 12220 17392
rect 12254 17358 12310 17392
rect 12344 17358 12400 17392
rect 12434 17358 12564 17392
rect 11276 17323 12564 17358
rect 11276 17308 11377 17323
rect 11276 17274 11309 17308
rect 11343 17274 11377 17308
rect 11276 17218 11377 17274
rect 12463 17308 12564 17323
rect 12463 17274 12496 17308
rect 12530 17274 12564 17308
rect 11276 17184 11309 17218
rect 11343 17184 11377 17218
rect 11276 17128 11377 17184
rect 11276 17094 11309 17128
rect 11343 17094 11377 17128
rect 11276 17038 11377 17094
rect 11276 17004 11309 17038
rect 11343 17004 11377 17038
rect 11276 16948 11377 17004
rect 11276 16914 11309 16948
rect 11343 16914 11377 16948
rect 11276 16858 11377 16914
rect 11276 16824 11309 16858
rect 11343 16824 11377 16858
rect 11276 16768 11377 16824
rect 11276 16734 11309 16768
rect 11343 16734 11377 16768
rect 11276 16678 11377 16734
rect 11276 16644 11309 16678
rect 11343 16644 11377 16678
rect 11276 16588 11377 16644
rect 11276 16554 11309 16588
rect 11343 16554 11377 16588
rect 11276 16498 11377 16554
rect 11276 16464 11309 16498
rect 11343 16464 11377 16498
rect 11276 16408 11377 16464
rect 11276 16374 11309 16408
rect 11343 16374 11377 16408
rect 11276 16318 11377 16374
rect 11276 16284 11309 16318
rect 11343 16284 11377 16318
rect 12463 17218 12564 17274
rect 12463 17184 12496 17218
rect 12530 17184 12564 17218
rect 12463 17128 12564 17184
rect 12463 17094 12496 17128
rect 12530 17094 12564 17128
rect 12463 17038 12564 17094
rect 12463 17004 12496 17038
rect 12530 17004 12564 17038
rect 12463 16948 12564 17004
rect 12463 16914 12496 16948
rect 12530 16914 12564 16948
rect 12463 16858 12564 16914
rect 12463 16824 12496 16858
rect 12530 16824 12564 16858
rect 12463 16768 12564 16824
rect 12463 16734 12496 16768
rect 12530 16734 12564 16768
rect 12463 16678 12564 16734
rect 12463 16644 12496 16678
rect 12530 16644 12564 16678
rect 12463 16588 12564 16644
rect 12463 16554 12496 16588
rect 12530 16554 12564 16588
rect 12463 16498 12564 16554
rect 12463 16464 12496 16498
rect 12530 16464 12564 16498
rect 12463 16408 12564 16464
rect 12463 16374 12496 16408
rect 12530 16374 12564 16408
rect 12463 16318 12564 16374
rect 11276 16237 11377 16284
rect 12463 16284 12496 16318
rect 12530 16284 12564 16318
rect 12463 16237 12564 16284
rect 11276 16228 12564 16237
rect 11276 16194 11309 16228
rect 11343 16205 12496 16228
rect 11343 16194 11410 16205
rect 11276 16171 11410 16194
rect 11444 16171 11500 16205
rect 11534 16171 11590 16205
rect 11624 16171 11680 16205
rect 11714 16171 11770 16205
rect 11804 16171 11860 16205
rect 11894 16171 11950 16205
rect 11984 16171 12040 16205
rect 12074 16171 12130 16205
rect 12164 16171 12220 16205
rect 12254 16171 12310 16205
rect 12344 16171 12400 16205
rect 12434 16194 12496 16205
rect 12530 16194 12564 16228
rect 12434 16171 12564 16194
rect 11276 16136 12564 16171
rect 12636 17392 13924 17424
rect 12636 17358 12770 17392
rect 12804 17358 12860 17392
rect 12894 17358 12950 17392
rect 12984 17358 13040 17392
rect 13074 17358 13130 17392
rect 13164 17358 13220 17392
rect 13254 17358 13310 17392
rect 13344 17358 13400 17392
rect 13434 17358 13490 17392
rect 13524 17358 13580 17392
rect 13614 17358 13670 17392
rect 13704 17358 13760 17392
rect 13794 17358 13924 17392
rect 12636 17323 13924 17358
rect 12636 17308 12737 17323
rect 12636 17274 12669 17308
rect 12703 17274 12737 17308
rect 12636 17218 12737 17274
rect 13823 17308 13924 17323
rect 13823 17274 13856 17308
rect 13890 17274 13924 17308
rect 12636 17184 12669 17218
rect 12703 17184 12737 17218
rect 12636 17128 12737 17184
rect 12636 17094 12669 17128
rect 12703 17094 12737 17128
rect 12636 17038 12737 17094
rect 12636 17004 12669 17038
rect 12703 17004 12737 17038
rect 12636 16948 12737 17004
rect 12636 16914 12669 16948
rect 12703 16914 12737 16948
rect 12636 16858 12737 16914
rect 12636 16824 12669 16858
rect 12703 16824 12737 16858
rect 12636 16768 12737 16824
rect 12636 16734 12669 16768
rect 12703 16734 12737 16768
rect 12636 16678 12737 16734
rect 12636 16644 12669 16678
rect 12703 16644 12737 16678
rect 12636 16588 12737 16644
rect 12636 16554 12669 16588
rect 12703 16554 12737 16588
rect 12636 16498 12737 16554
rect 12636 16464 12669 16498
rect 12703 16464 12737 16498
rect 12636 16408 12737 16464
rect 12636 16374 12669 16408
rect 12703 16374 12737 16408
rect 12636 16318 12737 16374
rect 12636 16284 12669 16318
rect 12703 16284 12737 16318
rect 13823 17218 13924 17274
rect 13823 17184 13856 17218
rect 13890 17184 13924 17218
rect 13823 17128 13924 17184
rect 13823 17094 13856 17128
rect 13890 17094 13924 17128
rect 13823 17038 13924 17094
rect 13823 17004 13856 17038
rect 13890 17004 13924 17038
rect 13823 16948 13924 17004
rect 13823 16914 13856 16948
rect 13890 16914 13924 16948
rect 13823 16858 13924 16914
rect 13823 16824 13856 16858
rect 13890 16824 13924 16858
rect 13823 16768 13924 16824
rect 13823 16734 13856 16768
rect 13890 16734 13924 16768
rect 13823 16678 13924 16734
rect 13823 16644 13856 16678
rect 13890 16644 13924 16678
rect 13823 16588 13924 16644
rect 13823 16554 13856 16588
rect 13890 16554 13924 16588
rect 13823 16498 13924 16554
rect 13823 16464 13856 16498
rect 13890 16464 13924 16498
rect 13823 16408 13924 16464
rect 13823 16374 13856 16408
rect 13890 16374 13924 16408
rect 13823 16318 13924 16374
rect 12636 16237 12737 16284
rect 13823 16284 13856 16318
rect 13890 16284 13924 16318
rect 13823 16237 13924 16284
rect 12636 16228 13924 16237
rect 12636 16194 12669 16228
rect 12703 16205 13856 16228
rect 12703 16194 12770 16205
rect 12636 16171 12770 16194
rect 12804 16171 12860 16205
rect 12894 16171 12950 16205
rect 12984 16171 13040 16205
rect 13074 16171 13130 16205
rect 13164 16171 13220 16205
rect 13254 16171 13310 16205
rect 13344 16171 13400 16205
rect 13434 16171 13490 16205
rect 13524 16171 13580 16205
rect 13614 16171 13670 16205
rect 13704 16171 13760 16205
rect 13794 16194 13856 16205
rect 13890 16194 13924 16228
rect 13794 16171 13924 16194
rect 12636 16136 13924 16171
rect 13996 17392 15284 17424
rect 13996 17358 14130 17392
rect 14164 17358 14220 17392
rect 14254 17358 14310 17392
rect 14344 17358 14400 17392
rect 14434 17358 14490 17392
rect 14524 17358 14580 17392
rect 14614 17358 14670 17392
rect 14704 17358 14760 17392
rect 14794 17358 14850 17392
rect 14884 17358 14940 17392
rect 14974 17358 15030 17392
rect 15064 17358 15120 17392
rect 15154 17358 15284 17392
rect 13996 17323 15284 17358
rect 13996 17308 14097 17323
rect 13996 17274 14029 17308
rect 14063 17274 14097 17308
rect 13996 17218 14097 17274
rect 15183 17308 15284 17323
rect 15183 17274 15216 17308
rect 15250 17274 15284 17308
rect 13996 17184 14029 17218
rect 14063 17184 14097 17218
rect 13996 17128 14097 17184
rect 13996 17094 14029 17128
rect 14063 17094 14097 17128
rect 13996 17038 14097 17094
rect 13996 17004 14029 17038
rect 14063 17004 14097 17038
rect 13996 16948 14097 17004
rect 13996 16914 14029 16948
rect 14063 16914 14097 16948
rect 13996 16858 14097 16914
rect 13996 16824 14029 16858
rect 14063 16824 14097 16858
rect 13996 16768 14097 16824
rect 13996 16734 14029 16768
rect 14063 16734 14097 16768
rect 13996 16678 14097 16734
rect 13996 16644 14029 16678
rect 14063 16644 14097 16678
rect 13996 16588 14097 16644
rect 13996 16554 14029 16588
rect 14063 16554 14097 16588
rect 13996 16498 14097 16554
rect 13996 16464 14029 16498
rect 14063 16464 14097 16498
rect 13996 16408 14097 16464
rect 13996 16374 14029 16408
rect 14063 16374 14097 16408
rect 13996 16318 14097 16374
rect 13996 16284 14029 16318
rect 14063 16284 14097 16318
rect 15183 17218 15284 17274
rect 15183 17184 15216 17218
rect 15250 17184 15284 17218
rect 15183 17128 15284 17184
rect 15183 17094 15216 17128
rect 15250 17094 15284 17128
rect 15183 17038 15284 17094
rect 15183 17004 15216 17038
rect 15250 17004 15284 17038
rect 15183 16948 15284 17004
rect 15183 16914 15216 16948
rect 15250 16914 15284 16948
rect 15183 16858 15284 16914
rect 15183 16824 15216 16858
rect 15250 16824 15284 16858
rect 15183 16768 15284 16824
rect 15183 16734 15216 16768
rect 15250 16734 15284 16768
rect 15183 16678 15284 16734
rect 15183 16644 15216 16678
rect 15250 16644 15284 16678
rect 15183 16588 15284 16644
rect 15183 16554 15216 16588
rect 15250 16554 15284 16588
rect 15183 16498 15284 16554
rect 15183 16464 15216 16498
rect 15250 16464 15284 16498
rect 15183 16408 15284 16464
rect 15183 16374 15216 16408
rect 15250 16374 15284 16408
rect 15183 16318 15284 16374
rect 13996 16237 14097 16284
rect 15183 16284 15216 16318
rect 15250 16284 15284 16318
rect 15183 16237 15284 16284
rect 13996 16228 15284 16237
rect 13996 16194 14029 16228
rect 14063 16205 15216 16228
rect 14063 16194 14130 16205
rect 13996 16171 14130 16194
rect 14164 16171 14220 16205
rect 14254 16171 14310 16205
rect 14344 16171 14400 16205
rect 14434 16171 14490 16205
rect 14524 16171 14580 16205
rect 14614 16171 14670 16205
rect 14704 16171 14760 16205
rect 14794 16171 14850 16205
rect 14884 16171 14940 16205
rect 14974 16171 15030 16205
rect 15064 16171 15120 16205
rect 15154 16194 15216 16205
rect 15250 16194 15284 16228
rect 15154 16171 15284 16194
rect 13996 16136 15284 16171
rect 11276 16032 12564 16064
rect 11276 15998 11410 16032
rect 11444 15998 11500 16032
rect 11534 15998 11590 16032
rect 11624 15998 11680 16032
rect 11714 15998 11770 16032
rect 11804 15998 11860 16032
rect 11894 15998 11950 16032
rect 11984 15998 12040 16032
rect 12074 15998 12130 16032
rect 12164 15998 12220 16032
rect 12254 15998 12310 16032
rect 12344 15998 12400 16032
rect 12434 15998 12564 16032
rect 11276 15963 12564 15998
rect 11276 15948 11377 15963
rect 11276 15914 11309 15948
rect 11343 15914 11377 15948
rect 11276 15858 11377 15914
rect 12463 15948 12564 15963
rect 12463 15914 12496 15948
rect 12530 15914 12564 15948
rect 11276 15824 11309 15858
rect 11343 15824 11377 15858
rect 11276 15768 11377 15824
rect 11276 15734 11309 15768
rect 11343 15734 11377 15768
rect 11276 15678 11377 15734
rect 11276 15644 11309 15678
rect 11343 15644 11377 15678
rect 11276 15588 11377 15644
rect 11276 15554 11309 15588
rect 11343 15554 11377 15588
rect 11276 15498 11377 15554
rect 11276 15464 11309 15498
rect 11343 15464 11377 15498
rect 11276 15408 11377 15464
rect 11276 15374 11309 15408
rect 11343 15374 11377 15408
rect 11276 15318 11377 15374
rect 11276 15284 11309 15318
rect 11343 15284 11377 15318
rect 11276 15228 11377 15284
rect 11276 15194 11309 15228
rect 11343 15194 11377 15228
rect 11276 15138 11377 15194
rect 11276 15104 11309 15138
rect 11343 15104 11377 15138
rect 11276 15048 11377 15104
rect 11276 15014 11309 15048
rect 11343 15014 11377 15048
rect 11276 14958 11377 15014
rect 11276 14924 11309 14958
rect 11343 14924 11377 14958
rect 12463 15858 12564 15914
rect 12463 15824 12496 15858
rect 12530 15824 12564 15858
rect 12463 15768 12564 15824
rect 12463 15734 12496 15768
rect 12530 15734 12564 15768
rect 12463 15678 12564 15734
rect 12463 15644 12496 15678
rect 12530 15644 12564 15678
rect 12463 15588 12564 15644
rect 12463 15554 12496 15588
rect 12530 15554 12564 15588
rect 12463 15498 12564 15554
rect 12463 15464 12496 15498
rect 12530 15464 12564 15498
rect 12463 15408 12564 15464
rect 12463 15374 12496 15408
rect 12530 15374 12564 15408
rect 12463 15318 12564 15374
rect 12463 15284 12496 15318
rect 12530 15284 12564 15318
rect 12463 15228 12564 15284
rect 12463 15194 12496 15228
rect 12530 15194 12564 15228
rect 12463 15138 12564 15194
rect 12463 15104 12496 15138
rect 12530 15104 12564 15138
rect 12463 15048 12564 15104
rect 12463 15014 12496 15048
rect 12530 15014 12564 15048
rect 12463 14958 12564 15014
rect 11276 14877 11377 14924
rect 12463 14924 12496 14958
rect 12530 14924 12564 14958
rect 12463 14877 12564 14924
rect 11276 14868 12564 14877
rect 11276 14834 11309 14868
rect 11343 14845 12496 14868
rect 11343 14834 11410 14845
rect 11276 14811 11410 14834
rect 11444 14811 11500 14845
rect 11534 14811 11590 14845
rect 11624 14811 11680 14845
rect 11714 14811 11770 14845
rect 11804 14811 11860 14845
rect 11894 14811 11950 14845
rect 11984 14811 12040 14845
rect 12074 14811 12130 14845
rect 12164 14811 12220 14845
rect 12254 14811 12310 14845
rect 12344 14811 12400 14845
rect 12434 14834 12496 14845
rect 12530 14834 12564 14868
rect 12434 14811 12564 14834
rect 11276 14776 12564 14811
rect 12636 16032 13924 16064
rect 12636 15998 12770 16032
rect 12804 15998 12860 16032
rect 12894 15998 12950 16032
rect 12984 15998 13040 16032
rect 13074 15998 13130 16032
rect 13164 15998 13220 16032
rect 13254 15998 13310 16032
rect 13344 15998 13400 16032
rect 13434 15998 13490 16032
rect 13524 15998 13580 16032
rect 13614 15998 13670 16032
rect 13704 15998 13760 16032
rect 13794 15998 13924 16032
rect 12636 15963 13924 15998
rect 12636 15948 12737 15963
rect 12636 15914 12669 15948
rect 12703 15914 12737 15948
rect 12636 15858 12737 15914
rect 13823 15948 13924 15963
rect 13823 15914 13856 15948
rect 13890 15914 13924 15948
rect 12636 15824 12669 15858
rect 12703 15824 12737 15858
rect 12636 15768 12737 15824
rect 12636 15734 12669 15768
rect 12703 15734 12737 15768
rect 12636 15678 12737 15734
rect 12636 15644 12669 15678
rect 12703 15644 12737 15678
rect 12636 15588 12737 15644
rect 12636 15554 12669 15588
rect 12703 15554 12737 15588
rect 12636 15498 12737 15554
rect 12636 15464 12669 15498
rect 12703 15464 12737 15498
rect 12636 15408 12737 15464
rect 12636 15374 12669 15408
rect 12703 15374 12737 15408
rect 12636 15318 12737 15374
rect 12636 15284 12669 15318
rect 12703 15284 12737 15318
rect 12636 15228 12737 15284
rect 12636 15194 12669 15228
rect 12703 15194 12737 15228
rect 12636 15138 12737 15194
rect 12636 15104 12669 15138
rect 12703 15104 12737 15138
rect 12636 15048 12737 15104
rect 12636 15014 12669 15048
rect 12703 15014 12737 15048
rect 12636 14958 12737 15014
rect 12636 14924 12669 14958
rect 12703 14924 12737 14958
rect 13823 15858 13924 15914
rect 13823 15824 13856 15858
rect 13890 15824 13924 15858
rect 13823 15768 13924 15824
rect 13823 15734 13856 15768
rect 13890 15734 13924 15768
rect 13823 15678 13924 15734
rect 13823 15644 13856 15678
rect 13890 15644 13924 15678
rect 13823 15588 13924 15644
rect 13823 15554 13856 15588
rect 13890 15554 13924 15588
rect 13823 15498 13924 15554
rect 13823 15464 13856 15498
rect 13890 15464 13924 15498
rect 13823 15408 13924 15464
rect 13823 15374 13856 15408
rect 13890 15374 13924 15408
rect 13823 15318 13924 15374
rect 13823 15284 13856 15318
rect 13890 15284 13924 15318
rect 13823 15228 13924 15284
rect 13823 15194 13856 15228
rect 13890 15194 13924 15228
rect 13823 15138 13924 15194
rect 13823 15104 13856 15138
rect 13890 15104 13924 15138
rect 13823 15048 13924 15104
rect 13823 15014 13856 15048
rect 13890 15014 13924 15048
rect 13823 14958 13924 15014
rect 12636 14877 12737 14924
rect 13823 14924 13856 14958
rect 13890 14924 13924 14958
rect 13823 14877 13924 14924
rect 12636 14868 13924 14877
rect 12636 14834 12669 14868
rect 12703 14845 13856 14868
rect 12703 14834 12770 14845
rect 12636 14811 12770 14834
rect 12804 14811 12860 14845
rect 12894 14811 12950 14845
rect 12984 14811 13040 14845
rect 13074 14811 13130 14845
rect 13164 14811 13220 14845
rect 13254 14811 13310 14845
rect 13344 14811 13400 14845
rect 13434 14811 13490 14845
rect 13524 14811 13580 14845
rect 13614 14811 13670 14845
rect 13704 14811 13760 14845
rect 13794 14834 13856 14845
rect 13890 14834 13924 14868
rect 13794 14811 13924 14834
rect 12636 14776 13924 14811
rect 13996 16032 15284 16064
rect 13996 15998 14130 16032
rect 14164 15998 14220 16032
rect 14254 15998 14310 16032
rect 14344 15998 14400 16032
rect 14434 15998 14490 16032
rect 14524 15998 14580 16032
rect 14614 15998 14670 16032
rect 14704 15998 14760 16032
rect 14794 15998 14850 16032
rect 14884 15998 14940 16032
rect 14974 15998 15030 16032
rect 15064 15998 15120 16032
rect 15154 15998 15284 16032
rect 13996 15963 15284 15998
rect 13996 15948 14097 15963
rect 13996 15914 14029 15948
rect 14063 15914 14097 15948
rect 13996 15858 14097 15914
rect 15183 15948 15284 15963
rect 15183 15914 15216 15948
rect 15250 15914 15284 15948
rect 13996 15824 14029 15858
rect 14063 15824 14097 15858
rect 13996 15768 14097 15824
rect 13996 15734 14029 15768
rect 14063 15734 14097 15768
rect 13996 15678 14097 15734
rect 13996 15644 14029 15678
rect 14063 15644 14097 15678
rect 13996 15588 14097 15644
rect 13996 15554 14029 15588
rect 14063 15554 14097 15588
rect 13996 15498 14097 15554
rect 13996 15464 14029 15498
rect 14063 15464 14097 15498
rect 13996 15408 14097 15464
rect 13996 15374 14029 15408
rect 14063 15374 14097 15408
rect 13996 15318 14097 15374
rect 13996 15284 14029 15318
rect 14063 15284 14097 15318
rect 13996 15228 14097 15284
rect 13996 15194 14029 15228
rect 14063 15194 14097 15228
rect 13996 15138 14097 15194
rect 13996 15104 14029 15138
rect 14063 15104 14097 15138
rect 13996 15048 14097 15104
rect 13996 15014 14029 15048
rect 14063 15014 14097 15048
rect 13996 14958 14097 15014
rect 13996 14924 14029 14958
rect 14063 14924 14097 14958
rect 15183 15858 15284 15914
rect 15183 15824 15216 15858
rect 15250 15824 15284 15858
rect 15183 15768 15284 15824
rect 15183 15734 15216 15768
rect 15250 15734 15284 15768
rect 15183 15678 15284 15734
rect 15183 15644 15216 15678
rect 15250 15644 15284 15678
rect 15183 15588 15284 15644
rect 15183 15554 15216 15588
rect 15250 15554 15284 15588
rect 15183 15498 15284 15554
rect 15183 15464 15216 15498
rect 15250 15464 15284 15498
rect 15183 15408 15284 15464
rect 15183 15374 15216 15408
rect 15250 15374 15284 15408
rect 15183 15318 15284 15374
rect 15183 15284 15216 15318
rect 15250 15284 15284 15318
rect 15183 15228 15284 15284
rect 15183 15194 15216 15228
rect 15250 15194 15284 15228
rect 15183 15138 15284 15194
rect 15183 15104 15216 15138
rect 15250 15104 15284 15138
rect 15183 15048 15284 15104
rect 15183 15014 15216 15048
rect 15250 15014 15284 15048
rect 15183 14958 15284 15014
rect 13996 14877 14097 14924
rect 15183 14924 15216 14958
rect 15250 14924 15284 14958
rect 15183 14877 15284 14924
rect 13996 14868 15284 14877
rect 13996 14834 14029 14868
rect 14063 14845 15216 14868
rect 14063 14834 14130 14845
rect 13996 14811 14130 14834
rect 14164 14811 14220 14845
rect 14254 14811 14310 14845
rect 14344 14811 14400 14845
rect 14434 14811 14490 14845
rect 14524 14811 14580 14845
rect 14614 14811 14670 14845
rect 14704 14811 14760 14845
rect 14794 14811 14850 14845
rect 14884 14811 14940 14845
rect 14974 14811 15030 14845
rect 15064 14811 15120 14845
rect 15154 14834 15216 14845
rect 15250 14834 15284 14868
rect 15154 14811 15284 14834
rect 13996 14776 15284 14811
rect 15400 14250 15480 14280
rect 15400 14210 15420 14250
rect 15460 14210 15480 14250
rect 15400 14150 15480 14210
rect 15400 14110 15420 14150
rect 15460 14110 15480 14150
rect 15400 14080 15480 14110
rect 11900 13640 11980 13670
rect 11900 13600 11920 13640
rect 11960 13600 11980 13640
rect 11900 13540 11980 13600
rect 11900 13500 11920 13540
rect 11960 13500 11980 13540
rect 11900 13440 11980 13500
rect 11900 13400 11920 13440
rect 11960 13400 11980 13440
rect 11900 13340 11980 13400
rect 11900 13300 11920 13340
rect 11960 13300 11980 13340
rect 11900 13240 11980 13300
rect 11900 13200 11920 13240
rect 11960 13200 11980 13240
rect 11900 13170 11980 13200
rect 14580 13640 14660 13670
rect 14580 13600 14600 13640
rect 14640 13600 14660 13640
rect 14580 13540 14660 13600
rect 14580 13500 14600 13540
rect 14640 13500 14660 13540
rect 14580 13440 14660 13500
rect 14580 13400 14600 13440
rect 14640 13400 14660 13440
rect 14580 13340 14660 13400
rect 14580 13300 14600 13340
rect 14640 13300 14660 13340
rect 14580 13240 14660 13300
rect 14580 13200 14600 13240
rect 14640 13200 14660 13240
rect 14580 13170 14660 13200
rect 12800 12720 12880 12750
rect 12800 12680 12820 12720
rect 12860 12680 12880 12720
rect 12800 12640 12880 12680
rect 12800 12600 12820 12640
rect 12860 12600 12880 12640
rect 12800 12560 12880 12600
rect 12800 12520 12820 12560
rect 12860 12520 12880 12560
rect 12800 12490 12880 12520
rect 13680 12720 13760 12750
rect 13680 12680 13700 12720
rect 13740 12680 13760 12720
rect 13680 12640 13760 12680
rect 13680 12600 13700 12640
rect 13740 12600 13760 12640
rect 13680 12560 13760 12600
rect 13680 12520 13700 12560
rect 13740 12520 13760 12560
rect 13680 12490 13760 12520
<< nsubdiff >>
rect 8263 18563 8359 18597
rect 8619 18563 8715 18597
rect 8263 18501 8297 18563
rect 8681 18501 8715 18563
rect 8263 17111 8297 17173
rect 8681 17111 8715 17173
rect 8263 17077 8359 17111
rect 8619 17077 8715 17111
rect 9050 18566 9146 18600
rect 9738 18566 9834 18600
rect 9050 18504 9084 18566
rect 9800 18504 9834 18566
rect 9050 16712 9084 16774
rect 9800 16712 9834 16774
rect 9050 16678 9146 16712
rect 9738 16678 9834 16712
rect 10163 18563 10259 18597
rect 10851 18563 10947 18597
rect 10163 18501 10197 18563
rect 10913 18501 10947 18563
rect 10163 16181 10197 16243
rect 11439 18602 12401 18621
rect 11439 18568 11550 18602
rect 11584 18568 11640 18602
rect 11674 18568 11730 18602
rect 11764 18568 11820 18602
rect 11854 18568 11910 18602
rect 11944 18568 12000 18602
rect 12034 18568 12090 18602
rect 12124 18568 12180 18602
rect 12214 18568 12270 18602
rect 12304 18568 12401 18602
rect 11439 18549 12401 18568
rect 11439 18508 11511 18549
rect 11439 18474 11458 18508
rect 11492 18474 11511 18508
rect 12329 18489 12401 18549
rect 11439 18418 11511 18474
rect 11439 18384 11458 18418
rect 11492 18384 11511 18418
rect 11439 18328 11511 18384
rect 11439 18294 11458 18328
rect 11492 18294 11511 18328
rect 11439 18238 11511 18294
rect 11439 18204 11458 18238
rect 11492 18204 11511 18238
rect 11439 18148 11511 18204
rect 11439 18114 11458 18148
rect 11492 18114 11511 18148
rect 11439 18058 11511 18114
rect 11439 18024 11458 18058
rect 11492 18024 11511 18058
rect 11439 17968 11511 18024
rect 11439 17934 11458 17968
rect 11492 17934 11511 17968
rect 11439 17878 11511 17934
rect 11439 17844 11458 17878
rect 11492 17844 11511 17878
rect 11439 17788 11511 17844
rect 12329 18455 12348 18489
rect 12382 18455 12401 18489
rect 12329 18399 12401 18455
rect 12329 18365 12348 18399
rect 12382 18365 12401 18399
rect 12329 18309 12401 18365
rect 12329 18275 12348 18309
rect 12382 18275 12401 18309
rect 12329 18219 12401 18275
rect 12329 18185 12348 18219
rect 12382 18185 12401 18219
rect 12329 18129 12401 18185
rect 12329 18095 12348 18129
rect 12382 18095 12401 18129
rect 12329 18039 12401 18095
rect 12329 18005 12348 18039
rect 12382 18005 12401 18039
rect 12329 17949 12401 18005
rect 12329 17915 12348 17949
rect 12382 17915 12401 17949
rect 12329 17859 12401 17915
rect 12329 17825 12348 17859
rect 12382 17825 12401 17859
rect 11439 17754 11458 17788
rect 11492 17754 11511 17788
rect 11439 17731 11511 17754
rect 12329 17769 12401 17825
rect 12329 17735 12348 17769
rect 12382 17735 12401 17769
rect 12329 17731 12401 17735
rect 11439 17712 12401 17731
rect 11439 17678 11516 17712
rect 11550 17678 11606 17712
rect 11640 17678 11696 17712
rect 11730 17678 11786 17712
rect 11820 17678 11876 17712
rect 11910 17678 11966 17712
rect 12000 17678 12056 17712
rect 12090 17678 12146 17712
rect 12180 17678 12236 17712
rect 12270 17678 12401 17712
rect 11439 17659 12401 17678
rect 12799 18602 13761 18621
rect 12799 18568 12910 18602
rect 12944 18568 13000 18602
rect 13034 18568 13090 18602
rect 13124 18568 13180 18602
rect 13214 18568 13270 18602
rect 13304 18568 13360 18602
rect 13394 18568 13450 18602
rect 13484 18568 13540 18602
rect 13574 18568 13630 18602
rect 13664 18568 13761 18602
rect 12799 18549 13761 18568
rect 12799 18508 12871 18549
rect 12799 18474 12818 18508
rect 12852 18474 12871 18508
rect 13689 18489 13761 18549
rect 12799 18418 12871 18474
rect 12799 18384 12818 18418
rect 12852 18384 12871 18418
rect 12799 18328 12871 18384
rect 12799 18294 12818 18328
rect 12852 18294 12871 18328
rect 12799 18238 12871 18294
rect 12799 18204 12818 18238
rect 12852 18204 12871 18238
rect 12799 18148 12871 18204
rect 12799 18114 12818 18148
rect 12852 18114 12871 18148
rect 12799 18058 12871 18114
rect 12799 18024 12818 18058
rect 12852 18024 12871 18058
rect 12799 17968 12871 18024
rect 12799 17934 12818 17968
rect 12852 17934 12871 17968
rect 12799 17878 12871 17934
rect 12799 17844 12818 17878
rect 12852 17844 12871 17878
rect 12799 17788 12871 17844
rect 13689 18455 13708 18489
rect 13742 18455 13761 18489
rect 13689 18399 13761 18455
rect 13689 18365 13708 18399
rect 13742 18365 13761 18399
rect 13689 18309 13761 18365
rect 13689 18275 13708 18309
rect 13742 18275 13761 18309
rect 13689 18219 13761 18275
rect 13689 18185 13708 18219
rect 13742 18185 13761 18219
rect 13689 18129 13761 18185
rect 13689 18095 13708 18129
rect 13742 18095 13761 18129
rect 13689 18039 13761 18095
rect 13689 18005 13708 18039
rect 13742 18005 13761 18039
rect 13689 17949 13761 18005
rect 13689 17915 13708 17949
rect 13742 17915 13761 17949
rect 13689 17859 13761 17915
rect 13689 17825 13708 17859
rect 13742 17825 13761 17859
rect 12799 17754 12818 17788
rect 12852 17754 12871 17788
rect 12799 17731 12871 17754
rect 13689 17769 13761 17825
rect 13689 17735 13708 17769
rect 13742 17735 13761 17769
rect 13689 17731 13761 17735
rect 12799 17712 13761 17731
rect 12799 17678 12876 17712
rect 12910 17678 12966 17712
rect 13000 17678 13056 17712
rect 13090 17678 13146 17712
rect 13180 17678 13236 17712
rect 13270 17678 13326 17712
rect 13360 17678 13416 17712
rect 13450 17678 13506 17712
rect 13540 17678 13596 17712
rect 13630 17678 13761 17712
rect 12799 17659 13761 17678
rect 14159 18602 15121 18621
rect 14159 18568 14270 18602
rect 14304 18568 14360 18602
rect 14394 18568 14450 18602
rect 14484 18568 14540 18602
rect 14574 18568 14630 18602
rect 14664 18568 14720 18602
rect 14754 18568 14810 18602
rect 14844 18568 14900 18602
rect 14934 18568 14990 18602
rect 15024 18568 15121 18602
rect 14159 18549 15121 18568
rect 14159 18508 14231 18549
rect 14159 18474 14178 18508
rect 14212 18474 14231 18508
rect 15049 18489 15121 18549
rect 14159 18418 14231 18474
rect 14159 18384 14178 18418
rect 14212 18384 14231 18418
rect 14159 18328 14231 18384
rect 14159 18294 14178 18328
rect 14212 18294 14231 18328
rect 14159 18238 14231 18294
rect 14159 18204 14178 18238
rect 14212 18204 14231 18238
rect 14159 18148 14231 18204
rect 14159 18114 14178 18148
rect 14212 18114 14231 18148
rect 14159 18058 14231 18114
rect 14159 18024 14178 18058
rect 14212 18024 14231 18058
rect 14159 17968 14231 18024
rect 14159 17934 14178 17968
rect 14212 17934 14231 17968
rect 14159 17878 14231 17934
rect 14159 17844 14178 17878
rect 14212 17844 14231 17878
rect 14159 17788 14231 17844
rect 15049 18455 15068 18489
rect 15102 18455 15121 18489
rect 15049 18399 15121 18455
rect 15049 18365 15068 18399
rect 15102 18365 15121 18399
rect 15049 18309 15121 18365
rect 15049 18275 15068 18309
rect 15102 18275 15121 18309
rect 15049 18219 15121 18275
rect 15049 18185 15068 18219
rect 15102 18185 15121 18219
rect 15049 18129 15121 18185
rect 15049 18095 15068 18129
rect 15102 18095 15121 18129
rect 15049 18039 15121 18095
rect 15049 18005 15068 18039
rect 15102 18005 15121 18039
rect 15049 17949 15121 18005
rect 15049 17915 15068 17949
rect 15102 17915 15121 17949
rect 15049 17859 15121 17915
rect 15049 17825 15068 17859
rect 15102 17825 15121 17859
rect 14159 17754 14178 17788
rect 14212 17754 14231 17788
rect 14159 17731 14231 17754
rect 15049 17769 15121 17825
rect 15049 17735 15068 17769
rect 15102 17735 15121 17769
rect 15049 17731 15121 17735
rect 14159 17712 15121 17731
rect 14159 17678 14236 17712
rect 14270 17678 14326 17712
rect 14360 17678 14416 17712
rect 14450 17678 14506 17712
rect 14540 17678 14596 17712
rect 14630 17678 14686 17712
rect 14720 17678 14776 17712
rect 14810 17678 14866 17712
rect 14900 17678 14956 17712
rect 14990 17678 15121 17712
rect 14159 17659 15121 17678
rect 15483 18563 15579 18597
rect 16171 18563 16267 18597
rect 15483 18501 15517 18563
rect 10913 16181 10947 16243
rect 10163 16147 10259 16181
rect 10851 16147 10947 16181
rect 11439 17242 12401 17261
rect 11439 17208 11550 17242
rect 11584 17208 11640 17242
rect 11674 17208 11730 17242
rect 11764 17208 11820 17242
rect 11854 17208 11910 17242
rect 11944 17208 12000 17242
rect 12034 17208 12090 17242
rect 12124 17208 12180 17242
rect 12214 17208 12270 17242
rect 12304 17208 12401 17242
rect 11439 17189 12401 17208
rect 11439 17148 11511 17189
rect 11439 17114 11458 17148
rect 11492 17114 11511 17148
rect 12329 17129 12401 17189
rect 11439 17058 11511 17114
rect 11439 17024 11458 17058
rect 11492 17024 11511 17058
rect 11439 16968 11511 17024
rect 11439 16934 11458 16968
rect 11492 16934 11511 16968
rect 11439 16878 11511 16934
rect 11439 16844 11458 16878
rect 11492 16844 11511 16878
rect 11439 16788 11511 16844
rect 11439 16754 11458 16788
rect 11492 16754 11511 16788
rect 11439 16698 11511 16754
rect 11439 16664 11458 16698
rect 11492 16664 11511 16698
rect 11439 16608 11511 16664
rect 11439 16574 11458 16608
rect 11492 16574 11511 16608
rect 11439 16518 11511 16574
rect 11439 16484 11458 16518
rect 11492 16484 11511 16518
rect 11439 16428 11511 16484
rect 12329 17095 12348 17129
rect 12382 17095 12401 17129
rect 12329 17039 12401 17095
rect 12329 17005 12348 17039
rect 12382 17005 12401 17039
rect 12329 16949 12401 17005
rect 12329 16915 12348 16949
rect 12382 16915 12401 16949
rect 12329 16859 12401 16915
rect 12329 16825 12348 16859
rect 12382 16825 12401 16859
rect 12329 16769 12401 16825
rect 12329 16735 12348 16769
rect 12382 16735 12401 16769
rect 12329 16679 12401 16735
rect 12329 16645 12348 16679
rect 12382 16645 12401 16679
rect 12329 16589 12401 16645
rect 12329 16555 12348 16589
rect 12382 16555 12401 16589
rect 12329 16499 12401 16555
rect 12329 16465 12348 16499
rect 12382 16465 12401 16499
rect 11439 16394 11458 16428
rect 11492 16394 11511 16428
rect 11439 16371 11511 16394
rect 12329 16409 12401 16465
rect 12329 16375 12348 16409
rect 12382 16375 12401 16409
rect 12329 16371 12401 16375
rect 11439 16352 12401 16371
rect 11439 16318 11516 16352
rect 11550 16318 11606 16352
rect 11640 16318 11696 16352
rect 11730 16318 11786 16352
rect 11820 16318 11876 16352
rect 11910 16318 11966 16352
rect 12000 16318 12056 16352
rect 12090 16318 12146 16352
rect 12180 16318 12236 16352
rect 12270 16318 12401 16352
rect 11439 16299 12401 16318
rect 12799 17242 13761 17261
rect 12799 17208 12910 17242
rect 12944 17208 13000 17242
rect 13034 17208 13090 17242
rect 13124 17208 13180 17242
rect 13214 17208 13270 17242
rect 13304 17208 13360 17242
rect 13394 17208 13450 17242
rect 13484 17208 13540 17242
rect 13574 17208 13630 17242
rect 13664 17208 13761 17242
rect 12799 17189 13761 17208
rect 12799 17148 12871 17189
rect 12799 17114 12818 17148
rect 12852 17114 12871 17148
rect 13689 17129 13761 17189
rect 12799 17058 12871 17114
rect 12799 17024 12818 17058
rect 12852 17024 12871 17058
rect 12799 16968 12871 17024
rect 12799 16934 12818 16968
rect 12852 16934 12871 16968
rect 12799 16878 12871 16934
rect 12799 16844 12818 16878
rect 12852 16844 12871 16878
rect 12799 16788 12871 16844
rect 12799 16754 12818 16788
rect 12852 16754 12871 16788
rect 12799 16698 12871 16754
rect 12799 16664 12818 16698
rect 12852 16664 12871 16698
rect 12799 16608 12871 16664
rect 12799 16574 12818 16608
rect 12852 16574 12871 16608
rect 12799 16518 12871 16574
rect 12799 16484 12818 16518
rect 12852 16484 12871 16518
rect 12799 16428 12871 16484
rect 13689 17095 13708 17129
rect 13742 17095 13761 17129
rect 13689 17039 13761 17095
rect 13689 17005 13708 17039
rect 13742 17005 13761 17039
rect 13689 16949 13761 17005
rect 13689 16915 13708 16949
rect 13742 16915 13761 16949
rect 13689 16859 13761 16915
rect 13689 16825 13708 16859
rect 13742 16825 13761 16859
rect 13689 16769 13761 16825
rect 13689 16735 13708 16769
rect 13742 16735 13761 16769
rect 13689 16679 13761 16735
rect 13689 16645 13708 16679
rect 13742 16645 13761 16679
rect 13689 16589 13761 16645
rect 13689 16555 13708 16589
rect 13742 16555 13761 16589
rect 13689 16499 13761 16555
rect 13689 16465 13708 16499
rect 13742 16465 13761 16499
rect 12799 16394 12818 16428
rect 12852 16394 12871 16428
rect 12799 16371 12871 16394
rect 13689 16409 13761 16465
rect 13689 16375 13708 16409
rect 13742 16375 13761 16409
rect 13689 16371 13761 16375
rect 12799 16352 13761 16371
rect 12799 16318 12876 16352
rect 12910 16318 12966 16352
rect 13000 16318 13056 16352
rect 13090 16318 13146 16352
rect 13180 16318 13236 16352
rect 13270 16318 13326 16352
rect 13360 16318 13416 16352
rect 13450 16318 13506 16352
rect 13540 16318 13596 16352
rect 13630 16318 13761 16352
rect 12799 16299 13761 16318
rect 14159 17242 15121 17261
rect 14159 17208 14270 17242
rect 14304 17208 14360 17242
rect 14394 17208 14450 17242
rect 14484 17208 14540 17242
rect 14574 17208 14630 17242
rect 14664 17208 14720 17242
rect 14754 17208 14810 17242
rect 14844 17208 14900 17242
rect 14934 17208 14990 17242
rect 15024 17208 15121 17242
rect 14159 17189 15121 17208
rect 14159 17148 14231 17189
rect 14159 17114 14178 17148
rect 14212 17114 14231 17148
rect 15049 17129 15121 17189
rect 14159 17058 14231 17114
rect 14159 17024 14178 17058
rect 14212 17024 14231 17058
rect 14159 16968 14231 17024
rect 14159 16934 14178 16968
rect 14212 16934 14231 16968
rect 14159 16878 14231 16934
rect 14159 16844 14178 16878
rect 14212 16844 14231 16878
rect 14159 16788 14231 16844
rect 14159 16754 14178 16788
rect 14212 16754 14231 16788
rect 14159 16698 14231 16754
rect 14159 16664 14178 16698
rect 14212 16664 14231 16698
rect 14159 16608 14231 16664
rect 14159 16574 14178 16608
rect 14212 16574 14231 16608
rect 14159 16518 14231 16574
rect 14159 16484 14178 16518
rect 14212 16484 14231 16518
rect 14159 16428 14231 16484
rect 15049 17095 15068 17129
rect 15102 17095 15121 17129
rect 15049 17039 15121 17095
rect 15049 17005 15068 17039
rect 15102 17005 15121 17039
rect 15049 16949 15121 17005
rect 15049 16915 15068 16949
rect 15102 16915 15121 16949
rect 15049 16859 15121 16915
rect 15049 16825 15068 16859
rect 15102 16825 15121 16859
rect 15049 16769 15121 16825
rect 15049 16735 15068 16769
rect 15102 16735 15121 16769
rect 15049 16679 15121 16735
rect 15049 16645 15068 16679
rect 15102 16645 15121 16679
rect 15049 16589 15121 16645
rect 15049 16555 15068 16589
rect 15102 16555 15121 16589
rect 15049 16499 15121 16555
rect 15049 16465 15068 16499
rect 15102 16465 15121 16499
rect 14159 16394 14178 16428
rect 14212 16394 14231 16428
rect 14159 16371 14231 16394
rect 15049 16409 15121 16465
rect 15049 16375 15068 16409
rect 15102 16375 15121 16409
rect 15049 16371 15121 16375
rect 14159 16352 15121 16371
rect 14159 16318 14236 16352
rect 14270 16318 14326 16352
rect 14360 16318 14416 16352
rect 14450 16318 14506 16352
rect 14540 16318 14596 16352
rect 14630 16318 14686 16352
rect 14720 16318 14776 16352
rect 14810 16318 14866 16352
rect 14900 16318 14956 16352
rect 14990 16318 15121 16352
rect 14159 16299 15121 16318
rect 16233 18501 16267 18563
rect 15483 16181 15517 16243
rect 16596 18560 16692 18594
rect 16952 18560 17048 18594
rect 16596 18498 16630 18560
rect 17014 18498 17048 18560
rect 16596 17318 16630 17380
rect 17014 17318 17048 17380
rect 16596 17284 16692 17318
rect 16952 17284 17048 17318
rect 17383 18563 17479 18597
rect 17739 18563 17835 18597
rect 17383 18501 17417 18563
rect 17801 18501 17835 18563
rect 17383 17111 17417 17173
rect 17801 17111 17835 17173
rect 17383 17077 17479 17111
rect 17739 17077 17835 17111
rect 16233 16181 16267 16243
rect 15483 16147 15579 16181
rect 16171 16147 16267 16181
rect 11439 15882 12401 15901
rect 11439 15848 11550 15882
rect 11584 15848 11640 15882
rect 11674 15848 11730 15882
rect 11764 15848 11820 15882
rect 11854 15848 11910 15882
rect 11944 15848 12000 15882
rect 12034 15848 12090 15882
rect 12124 15848 12180 15882
rect 12214 15848 12270 15882
rect 12304 15848 12401 15882
rect 11439 15829 12401 15848
rect 11439 15788 11511 15829
rect 11439 15754 11458 15788
rect 11492 15754 11511 15788
rect 12329 15769 12401 15829
rect 11439 15698 11511 15754
rect 11439 15664 11458 15698
rect 11492 15664 11511 15698
rect 11439 15608 11511 15664
rect 11439 15574 11458 15608
rect 11492 15574 11511 15608
rect 11439 15518 11511 15574
rect 11439 15484 11458 15518
rect 11492 15484 11511 15518
rect 11439 15428 11511 15484
rect 11439 15394 11458 15428
rect 11492 15394 11511 15428
rect 11439 15338 11511 15394
rect 11439 15304 11458 15338
rect 11492 15304 11511 15338
rect 11439 15248 11511 15304
rect 11439 15214 11458 15248
rect 11492 15214 11511 15248
rect 11439 15158 11511 15214
rect 11439 15124 11458 15158
rect 11492 15124 11511 15158
rect 11439 15068 11511 15124
rect 12329 15735 12348 15769
rect 12382 15735 12401 15769
rect 12329 15679 12401 15735
rect 12329 15645 12348 15679
rect 12382 15645 12401 15679
rect 12329 15589 12401 15645
rect 12329 15555 12348 15589
rect 12382 15555 12401 15589
rect 12329 15499 12401 15555
rect 12329 15465 12348 15499
rect 12382 15465 12401 15499
rect 12329 15409 12401 15465
rect 12329 15375 12348 15409
rect 12382 15375 12401 15409
rect 12329 15319 12401 15375
rect 12329 15285 12348 15319
rect 12382 15285 12401 15319
rect 12329 15229 12401 15285
rect 12329 15195 12348 15229
rect 12382 15195 12401 15229
rect 12329 15139 12401 15195
rect 12329 15105 12348 15139
rect 12382 15105 12401 15139
rect 11439 15034 11458 15068
rect 11492 15034 11511 15068
rect 11439 15011 11511 15034
rect 12329 15049 12401 15105
rect 12329 15015 12348 15049
rect 12382 15015 12401 15049
rect 12329 15011 12401 15015
rect 11439 14992 12401 15011
rect 11439 14958 11516 14992
rect 11550 14958 11606 14992
rect 11640 14958 11696 14992
rect 11730 14958 11786 14992
rect 11820 14958 11876 14992
rect 11910 14958 11966 14992
rect 12000 14958 12056 14992
rect 12090 14958 12146 14992
rect 12180 14958 12236 14992
rect 12270 14958 12401 14992
rect 11439 14939 12401 14958
rect 12799 15882 13761 15901
rect 12799 15848 12910 15882
rect 12944 15848 13000 15882
rect 13034 15848 13090 15882
rect 13124 15848 13180 15882
rect 13214 15848 13270 15882
rect 13304 15848 13360 15882
rect 13394 15848 13450 15882
rect 13484 15848 13540 15882
rect 13574 15848 13630 15882
rect 13664 15848 13761 15882
rect 12799 15829 13761 15848
rect 12799 15788 12871 15829
rect 12799 15754 12818 15788
rect 12852 15754 12871 15788
rect 13689 15769 13761 15829
rect 12799 15698 12871 15754
rect 12799 15664 12818 15698
rect 12852 15664 12871 15698
rect 12799 15608 12871 15664
rect 12799 15574 12818 15608
rect 12852 15574 12871 15608
rect 12799 15518 12871 15574
rect 12799 15484 12818 15518
rect 12852 15484 12871 15518
rect 12799 15428 12871 15484
rect 12799 15394 12818 15428
rect 12852 15394 12871 15428
rect 12799 15338 12871 15394
rect 12799 15304 12818 15338
rect 12852 15304 12871 15338
rect 12799 15248 12871 15304
rect 12799 15214 12818 15248
rect 12852 15214 12871 15248
rect 12799 15158 12871 15214
rect 12799 15124 12818 15158
rect 12852 15124 12871 15158
rect 12799 15068 12871 15124
rect 13689 15735 13708 15769
rect 13742 15735 13761 15769
rect 13689 15679 13761 15735
rect 13689 15645 13708 15679
rect 13742 15645 13761 15679
rect 13689 15589 13761 15645
rect 13689 15555 13708 15589
rect 13742 15555 13761 15589
rect 13689 15499 13761 15555
rect 13689 15465 13708 15499
rect 13742 15465 13761 15499
rect 13689 15409 13761 15465
rect 13689 15375 13708 15409
rect 13742 15375 13761 15409
rect 13689 15319 13761 15375
rect 13689 15285 13708 15319
rect 13742 15285 13761 15319
rect 13689 15229 13761 15285
rect 13689 15195 13708 15229
rect 13742 15195 13761 15229
rect 13689 15139 13761 15195
rect 13689 15105 13708 15139
rect 13742 15105 13761 15139
rect 12799 15034 12818 15068
rect 12852 15034 12871 15068
rect 12799 15011 12871 15034
rect 13689 15049 13761 15105
rect 13689 15015 13708 15049
rect 13742 15015 13761 15049
rect 13689 15011 13761 15015
rect 12799 14992 13761 15011
rect 12799 14958 12876 14992
rect 12910 14958 12966 14992
rect 13000 14958 13056 14992
rect 13090 14958 13146 14992
rect 13180 14958 13236 14992
rect 13270 14958 13326 14992
rect 13360 14958 13416 14992
rect 13450 14958 13506 14992
rect 13540 14958 13596 14992
rect 13630 14958 13761 14992
rect 12799 14939 13761 14958
rect 14159 15882 15121 15901
rect 14159 15848 14270 15882
rect 14304 15848 14360 15882
rect 14394 15848 14450 15882
rect 14484 15848 14540 15882
rect 14574 15848 14630 15882
rect 14664 15848 14720 15882
rect 14754 15848 14810 15882
rect 14844 15848 14900 15882
rect 14934 15848 14990 15882
rect 15024 15848 15121 15882
rect 14159 15829 15121 15848
rect 14159 15788 14231 15829
rect 14159 15754 14178 15788
rect 14212 15754 14231 15788
rect 15049 15769 15121 15829
rect 14159 15698 14231 15754
rect 14159 15664 14178 15698
rect 14212 15664 14231 15698
rect 14159 15608 14231 15664
rect 14159 15574 14178 15608
rect 14212 15574 14231 15608
rect 14159 15518 14231 15574
rect 14159 15484 14178 15518
rect 14212 15484 14231 15518
rect 14159 15428 14231 15484
rect 14159 15394 14178 15428
rect 14212 15394 14231 15428
rect 14159 15338 14231 15394
rect 14159 15304 14178 15338
rect 14212 15304 14231 15338
rect 14159 15248 14231 15304
rect 14159 15214 14178 15248
rect 14212 15214 14231 15248
rect 14159 15158 14231 15214
rect 14159 15124 14178 15158
rect 14212 15124 14231 15158
rect 14159 15068 14231 15124
rect 15049 15735 15068 15769
rect 15102 15735 15121 15769
rect 15049 15679 15121 15735
rect 15049 15645 15068 15679
rect 15102 15645 15121 15679
rect 15049 15589 15121 15645
rect 15049 15555 15068 15589
rect 15102 15555 15121 15589
rect 15049 15499 15121 15555
rect 15049 15465 15068 15499
rect 15102 15465 15121 15499
rect 15049 15409 15121 15465
rect 15049 15375 15068 15409
rect 15102 15375 15121 15409
rect 15049 15319 15121 15375
rect 15049 15285 15068 15319
rect 15102 15285 15121 15319
rect 15049 15229 15121 15285
rect 15049 15195 15068 15229
rect 15102 15195 15121 15229
rect 15049 15139 15121 15195
rect 15049 15105 15068 15139
rect 15102 15105 15121 15139
rect 14159 15034 14178 15068
rect 14212 15034 14231 15068
rect 14159 15011 14231 15034
rect 15049 15049 15121 15105
rect 15049 15015 15068 15049
rect 15102 15015 15121 15049
rect 15049 15011 15121 15015
rect 14159 14992 15121 15011
rect 14159 14958 14236 14992
rect 14270 14958 14326 14992
rect 14360 14958 14416 14992
rect 14450 14958 14506 14992
rect 14540 14958 14596 14992
rect 14630 14958 14686 14992
rect 14720 14958 14776 14992
rect 14810 14958 14866 14992
rect 14900 14958 14956 14992
rect 14990 14958 15121 14992
rect 14159 14939 15121 14958
rect 10440 11790 10520 11820
rect 10440 11750 10460 11790
rect 10500 11750 10520 11790
rect 10440 11690 10520 11750
rect 10440 11650 10460 11690
rect 10500 11650 10520 11690
rect 10440 11620 10520 11650
rect 13000 11790 13080 11820
rect 13000 11750 13020 11790
rect 13060 11750 13080 11790
rect 13000 11690 13080 11750
rect 13000 11650 13020 11690
rect 13060 11650 13080 11690
rect 13000 11620 13080 11650
rect 13480 11790 13560 11820
rect 13480 11750 13500 11790
rect 13540 11750 13560 11790
rect 13480 11690 13560 11750
rect 13480 11650 13500 11690
rect 13540 11650 13560 11690
rect 13480 11620 13560 11650
rect 16040 11790 16120 11820
rect 16040 11750 16060 11790
rect 16100 11750 16120 11790
rect 16040 11690 16120 11750
rect 16040 11650 16060 11690
rect 16100 11650 16120 11690
rect 16040 11620 16120 11650
rect 11540 10630 11620 10660
rect 11540 10590 11560 10630
rect 11600 10590 11620 10630
rect 11540 10530 11620 10590
rect 11540 10490 11560 10530
rect 11600 10490 11620 10530
rect 11540 10430 11620 10490
rect 11540 10390 11560 10430
rect 11600 10390 11620 10430
rect 11540 10330 11620 10390
rect 11540 10290 11560 10330
rect 11600 10290 11620 10330
rect 11540 10230 11620 10290
rect 11540 10190 11560 10230
rect 11600 10190 11620 10230
rect 11540 10130 11620 10190
rect 11540 10090 11560 10130
rect 11600 10090 11620 10130
rect 11540 10060 11620 10090
rect 14940 10630 15020 10660
rect 14940 10590 14960 10630
rect 15000 10590 15020 10630
rect 14940 10530 15020 10590
rect 14940 10490 14960 10530
rect 15000 10490 15020 10530
rect 14940 10430 15020 10490
rect 14940 10390 14960 10430
rect 15000 10390 15020 10430
rect 14940 10330 15020 10390
rect 14940 10290 14960 10330
rect 15000 10290 15020 10330
rect 14940 10230 15020 10290
rect 15400 10430 15480 10460
rect 15400 10390 15420 10430
rect 15460 10390 15480 10430
rect 15400 10330 15480 10390
rect 15400 10290 15420 10330
rect 15460 10290 15480 10330
rect 15400 10260 15480 10290
rect 16010 10430 16090 10460
rect 16010 10390 16030 10430
rect 16070 10390 16090 10430
rect 16010 10330 16090 10390
rect 16010 10290 16030 10330
rect 16070 10290 16090 10330
rect 16010 10260 16090 10290
rect 14940 10190 14960 10230
rect 15000 10190 15020 10230
rect 14940 10130 15020 10190
rect 14940 10090 14960 10130
rect 15000 10090 15020 10130
rect 14940 10060 15020 10090
rect 11550 9630 11630 9660
rect 11550 9590 11570 9630
rect 11610 9590 11630 9630
rect 11550 9530 11630 9590
rect 11550 9490 11570 9530
rect 11610 9490 11630 9530
rect 11550 9460 11630 9490
rect 13030 9630 13110 9660
rect 13030 9590 13050 9630
rect 13090 9590 13110 9630
rect 13030 9530 13110 9590
rect 13030 9490 13050 9530
rect 13090 9490 13110 9530
rect 13030 9460 13110 9490
rect 13450 9630 13530 9660
rect 13450 9590 13470 9630
rect 13510 9590 13530 9630
rect 13450 9530 13530 9590
rect 13450 9490 13470 9530
rect 13510 9490 13530 9530
rect 13450 9460 13530 9490
rect 14930 9630 15010 9660
rect 14930 9590 14950 9630
rect 14990 9590 15010 9630
rect 14930 9530 15010 9590
rect 14930 9490 14950 9530
rect 14990 9490 15010 9530
rect 14930 9460 15010 9490
<< psubdiffcont >>
rect 13260 19030 13300 19070
rect 13260 18950 13300 18990
rect 13260 18870 13300 18910
rect 11410 18718 11444 18752
rect 11500 18718 11534 18752
rect 11590 18718 11624 18752
rect 11680 18718 11714 18752
rect 11770 18718 11804 18752
rect 11860 18718 11894 18752
rect 11950 18718 11984 18752
rect 12040 18718 12074 18752
rect 12130 18718 12164 18752
rect 12220 18718 12254 18752
rect 12310 18718 12344 18752
rect 12400 18718 12434 18752
rect 11309 18634 11343 18668
rect 12496 18634 12530 18668
rect 11309 18544 11343 18578
rect 11309 18454 11343 18488
rect 11309 18364 11343 18398
rect 11309 18274 11343 18308
rect 11309 18184 11343 18218
rect 11309 18094 11343 18128
rect 11309 18004 11343 18038
rect 11309 17914 11343 17948
rect 11309 17824 11343 17858
rect 11309 17734 11343 17768
rect 11309 17644 11343 17678
rect 12496 18544 12530 18578
rect 12496 18454 12530 18488
rect 12496 18364 12530 18398
rect 12496 18274 12530 18308
rect 12496 18184 12530 18218
rect 12496 18094 12530 18128
rect 12496 18004 12530 18038
rect 12496 17914 12530 17948
rect 12496 17824 12530 17858
rect 12496 17734 12530 17768
rect 12496 17644 12530 17678
rect 11309 17554 11343 17588
rect 11410 17531 11444 17565
rect 11500 17531 11534 17565
rect 11590 17531 11624 17565
rect 11680 17531 11714 17565
rect 11770 17531 11804 17565
rect 11860 17531 11894 17565
rect 11950 17531 11984 17565
rect 12040 17531 12074 17565
rect 12130 17531 12164 17565
rect 12220 17531 12254 17565
rect 12310 17531 12344 17565
rect 12400 17531 12434 17565
rect 12496 17554 12530 17588
rect 12770 18718 12804 18752
rect 12860 18718 12894 18752
rect 12950 18718 12984 18752
rect 13040 18718 13074 18752
rect 13130 18718 13164 18752
rect 13220 18718 13254 18752
rect 13310 18718 13344 18752
rect 13400 18718 13434 18752
rect 13490 18718 13524 18752
rect 13580 18718 13614 18752
rect 13670 18718 13704 18752
rect 13760 18718 13794 18752
rect 12669 18634 12703 18668
rect 13856 18634 13890 18668
rect 12669 18544 12703 18578
rect 12669 18454 12703 18488
rect 12669 18364 12703 18398
rect 12669 18274 12703 18308
rect 12669 18184 12703 18218
rect 12669 18094 12703 18128
rect 12669 18004 12703 18038
rect 12669 17914 12703 17948
rect 12669 17824 12703 17858
rect 12669 17734 12703 17768
rect 12669 17644 12703 17678
rect 13856 18544 13890 18578
rect 13856 18454 13890 18488
rect 13856 18364 13890 18398
rect 13856 18274 13890 18308
rect 13856 18184 13890 18218
rect 13856 18094 13890 18128
rect 13856 18004 13890 18038
rect 13856 17914 13890 17948
rect 13856 17824 13890 17858
rect 13856 17734 13890 17768
rect 13856 17644 13890 17678
rect 12669 17554 12703 17588
rect 12770 17531 12804 17565
rect 12860 17531 12894 17565
rect 12950 17531 12984 17565
rect 13040 17531 13074 17565
rect 13130 17531 13164 17565
rect 13220 17531 13254 17565
rect 13310 17531 13344 17565
rect 13400 17531 13434 17565
rect 13490 17531 13524 17565
rect 13580 17531 13614 17565
rect 13670 17531 13704 17565
rect 13760 17531 13794 17565
rect 13856 17554 13890 17588
rect 14130 18718 14164 18752
rect 14220 18718 14254 18752
rect 14310 18718 14344 18752
rect 14400 18718 14434 18752
rect 14490 18718 14524 18752
rect 14580 18718 14614 18752
rect 14670 18718 14704 18752
rect 14760 18718 14794 18752
rect 14850 18718 14884 18752
rect 14940 18718 14974 18752
rect 15030 18718 15064 18752
rect 15120 18718 15154 18752
rect 14029 18634 14063 18668
rect 15216 18634 15250 18668
rect 14029 18544 14063 18578
rect 14029 18454 14063 18488
rect 14029 18364 14063 18398
rect 14029 18274 14063 18308
rect 14029 18184 14063 18218
rect 14029 18094 14063 18128
rect 14029 18004 14063 18038
rect 14029 17914 14063 17948
rect 14029 17824 14063 17858
rect 14029 17734 14063 17768
rect 14029 17644 14063 17678
rect 15216 18544 15250 18578
rect 15216 18454 15250 18488
rect 15216 18364 15250 18398
rect 15216 18274 15250 18308
rect 15216 18184 15250 18218
rect 15216 18094 15250 18128
rect 15216 18004 15250 18038
rect 15216 17914 15250 17948
rect 15216 17824 15250 17858
rect 15216 17734 15250 17768
rect 15216 17644 15250 17678
rect 14029 17554 14063 17588
rect 14130 17531 14164 17565
rect 14220 17531 14254 17565
rect 14310 17531 14344 17565
rect 14400 17531 14434 17565
rect 14490 17531 14524 17565
rect 14580 17531 14614 17565
rect 14670 17531 14704 17565
rect 14760 17531 14794 17565
rect 14850 17531 14884 17565
rect 14940 17531 14974 17565
rect 15030 17531 15064 17565
rect 15120 17531 15154 17565
rect 15216 17554 15250 17588
rect 11410 17358 11444 17392
rect 11500 17358 11534 17392
rect 11590 17358 11624 17392
rect 11680 17358 11714 17392
rect 11770 17358 11804 17392
rect 11860 17358 11894 17392
rect 11950 17358 11984 17392
rect 12040 17358 12074 17392
rect 12130 17358 12164 17392
rect 12220 17358 12254 17392
rect 12310 17358 12344 17392
rect 12400 17358 12434 17392
rect 11309 17274 11343 17308
rect 12496 17274 12530 17308
rect 11309 17184 11343 17218
rect 11309 17094 11343 17128
rect 11309 17004 11343 17038
rect 11309 16914 11343 16948
rect 11309 16824 11343 16858
rect 11309 16734 11343 16768
rect 11309 16644 11343 16678
rect 11309 16554 11343 16588
rect 11309 16464 11343 16498
rect 11309 16374 11343 16408
rect 11309 16284 11343 16318
rect 12496 17184 12530 17218
rect 12496 17094 12530 17128
rect 12496 17004 12530 17038
rect 12496 16914 12530 16948
rect 12496 16824 12530 16858
rect 12496 16734 12530 16768
rect 12496 16644 12530 16678
rect 12496 16554 12530 16588
rect 12496 16464 12530 16498
rect 12496 16374 12530 16408
rect 12496 16284 12530 16318
rect 11309 16194 11343 16228
rect 11410 16171 11444 16205
rect 11500 16171 11534 16205
rect 11590 16171 11624 16205
rect 11680 16171 11714 16205
rect 11770 16171 11804 16205
rect 11860 16171 11894 16205
rect 11950 16171 11984 16205
rect 12040 16171 12074 16205
rect 12130 16171 12164 16205
rect 12220 16171 12254 16205
rect 12310 16171 12344 16205
rect 12400 16171 12434 16205
rect 12496 16194 12530 16228
rect 12770 17358 12804 17392
rect 12860 17358 12894 17392
rect 12950 17358 12984 17392
rect 13040 17358 13074 17392
rect 13130 17358 13164 17392
rect 13220 17358 13254 17392
rect 13310 17358 13344 17392
rect 13400 17358 13434 17392
rect 13490 17358 13524 17392
rect 13580 17358 13614 17392
rect 13670 17358 13704 17392
rect 13760 17358 13794 17392
rect 12669 17274 12703 17308
rect 13856 17274 13890 17308
rect 12669 17184 12703 17218
rect 12669 17094 12703 17128
rect 12669 17004 12703 17038
rect 12669 16914 12703 16948
rect 12669 16824 12703 16858
rect 12669 16734 12703 16768
rect 12669 16644 12703 16678
rect 12669 16554 12703 16588
rect 12669 16464 12703 16498
rect 12669 16374 12703 16408
rect 12669 16284 12703 16318
rect 13856 17184 13890 17218
rect 13856 17094 13890 17128
rect 13856 17004 13890 17038
rect 13856 16914 13890 16948
rect 13856 16824 13890 16858
rect 13856 16734 13890 16768
rect 13856 16644 13890 16678
rect 13856 16554 13890 16588
rect 13856 16464 13890 16498
rect 13856 16374 13890 16408
rect 13856 16284 13890 16318
rect 12669 16194 12703 16228
rect 12770 16171 12804 16205
rect 12860 16171 12894 16205
rect 12950 16171 12984 16205
rect 13040 16171 13074 16205
rect 13130 16171 13164 16205
rect 13220 16171 13254 16205
rect 13310 16171 13344 16205
rect 13400 16171 13434 16205
rect 13490 16171 13524 16205
rect 13580 16171 13614 16205
rect 13670 16171 13704 16205
rect 13760 16171 13794 16205
rect 13856 16194 13890 16228
rect 14130 17358 14164 17392
rect 14220 17358 14254 17392
rect 14310 17358 14344 17392
rect 14400 17358 14434 17392
rect 14490 17358 14524 17392
rect 14580 17358 14614 17392
rect 14670 17358 14704 17392
rect 14760 17358 14794 17392
rect 14850 17358 14884 17392
rect 14940 17358 14974 17392
rect 15030 17358 15064 17392
rect 15120 17358 15154 17392
rect 14029 17274 14063 17308
rect 15216 17274 15250 17308
rect 14029 17184 14063 17218
rect 14029 17094 14063 17128
rect 14029 17004 14063 17038
rect 14029 16914 14063 16948
rect 14029 16824 14063 16858
rect 14029 16734 14063 16768
rect 14029 16644 14063 16678
rect 14029 16554 14063 16588
rect 14029 16464 14063 16498
rect 14029 16374 14063 16408
rect 14029 16284 14063 16318
rect 15216 17184 15250 17218
rect 15216 17094 15250 17128
rect 15216 17004 15250 17038
rect 15216 16914 15250 16948
rect 15216 16824 15250 16858
rect 15216 16734 15250 16768
rect 15216 16644 15250 16678
rect 15216 16554 15250 16588
rect 15216 16464 15250 16498
rect 15216 16374 15250 16408
rect 15216 16284 15250 16318
rect 14029 16194 14063 16228
rect 14130 16171 14164 16205
rect 14220 16171 14254 16205
rect 14310 16171 14344 16205
rect 14400 16171 14434 16205
rect 14490 16171 14524 16205
rect 14580 16171 14614 16205
rect 14670 16171 14704 16205
rect 14760 16171 14794 16205
rect 14850 16171 14884 16205
rect 14940 16171 14974 16205
rect 15030 16171 15064 16205
rect 15120 16171 15154 16205
rect 15216 16194 15250 16228
rect 11410 15998 11444 16032
rect 11500 15998 11534 16032
rect 11590 15998 11624 16032
rect 11680 15998 11714 16032
rect 11770 15998 11804 16032
rect 11860 15998 11894 16032
rect 11950 15998 11984 16032
rect 12040 15998 12074 16032
rect 12130 15998 12164 16032
rect 12220 15998 12254 16032
rect 12310 15998 12344 16032
rect 12400 15998 12434 16032
rect 11309 15914 11343 15948
rect 12496 15914 12530 15948
rect 11309 15824 11343 15858
rect 11309 15734 11343 15768
rect 11309 15644 11343 15678
rect 11309 15554 11343 15588
rect 11309 15464 11343 15498
rect 11309 15374 11343 15408
rect 11309 15284 11343 15318
rect 11309 15194 11343 15228
rect 11309 15104 11343 15138
rect 11309 15014 11343 15048
rect 11309 14924 11343 14958
rect 12496 15824 12530 15858
rect 12496 15734 12530 15768
rect 12496 15644 12530 15678
rect 12496 15554 12530 15588
rect 12496 15464 12530 15498
rect 12496 15374 12530 15408
rect 12496 15284 12530 15318
rect 12496 15194 12530 15228
rect 12496 15104 12530 15138
rect 12496 15014 12530 15048
rect 12496 14924 12530 14958
rect 11309 14834 11343 14868
rect 11410 14811 11444 14845
rect 11500 14811 11534 14845
rect 11590 14811 11624 14845
rect 11680 14811 11714 14845
rect 11770 14811 11804 14845
rect 11860 14811 11894 14845
rect 11950 14811 11984 14845
rect 12040 14811 12074 14845
rect 12130 14811 12164 14845
rect 12220 14811 12254 14845
rect 12310 14811 12344 14845
rect 12400 14811 12434 14845
rect 12496 14834 12530 14868
rect 12770 15998 12804 16032
rect 12860 15998 12894 16032
rect 12950 15998 12984 16032
rect 13040 15998 13074 16032
rect 13130 15998 13164 16032
rect 13220 15998 13254 16032
rect 13310 15998 13344 16032
rect 13400 15998 13434 16032
rect 13490 15998 13524 16032
rect 13580 15998 13614 16032
rect 13670 15998 13704 16032
rect 13760 15998 13794 16032
rect 12669 15914 12703 15948
rect 13856 15914 13890 15948
rect 12669 15824 12703 15858
rect 12669 15734 12703 15768
rect 12669 15644 12703 15678
rect 12669 15554 12703 15588
rect 12669 15464 12703 15498
rect 12669 15374 12703 15408
rect 12669 15284 12703 15318
rect 12669 15194 12703 15228
rect 12669 15104 12703 15138
rect 12669 15014 12703 15048
rect 12669 14924 12703 14958
rect 13856 15824 13890 15858
rect 13856 15734 13890 15768
rect 13856 15644 13890 15678
rect 13856 15554 13890 15588
rect 13856 15464 13890 15498
rect 13856 15374 13890 15408
rect 13856 15284 13890 15318
rect 13856 15194 13890 15228
rect 13856 15104 13890 15138
rect 13856 15014 13890 15048
rect 13856 14924 13890 14958
rect 12669 14834 12703 14868
rect 12770 14811 12804 14845
rect 12860 14811 12894 14845
rect 12950 14811 12984 14845
rect 13040 14811 13074 14845
rect 13130 14811 13164 14845
rect 13220 14811 13254 14845
rect 13310 14811 13344 14845
rect 13400 14811 13434 14845
rect 13490 14811 13524 14845
rect 13580 14811 13614 14845
rect 13670 14811 13704 14845
rect 13760 14811 13794 14845
rect 13856 14834 13890 14868
rect 14130 15998 14164 16032
rect 14220 15998 14254 16032
rect 14310 15998 14344 16032
rect 14400 15998 14434 16032
rect 14490 15998 14524 16032
rect 14580 15998 14614 16032
rect 14670 15998 14704 16032
rect 14760 15998 14794 16032
rect 14850 15998 14884 16032
rect 14940 15998 14974 16032
rect 15030 15998 15064 16032
rect 15120 15998 15154 16032
rect 14029 15914 14063 15948
rect 15216 15914 15250 15948
rect 14029 15824 14063 15858
rect 14029 15734 14063 15768
rect 14029 15644 14063 15678
rect 14029 15554 14063 15588
rect 14029 15464 14063 15498
rect 14029 15374 14063 15408
rect 14029 15284 14063 15318
rect 14029 15194 14063 15228
rect 14029 15104 14063 15138
rect 14029 15014 14063 15048
rect 14029 14924 14063 14958
rect 15216 15824 15250 15858
rect 15216 15734 15250 15768
rect 15216 15644 15250 15678
rect 15216 15554 15250 15588
rect 15216 15464 15250 15498
rect 15216 15374 15250 15408
rect 15216 15284 15250 15318
rect 15216 15194 15250 15228
rect 15216 15104 15250 15138
rect 15216 15014 15250 15048
rect 15216 14924 15250 14958
rect 14029 14834 14063 14868
rect 14130 14811 14164 14845
rect 14220 14811 14254 14845
rect 14310 14811 14344 14845
rect 14400 14811 14434 14845
rect 14490 14811 14524 14845
rect 14580 14811 14614 14845
rect 14670 14811 14704 14845
rect 14760 14811 14794 14845
rect 14850 14811 14884 14845
rect 14940 14811 14974 14845
rect 15030 14811 15064 14845
rect 15120 14811 15154 14845
rect 15216 14834 15250 14868
rect 15420 14210 15460 14250
rect 15420 14110 15460 14150
rect 11920 13600 11960 13640
rect 11920 13500 11960 13540
rect 11920 13400 11960 13440
rect 11920 13300 11960 13340
rect 11920 13200 11960 13240
rect 14600 13600 14640 13640
rect 14600 13500 14640 13540
rect 14600 13400 14640 13440
rect 14600 13300 14640 13340
rect 14600 13200 14640 13240
rect 12820 12680 12860 12720
rect 12820 12600 12860 12640
rect 12820 12520 12860 12560
rect 13700 12680 13740 12720
rect 13700 12600 13740 12640
rect 13700 12520 13740 12560
<< nsubdiffcont >>
rect 8359 18563 8619 18597
rect 8263 17173 8297 18501
rect 8681 17173 8715 18501
rect 8359 17077 8619 17111
rect 9146 18566 9738 18600
rect 9050 16774 9084 18504
rect 9800 16774 9834 18504
rect 9146 16678 9738 16712
rect 10259 18563 10851 18597
rect 10163 16243 10197 18501
rect 10913 16243 10947 18501
rect 11550 18568 11584 18602
rect 11640 18568 11674 18602
rect 11730 18568 11764 18602
rect 11820 18568 11854 18602
rect 11910 18568 11944 18602
rect 12000 18568 12034 18602
rect 12090 18568 12124 18602
rect 12180 18568 12214 18602
rect 12270 18568 12304 18602
rect 11458 18474 11492 18508
rect 11458 18384 11492 18418
rect 11458 18294 11492 18328
rect 11458 18204 11492 18238
rect 11458 18114 11492 18148
rect 11458 18024 11492 18058
rect 11458 17934 11492 17968
rect 11458 17844 11492 17878
rect 12348 18455 12382 18489
rect 12348 18365 12382 18399
rect 12348 18275 12382 18309
rect 12348 18185 12382 18219
rect 12348 18095 12382 18129
rect 12348 18005 12382 18039
rect 12348 17915 12382 17949
rect 12348 17825 12382 17859
rect 11458 17754 11492 17788
rect 12348 17735 12382 17769
rect 11516 17678 11550 17712
rect 11606 17678 11640 17712
rect 11696 17678 11730 17712
rect 11786 17678 11820 17712
rect 11876 17678 11910 17712
rect 11966 17678 12000 17712
rect 12056 17678 12090 17712
rect 12146 17678 12180 17712
rect 12236 17678 12270 17712
rect 12910 18568 12944 18602
rect 13000 18568 13034 18602
rect 13090 18568 13124 18602
rect 13180 18568 13214 18602
rect 13270 18568 13304 18602
rect 13360 18568 13394 18602
rect 13450 18568 13484 18602
rect 13540 18568 13574 18602
rect 13630 18568 13664 18602
rect 12818 18474 12852 18508
rect 12818 18384 12852 18418
rect 12818 18294 12852 18328
rect 12818 18204 12852 18238
rect 12818 18114 12852 18148
rect 12818 18024 12852 18058
rect 12818 17934 12852 17968
rect 12818 17844 12852 17878
rect 13708 18455 13742 18489
rect 13708 18365 13742 18399
rect 13708 18275 13742 18309
rect 13708 18185 13742 18219
rect 13708 18095 13742 18129
rect 13708 18005 13742 18039
rect 13708 17915 13742 17949
rect 13708 17825 13742 17859
rect 12818 17754 12852 17788
rect 13708 17735 13742 17769
rect 12876 17678 12910 17712
rect 12966 17678 13000 17712
rect 13056 17678 13090 17712
rect 13146 17678 13180 17712
rect 13236 17678 13270 17712
rect 13326 17678 13360 17712
rect 13416 17678 13450 17712
rect 13506 17678 13540 17712
rect 13596 17678 13630 17712
rect 14270 18568 14304 18602
rect 14360 18568 14394 18602
rect 14450 18568 14484 18602
rect 14540 18568 14574 18602
rect 14630 18568 14664 18602
rect 14720 18568 14754 18602
rect 14810 18568 14844 18602
rect 14900 18568 14934 18602
rect 14990 18568 15024 18602
rect 14178 18474 14212 18508
rect 14178 18384 14212 18418
rect 14178 18294 14212 18328
rect 14178 18204 14212 18238
rect 14178 18114 14212 18148
rect 14178 18024 14212 18058
rect 14178 17934 14212 17968
rect 14178 17844 14212 17878
rect 15068 18455 15102 18489
rect 15068 18365 15102 18399
rect 15068 18275 15102 18309
rect 15068 18185 15102 18219
rect 15068 18095 15102 18129
rect 15068 18005 15102 18039
rect 15068 17915 15102 17949
rect 15068 17825 15102 17859
rect 14178 17754 14212 17788
rect 15068 17735 15102 17769
rect 14236 17678 14270 17712
rect 14326 17678 14360 17712
rect 14416 17678 14450 17712
rect 14506 17678 14540 17712
rect 14596 17678 14630 17712
rect 14686 17678 14720 17712
rect 14776 17678 14810 17712
rect 14866 17678 14900 17712
rect 14956 17678 14990 17712
rect 15579 18563 16171 18597
rect 10259 16147 10851 16181
rect 11550 17208 11584 17242
rect 11640 17208 11674 17242
rect 11730 17208 11764 17242
rect 11820 17208 11854 17242
rect 11910 17208 11944 17242
rect 12000 17208 12034 17242
rect 12090 17208 12124 17242
rect 12180 17208 12214 17242
rect 12270 17208 12304 17242
rect 11458 17114 11492 17148
rect 11458 17024 11492 17058
rect 11458 16934 11492 16968
rect 11458 16844 11492 16878
rect 11458 16754 11492 16788
rect 11458 16664 11492 16698
rect 11458 16574 11492 16608
rect 11458 16484 11492 16518
rect 12348 17095 12382 17129
rect 12348 17005 12382 17039
rect 12348 16915 12382 16949
rect 12348 16825 12382 16859
rect 12348 16735 12382 16769
rect 12348 16645 12382 16679
rect 12348 16555 12382 16589
rect 12348 16465 12382 16499
rect 11458 16394 11492 16428
rect 12348 16375 12382 16409
rect 11516 16318 11550 16352
rect 11606 16318 11640 16352
rect 11696 16318 11730 16352
rect 11786 16318 11820 16352
rect 11876 16318 11910 16352
rect 11966 16318 12000 16352
rect 12056 16318 12090 16352
rect 12146 16318 12180 16352
rect 12236 16318 12270 16352
rect 12910 17208 12944 17242
rect 13000 17208 13034 17242
rect 13090 17208 13124 17242
rect 13180 17208 13214 17242
rect 13270 17208 13304 17242
rect 13360 17208 13394 17242
rect 13450 17208 13484 17242
rect 13540 17208 13574 17242
rect 13630 17208 13664 17242
rect 12818 17114 12852 17148
rect 12818 17024 12852 17058
rect 12818 16934 12852 16968
rect 12818 16844 12852 16878
rect 12818 16754 12852 16788
rect 12818 16664 12852 16698
rect 12818 16574 12852 16608
rect 12818 16484 12852 16518
rect 13708 17095 13742 17129
rect 13708 17005 13742 17039
rect 13708 16915 13742 16949
rect 13708 16825 13742 16859
rect 13708 16735 13742 16769
rect 13708 16645 13742 16679
rect 13708 16555 13742 16589
rect 13708 16465 13742 16499
rect 12818 16394 12852 16428
rect 13708 16375 13742 16409
rect 12876 16318 12910 16352
rect 12966 16318 13000 16352
rect 13056 16318 13090 16352
rect 13146 16318 13180 16352
rect 13236 16318 13270 16352
rect 13326 16318 13360 16352
rect 13416 16318 13450 16352
rect 13506 16318 13540 16352
rect 13596 16318 13630 16352
rect 14270 17208 14304 17242
rect 14360 17208 14394 17242
rect 14450 17208 14484 17242
rect 14540 17208 14574 17242
rect 14630 17208 14664 17242
rect 14720 17208 14754 17242
rect 14810 17208 14844 17242
rect 14900 17208 14934 17242
rect 14990 17208 15024 17242
rect 14178 17114 14212 17148
rect 14178 17024 14212 17058
rect 14178 16934 14212 16968
rect 14178 16844 14212 16878
rect 14178 16754 14212 16788
rect 14178 16664 14212 16698
rect 14178 16574 14212 16608
rect 14178 16484 14212 16518
rect 15068 17095 15102 17129
rect 15068 17005 15102 17039
rect 15068 16915 15102 16949
rect 15068 16825 15102 16859
rect 15068 16735 15102 16769
rect 15068 16645 15102 16679
rect 15068 16555 15102 16589
rect 15068 16465 15102 16499
rect 14178 16394 14212 16428
rect 15068 16375 15102 16409
rect 14236 16318 14270 16352
rect 14326 16318 14360 16352
rect 14416 16318 14450 16352
rect 14506 16318 14540 16352
rect 14596 16318 14630 16352
rect 14686 16318 14720 16352
rect 14776 16318 14810 16352
rect 14866 16318 14900 16352
rect 14956 16318 14990 16352
rect 15483 16243 15517 18501
rect 16233 16243 16267 18501
rect 16692 18560 16952 18594
rect 16596 17380 16630 18498
rect 17014 17380 17048 18498
rect 16692 17284 16952 17318
rect 17479 18563 17739 18597
rect 17383 17173 17417 18501
rect 17801 17173 17835 18501
rect 17479 17077 17739 17111
rect 15579 16147 16171 16181
rect 11550 15848 11584 15882
rect 11640 15848 11674 15882
rect 11730 15848 11764 15882
rect 11820 15848 11854 15882
rect 11910 15848 11944 15882
rect 12000 15848 12034 15882
rect 12090 15848 12124 15882
rect 12180 15848 12214 15882
rect 12270 15848 12304 15882
rect 11458 15754 11492 15788
rect 11458 15664 11492 15698
rect 11458 15574 11492 15608
rect 11458 15484 11492 15518
rect 11458 15394 11492 15428
rect 11458 15304 11492 15338
rect 11458 15214 11492 15248
rect 11458 15124 11492 15158
rect 12348 15735 12382 15769
rect 12348 15645 12382 15679
rect 12348 15555 12382 15589
rect 12348 15465 12382 15499
rect 12348 15375 12382 15409
rect 12348 15285 12382 15319
rect 12348 15195 12382 15229
rect 12348 15105 12382 15139
rect 11458 15034 11492 15068
rect 12348 15015 12382 15049
rect 11516 14958 11550 14992
rect 11606 14958 11640 14992
rect 11696 14958 11730 14992
rect 11786 14958 11820 14992
rect 11876 14958 11910 14992
rect 11966 14958 12000 14992
rect 12056 14958 12090 14992
rect 12146 14958 12180 14992
rect 12236 14958 12270 14992
rect 12910 15848 12944 15882
rect 13000 15848 13034 15882
rect 13090 15848 13124 15882
rect 13180 15848 13214 15882
rect 13270 15848 13304 15882
rect 13360 15848 13394 15882
rect 13450 15848 13484 15882
rect 13540 15848 13574 15882
rect 13630 15848 13664 15882
rect 12818 15754 12852 15788
rect 12818 15664 12852 15698
rect 12818 15574 12852 15608
rect 12818 15484 12852 15518
rect 12818 15394 12852 15428
rect 12818 15304 12852 15338
rect 12818 15214 12852 15248
rect 12818 15124 12852 15158
rect 13708 15735 13742 15769
rect 13708 15645 13742 15679
rect 13708 15555 13742 15589
rect 13708 15465 13742 15499
rect 13708 15375 13742 15409
rect 13708 15285 13742 15319
rect 13708 15195 13742 15229
rect 13708 15105 13742 15139
rect 12818 15034 12852 15068
rect 13708 15015 13742 15049
rect 12876 14958 12910 14992
rect 12966 14958 13000 14992
rect 13056 14958 13090 14992
rect 13146 14958 13180 14992
rect 13236 14958 13270 14992
rect 13326 14958 13360 14992
rect 13416 14958 13450 14992
rect 13506 14958 13540 14992
rect 13596 14958 13630 14992
rect 14270 15848 14304 15882
rect 14360 15848 14394 15882
rect 14450 15848 14484 15882
rect 14540 15848 14574 15882
rect 14630 15848 14664 15882
rect 14720 15848 14754 15882
rect 14810 15848 14844 15882
rect 14900 15848 14934 15882
rect 14990 15848 15024 15882
rect 14178 15754 14212 15788
rect 14178 15664 14212 15698
rect 14178 15574 14212 15608
rect 14178 15484 14212 15518
rect 14178 15394 14212 15428
rect 14178 15304 14212 15338
rect 14178 15214 14212 15248
rect 14178 15124 14212 15158
rect 15068 15735 15102 15769
rect 15068 15645 15102 15679
rect 15068 15555 15102 15589
rect 15068 15465 15102 15499
rect 15068 15375 15102 15409
rect 15068 15285 15102 15319
rect 15068 15195 15102 15229
rect 15068 15105 15102 15139
rect 14178 15034 14212 15068
rect 15068 15015 15102 15049
rect 14236 14958 14270 14992
rect 14326 14958 14360 14992
rect 14416 14958 14450 14992
rect 14506 14958 14540 14992
rect 14596 14958 14630 14992
rect 14686 14958 14720 14992
rect 14776 14958 14810 14992
rect 14866 14958 14900 14992
rect 14956 14958 14990 14992
rect 10460 11750 10500 11790
rect 10460 11650 10500 11690
rect 13020 11750 13060 11790
rect 13020 11650 13060 11690
rect 13500 11750 13540 11790
rect 13500 11650 13540 11690
rect 16060 11750 16100 11790
rect 16060 11650 16100 11690
rect 11560 10590 11600 10630
rect 11560 10490 11600 10530
rect 11560 10390 11600 10430
rect 11560 10290 11600 10330
rect 11560 10190 11600 10230
rect 11560 10090 11600 10130
rect 14960 10590 15000 10630
rect 14960 10490 15000 10530
rect 14960 10390 15000 10430
rect 14960 10290 15000 10330
rect 15420 10390 15460 10430
rect 15420 10290 15460 10330
rect 16030 10390 16070 10430
rect 16030 10290 16070 10330
rect 14960 10190 15000 10230
rect 14960 10090 15000 10130
rect 11570 9590 11610 9630
rect 11570 9490 11610 9530
rect 13050 9590 13090 9630
rect 13050 9490 13090 9530
rect 13470 9590 13510 9630
rect 13470 9490 13510 9530
rect 14950 9590 14990 9630
rect 14950 9490 14990 9530
<< poly >>
rect 11240 14280 13240 14310
rect 13320 14280 15320 14310
rect 11240 14050 13240 14080
rect 13320 14050 15320 14080
rect 11320 14030 11400 14050
rect 11320 13990 11340 14030
rect 11380 13990 11400 14030
rect 11320 13970 11400 13990
rect 11480 14030 11560 14050
rect 11480 13990 11500 14030
rect 11540 13990 11560 14030
rect 11480 13970 11560 13990
rect 11640 14030 11720 14050
rect 11640 13990 11660 14030
rect 11700 13990 11720 14030
rect 11640 13970 11720 13990
rect 11800 14030 11880 14050
rect 11800 13990 11820 14030
rect 11860 13990 11880 14030
rect 11800 13970 11880 13990
rect 11960 14030 12040 14050
rect 11960 13990 11980 14030
rect 12020 13990 12040 14030
rect 11960 13970 12040 13990
rect 12120 14030 12200 14050
rect 12120 13990 12140 14030
rect 12180 13990 12200 14030
rect 12120 13970 12200 13990
rect 12280 14030 12360 14050
rect 12280 13990 12300 14030
rect 12340 13990 12360 14030
rect 12280 13970 12360 13990
rect 12440 14030 12520 14050
rect 12440 13990 12460 14030
rect 12500 13990 12520 14030
rect 12440 13970 12520 13990
rect 12600 14030 12680 14050
rect 12600 13990 12620 14030
rect 12660 13990 12680 14030
rect 12600 13970 12680 13990
rect 12760 14030 12840 14050
rect 12760 13990 12780 14030
rect 12820 13990 12840 14030
rect 12760 13970 12840 13990
rect 12920 14030 13000 14050
rect 12920 13990 12940 14030
rect 12980 13990 13000 14030
rect 12920 13970 13000 13990
rect 13080 14030 13160 14050
rect 13080 13990 13100 14030
rect 13140 13990 13160 14030
rect 13080 13970 13160 13990
rect 13400 14030 13480 14050
rect 13400 13990 13420 14030
rect 13460 13990 13480 14030
rect 13400 13970 13480 13990
rect 13560 14030 13640 14050
rect 13560 13990 13580 14030
rect 13620 13990 13640 14030
rect 13560 13970 13640 13990
rect 13720 14030 13800 14050
rect 13720 13990 13740 14030
rect 13780 13990 13800 14030
rect 13720 13970 13800 13990
rect 13880 14030 13960 14050
rect 13880 13990 13900 14030
rect 13940 13990 13960 14030
rect 13880 13970 13960 13990
rect 14040 14030 14120 14050
rect 14040 13990 14060 14030
rect 14100 13990 14120 14030
rect 14040 13970 14120 13990
rect 14200 14030 14280 14050
rect 14200 13990 14220 14030
rect 14260 13990 14280 14030
rect 14200 13970 14280 13990
rect 14360 14030 14440 14050
rect 14360 13990 14380 14030
rect 14420 13990 14440 14030
rect 14360 13970 14440 13990
rect 14520 14030 14600 14050
rect 14520 13990 14540 14030
rect 14580 13990 14600 14030
rect 14520 13970 14600 13990
rect 14680 14030 14760 14050
rect 14680 13990 14700 14030
rect 14740 13990 14760 14030
rect 14680 13970 14760 13990
rect 14840 14030 14920 14050
rect 14840 13990 14860 14030
rect 14900 13990 14920 14030
rect 14840 13970 14920 13990
rect 15000 14030 15080 14050
rect 15000 13990 15020 14030
rect 15060 13990 15080 14030
rect 15000 13970 15080 13990
rect 15160 14030 15240 14050
rect 15160 13990 15180 14030
rect 15220 13990 15240 14030
rect 15160 13970 15240 13990
rect 10820 13670 11820 13700
rect 12060 13670 13060 13700
rect 13500 13670 14500 13700
rect 14740 13670 15740 13700
rect 10820 13140 11820 13170
rect 12060 13140 13060 13170
rect 13500 13140 14500 13170
rect 14740 13140 15740 13170
rect 10920 13120 11000 13140
rect 10920 13080 10940 13120
rect 10980 13080 11000 13120
rect 10920 13060 11000 13080
rect 11160 13120 11240 13140
rect 11160 13080 11180 13120
rect 11220 13080 11240 13120
rect 11160 13060 11240 13080
rect 11400 13120 11480 13140
rect 11400 13080 11420 13120
rect 11460 13080 11480 13120
rect 11400 13060 11480 13080
rect 11640 13120 11720 13140
rect 11640 13080 11660 13120
rect 11700 13080 11720 13120
rect 11640 13060 11720 13080
rect 12280 13120 12360 13140
rect 12280 13080 12300 13120
rect 12340 13080 12360 13120
rect 12280 13060 12360 13080
rect 12520 13120 12600 13140
rect 12520 13080 12540 13120
rect 12580 13080 12600 13120
rect 12520 13060 12600 13080
rect 12760 13120 12840 13140
rect 12760 13080 12780 13120
rect 12820 13080 12840 13120
rect 12760 13060 12840 13080
rect 13720 13120 13800 13140
rect 13720 13080 13740 13120
rect 13780 13080 13800 13120
rect 13720 13060 13800 13080
rect 13960 13120 14040 13140
rect 13960 13080 13980 13120
rect 14020 13080 14040 13120
rect 13960 13060 14040 13080
rect 14200 13120 14280 13140
rect 14200 13080 14220 13120
rect 14260 13080 14280 13120
rect 14200 13060 14280 13080
rect 14840 13120 14920 13140
rect 14840 13080 14860 13120
rect 14900 13080 14920 13120
rect 14840 13060 14920 13080
rect 15080 13120 15160 13140
rect 15080 13080 15100 13120
rect 15140 13080 15160 13120
rect 15080 13060 15160 13080
rect 15320 13120 15400 13140
rect 15320 13080 15340 13120
rect 15380 13080 15400 13120
rect 15320 13060 15400 13080
rect 15560 13120 15640 13140
rect 15560 13080 15580 13120
rect 15620 13080 15640 13120
rect 15560 13060 15640 13080
rect 11431 12742 11489 12760
rect 11431 12708 11443 12742
rect 11477 12708 11489 12742
rect 11431 12690 11489 12708
rect 11791 12742 11849 12760
rect 11791 12708 11803 12742
rect 11837 12708 11849 12742
rect 11791 12690 11849 12708
rect 11911 12742 11969 12760
rect 11911 12708 11923 12742
rect 11957 12708 11969 12742
rect 11911 12690 11969 12708
rect 12271 12742 12329 12760
rect 12271 12708 12283 12742
rect 12317 12708 12329 12742
rect 12271 12690 12329 12708
rect 12391 12742 12449 12760
rect 12391 12708 12403 12742
rect 12437 12708 12449 12742
rect 12391 12690 12449 12708
rect 11440 12660 11480 12690
rect 11560 12660 11600 12690
rect 11680 12660 11720 12690
rect 11800 12660 11840 12690
rect 11920 12660 11960 12690
rect 12040 12660 12080 12690
rect 12160 12660 12200 12690
rect 12280 12660 12320 12690
rect 12400 12660 12440 12690
rect 12520 12660 12560 12690
rect 11440 12530 11480 12560
rect 11560 12530 11600 12560
rect 11532 12512 11600 12530
rect 11532 12478 11544 12512
rect 11578 12478 11600 12512
rect 11532 12460 11600 12478
rect 11680 12530 11720 12560
rect 11800 12530 11840 12560
rect 11920 12530 11960 12560
rect 12040 12530 12080 12560
rect 11680 12512 11748 12530
rect 11680 12478 11702 12512
rect 11736 12478 11748 12512
rect 11680 12460 11748 12478
rect 12014 12512 12080 12530
rect 12014 12478 12026 12512
rect 12060 12478 12080 12512
rect 12014 12460 12080 12478
rect 12160 12530 12200 12560
rect 12280 12530 12320 12560
rect 12400 12530 12440 12560
rect 12520 12530 12560 12560
rect 12160 12512 12226 12530
rect 12160 12478 12180 12512
rect 12214 12478 12226 12512
rect 12160 12460 12226 12478
rect 12492 12512 12560 12530
rect 12492 12478 12504 12512
rect 12538 12478 12560 12512
rect 14111 12742 14169 12760
rect 14111 12708 14123 12742
rect 14157 12708 14169 12742
rect 14111 12690 14169 12708
rect 14231 12742 14289 12760
rect 14231 12708 14243 12742
rect 14277 12708 14289 12742
rect 14231 12690 14289 12708
rect 14591 12742 14649 12760
rect 14591 12708 14603 12742
rect 14637 12708 14649 12742
rect 14591 12690 14649 12708
rect 14711 12742 14769 12760
rect 14711 12708 14723 12742
rect 14757 12708 14769 12742
rect 14711 12690 14769 12708
rect 15071 12742 15129 12760
rect 15071 12708 15083 12742
rect 15117 12708 15129 12742
rect 15071 12690 15129 12708
rect 14000 12660 14040 12690
rect 14120 12660 14160 12690
rect 14240 12660 14280 12690
rect 14360 12660 14400 12690
rect 14480 12660 14520 12690
rect 14600 12660 14640 12690
rect 14720 12660 14760 12690
rect 14840 12660 14880 12690
rect 14960 12660 15000 12690
rect 15080 12660 15120 12690
rect 14000 12530 14040 12560
rect 14120 12530 14160 12560
rect 14240 12530 14280 12560
rect 14360 12530 14400 12560
rect 14000 12512 14068 12530
rect 12492 12460 12560 12478
rect 14000 12478 14022 12512
rect 14056 12478 14068 12512
rect 14000 12460 14068 12478
rect 14334 12512 14400 12530
rect 14334 12478 14346 12512
rect 14380 12478 14400 12512
rect 14334 12460 14400 12478
rect 14480 12530 14520 12560
rect 14600 12530 14640 12560
rect 14720 12530 14760 12560
rect 14840 12530 14880 12560
rect 14480 12512 14546 12530
rect 14480 12478 14500 12512
rect 14534 12478 14546 12512
rect 14480 12460 14546 12478
rect 14812 12512 14880 12530
rect 14812 12478 14824 12512
rect 14858 12478 14880 12512
rect 14812 12460 14880 12478
rect 14960 12530 15000 12560
rect 15080 12530 15120 12560
rect 14960 12512 15028 12530
rect 14960 12478 14982 12512
rect 15016 12478 15028 12512
rect 14960 12460 15028 12478
rect 10710 11920 10770 11940
rect 10710 11880 10720 11920
rect 10760 11880 10770 11920
rect 10710 11860 10770 11880
rect 10880 11910 10960 11930
rect 10880 11870 10900 11910
rect 10940 11870 10960 11910
rect 11370 11910 11430 11930
rect 11370 11870 11380 11910
rect 11420 11870 11430 11910
rect 11600 11910 11680 11930
rect 11600 11870 11620 11910
rect 11660 11870 11680 11910
rect 12090 11910 12150 11930
rect 12090 11870 12100 11910
rect 12140 11870 12150 11910
rect 12320 11910 12400 11930
rect 12320 11870 12340 11910
rect 12380 11870 12400 11910
rect 12750 11910 12810 11930
rect 12750 11870 12760 11910
rect 12800 11870 12810 11910
rect 10600 11820 10640 11850
rect 10720 11820 10760 11860
rect 10840 11840 11240 11870
rect 10840 11820 10880 11840
rect 10960 11820 11000 11840
rect 11080 11820 11120 11840
rect 11200 11820 11240 11840
rect 11320 11840 11480 11870
rect 11320 11820 11360 11840
rect 11440 11820 11480 11840
rect 11560 11840 11960 11870
rect 11560 11820 11600 11840
rect 11680 11820 11720 11840
rect 11800 11820 11840 11840
rect 11920 11820 11960 11840
rect 12040 11840 12200 11870
rect 12040 11820 12080 11840
rect 12160 11820 12200 11840
rect 12280 11840 12680 11870
rect 12750 11850 12810 11870
rect 13750 11910 13810 11930
rect 13750 11870 13760 11910
rect 13800 11870 13810 11910
rect 14160 11910 14240 11930
rect 14160 11870 14180 11910
rect 14220 11870 14240 11910
rect 14410 11910 14470 11930
rect 14410 11870 14420 11910
rect 14460 11870 14470 11910
rect 14880 11910 14960 11930
rect 14880 11870 14900 11910
rect 14940 11870 14960 11910
rect 15130 11910 15190 11930
rect 15130 11870 15140 11910
rect 15180 11870 15190 11910
rect 15600 11910 15680 11930
rect 15600 11870 15620 11910
rect 15660 11870 15680 11910
rect 15790 11920 15850 11940
rect 15790 11880 15800 11920
rect 15840 11880 15850 11920
rect 13750 11850 13810 11870
rect 12280 11820 12320 11840
rect 12400 11820 12440 11840
rect 12520 11820 12560 11840
rect 12640 11820 12680 11840
rect 12760 11820 12800 11850
rect 12880 11820 12920 11850
rect 13640 11820 13680 11850
rect 13760 11820 13800 11850
rect 13880 11840 14280 11870
rect 13880 11820 13920 11840
rect 14000 11820 14040 11840
rect 14120 11820 14160 11840
rect 14240 11820 14280 11840
rect 14360 11840 14520 11870
rect 14360 11820 14400 11840
rect 14480 11820 14520 11840
rect 14600 11840 15000 11870
rect 14600 11820 14640 11840
rect 14720 11820 14760 11840
rect 14840 11820 14880 11840
rect 14960 11820 15000 11840
rect 15080 11840 15240 11870
rect 15080 11820 15120 11840
rect 15200 11820 15240 11840
rect 15320 11840 15720 11870
rect 15790 11860 15850 11880
rect 15320 11820 15360 11840
rect 15440 11820 15480 11840
rect 15560 11820 15600 11840
rect 15680 11820 15720 11840
rect 15800 11820 15840 11860
rect 15920 11820 15960 11850
rect 10600 11590 10640 11620
rect 10720 11590 10760 11620
rect 10840 11590 10880 11620
rect 10960 11590 11000 11620
rect 11080 11590 11120 11620
rect 11200 11590 11240 11620
rect 11320 11590 11360 11620
rect 11440 11590 11480 11620
rect 11560 11590 11600 11620
rect 11680 11590 11720 11620
rect 11800 11590 11840 11620
rect 11920 11590 11960 11620
rect 12040 11590 12080 11620
rect 12160 11590 12200 11620
rect 12280 11590 12320 11620
rect 12400 11590 12440 11620
rect 12520 11590 12560 11620
rect 12640 11590 12680 11620
rect 12760 11590 12800 11620
rect 12880 11590 12920 11620
rect 13640 11590 13680 11620
rect 13760 11590 13800 11620
rect 13880 11590 13920 11620
rect 14000 11590 14040 11620
rect 14120 11590 14160 11620
rect 14240 11590 14280 11620
rect 14360 11590 14400 11620
rect 14480 11590 14520 11620
rect 14600 11590 14640 11620
rect 14720 11590 14760 11620
rect 14840 11590 14880 11620
rect 14960 11590 15000 11620
rect 15080 11590 15120 11620
rect 15200 11590 15240 11620
rect 15320 11590 15360 11620
rect 15440 11590 15480 11620
rect 15560 11590 15600 11620
rect 15680 11590 15720 11620
rect 15800 11590 15840 11620
rect 15920 11590 15960 11620
rect 10530 11570 10640 11590
rect 10530 11530 10540 11570
rect 10580 11560 10640 11570
rect 12880 11570 12990 11590
rect 12880 11560 12940 11570
rect 10580 11530 10590 11560
rect 10530 11510 10590 11530
rect 12930 11530 12940 11560
rect 12980 11530 12990 11570
rect 12930 11510 12990 11530
rect 13570 11570 13680 11590
rect 13570 11530 13580 11570
rect 13620 11560 13680 11570
rect 15920 11570 16030 11590
rect 15920 11560 15980 11570
rect 13620 11530 13630 11560
rect 13570 11510 13630 11530
rect 15970 11530 15980 11560
rect 16020 11530 16030 11570
rect 15970 11510 16030 11530
rect 11900 10750 11970 10770
rect 11900 10710 11910 10750
rect 11950 10710 11970 10750
rect 11900 10690 11970 10710
rect 12070 10750 12150 10770
rect 12070 10710 12090 10750
rect 12130 10710 12150 10750
rect 12070 10690 12150 10710
rect 12250 10750 12330 10770
rect 12250 10710 12270 10750
rect 12310 10710 12330 10750
rect 12250 10690 12330 10710
rect 12430 10750 12510 10770
rect 12430 10710 12450 10750
rect 12490 10710 12510 10750
rect 12430 10690 12510 10710
rect 12610 10750 12690 10770
rect 12610 10710 12630 10750
rect 12670 10710 12690 10750
rect 12610 10690 12690 10710
rect 12790 10750 12870 10770
rect 12790 10710 12810 10750
rect 12850 10710 12870 10750
rect 12790 10690 12870 10710
rect 12970 10750 13050 10770
rect 12970 10710 12990 10750
rect 13030 10710 13050 10750
rect 12970 10690 13050 10710
rect 13150 10750 13220 10770
rect 13150 10710 13170 10750
rect 13210 10710 13220 10750
rect 13150 10690 13220 10710
rect 13340 10750 13410 10770
rect 13340 10710 13350 10750
rect 13390 10710 13410 10750
rect 13340 10690 13410 10710
rect 13510 10750 13590 10770
rect 13510 10710 13530 10750
rect 13570 10710 13590 10750
rect 13510 10690 13590 10710
rect 13690 10750 13770 10770
rect 13690 10710 13710 10750
rect 13750 10710 13770 10750
rect 13690 10690 13770 10710
rect 13870 10750 13950 10770
rect 13870 10710 13890 10750
rect 13930 10710 13950 10750
rect 13870 10690 13950 10710
rect 14050 10750 14130 10770
rect 14050 10710 14070 10750
rect 14110 10710 14130 10750
rect 14050 10690 14130 10710
rect 14230 10750 14310 10770
rect 14230 10710 14250 10750
rect 14290 10710 14310 10750
rect 14230 10690 14310 10710
rect 14410 10750 14490 10770
rect 14410 10710 14430 10750
rect 14470 10710 14490 10750
rect 14410 10690 14490 10710
rect 14590 10750 14660 10770
rect 14590 10710 14610 10750
rect 14650 10710 14660 10750
rect 14590 10700 14660 10710
rect 11700 10660 11800 10690
rect 11880 10660 11980 10690
rect 12060 10660 12160 10690
rect 12240 10660 12340 10690
rect 12420 10660 12520 10690
rect 12600 10660 12700 10690
rect 12780 10660 12880 10690
rect 12960 10660 13060 10690
rect 13140 10660 13240 10690
rect 13320 10660 13420 10690
rect 13500 10660 13600 10690
rect 13680 10660 13780 10690
rect 13860 10660 13960 10690
rect 14040 10660 14140 10690
rect 14220 10660 14320 10690
rect 14400 10660 14500 10690
rect 14580 10660 14680 10700
rect 14760 10660 14860 10690
rect 15710 10550 15790 10570
rect 15710 10510 15730 10550
rect 15770 10510 15790 10550
rect 15570 10460 15600 10490
rect 15680 10480 15820 10510
rect 15680 10460 15710 10480
rect 15790 10460 15820 10480
rect 15900 10460 15930 10490
rect 15570 10240 15600 10260
rect 15500 10210 15600 10240
rect 15680 10230 15710 10260
rect 15790 10230 15820 10260
rect 15900 10240 15930 10260
rect 15900 10210 16000 10240
rect 15500 10170 15510 10210
rect 15550 10170 15560 10210
rect 15500 10150 15560 10170
rect 15940 10170 15950 10210
rect 15990 10170 16000 10210
rect 15940 10150 16000 10170
rect 11700 10030 11800 10060
rect 11880 10030 11980 10060
rect 12060 10030 12160 10060
rect 12240 10030 12340 10060
rect 12420 10030 12520 10060
rect 12600 10030 12700 10060
rect 12780 10030 12880 10060
rect 12960 10030 13060 10060
rect 13140 10030 13240 10060
rect 13320 10030 13420 10060
rect 13500 10030 13600 10060
rect 13680 10030 13780 10060
rect 13860 10030 13960 10060
rect 14040 10030 14140 10060
rect 14220 10030 14320 10060
rect 14400 10030 14500 10060
rect 14580 10030 14680 10060
rect 14760 10030 14860 10060
rect 11620 10010 11800 10030
rect 11620 9970 11640 10010
rect 11680 10000 11800 10010
rect 14760 10010 14940 10030
rect 14760 10000 14880 10010
rect 11680 9970 11700 10000
rect 11620 9950 11700 9970
rect 14860 9970 14880 10000
rect 14920 9970 14940 10010
rect 14860 9950 14940 9970
rect 11806 9742 11864 9760
rect 11806 9708 11818 9742
rect 11852 9708 11864 9742
rect 11806 9690 11864 9708
rect 11916 9742 11974 9760
rect 11916 9708 11928 9742
rect 11962 9708 11974 9742
rect 11916 9690 11974 9708
rect 12026 9742 12084 9760
rect 12026 9708 12038 9742
rect 12072 9708 12084 9742
rect 12026 9690 12084 9708
rect 12136 9742 12194 9760
rect 12136 9708 12148 9742
rect 12182 9708 12194 9742
rect 12136 9690 12194 9708
rect 12246 9742 12304 9760
rect 12246 9708 12258 9742
rect 12292 9708 12304 9742
rect 12246 9690 12304 9708
rect 12356 9742 12414 9760
rect 12356 9708 12368 9742
rect 12402 9708 12414 9742
rect 12356 9690 12414 9708
rect 12466 9742 12524 9760
rect 12466 9708 12478 9742
rect 12512 9708 12524 9742
rect 12466 9690 12524 9708
rect 12576 9742 12634 9760
rect 12576 9708 12588 9742
rect 12622 9708 12634 9742
rect 12576 9690 12634 9708
rect 12686 9742 12744 9760
rect 12686 9708 12698 9742
rect 12732 9708 12744 9742
rect 12686 9690 12744 9708
rect 12796 9742 12854 9760
rect 12796 9708 12808 9742
rect 12842 9708 12854 9742
rect 12796 9690 12854 9708
rect 13706 9742 13764 9760
rect 13706 9708 13718 9742
rect 13752 9708 13764 9742
rect 13706 9690 13764 9708
rect 13816 9742 13874 9760
rect 13816 9708 13828 9742
rect 13862 9708 13874 9742
rect 13816 9690 13874 9708
rect 13926 9742 13984 9760
rect 13926 9708 13938 9742
rect 13972 9708 13984 9742
rect 13926 9690 13984 9708
rect 14036 9742 14094 9760
rect 14036 9708 14048 9742
rect 14082 9708 14094 9742
rect 14036 9690 14094 9708
rect 14146 9742 14204 9760
rect 14146 9708 14158 9742
rect 14192 9708 14204 9742
rect 14146 9690 14204 9708
rect 14256 9742 14314 9760
rect 14256 9708 14268 9742
rect 14302 9708 14314 9742
rect 14256 9690 14314 9708
rect 14366 9742 14424 9760
rect 14366 9708 14378 9742
rect 14412 9708 14424 9742
rect 14366 9690 14424 9708
rect 14476 9742 14534 9760
rect 14476 9708 14488 9742
rect 14522 9708 14534 9742
rect 14476 9690 14534 9708
rect 14586 9742 14644 9760
rect 14586 9708 14598 9742
rect 14632 9708 14644 9742
rect 14586 9690 14644 9708
rect 14696 9742 14754 9760
rect 14696 9708 14708 9742
rect 14742 9708 14754 9742
rect 14696 9690 14754 9708
rect 11710 9660 11740 9690
rect 11820 9660 11850 9690
rect 11930 9660 11960 9690
rect 12040 9660 12070 9690
rect 12150 9660 12180 9690
rect 12260 9660 12290 9690
rect 12370 9660 12400 9690
rect 12480 9660 12510 9690
rect 12590 9660 12620 9690
rect 12700 9660 12730 9690
rect 12810 9660 12840 9690
rect 12920 9660 12950 9690
rect 13610 9660 13640 9690
rect 13720 9660 13750 9690
rect 13830 9660 13860 9690
rect 13940 9660 13970 9690
rect 14050 9660 14080 9690
rect 14160 9660 14190 9690
rect 14270 9660 14300 9690
rect 14380 9660 14410 9690
rect 14490 9660 14520 9690
rect 14600 9660 14630 9690
rect 14710 9660 14740 9690
rect 14820 9660 14850 9690
rect 11710 9430 11740 9460
rect 11820 9430 11850 9460
rect 11930 9430 11960 9460
rect 12040 9430 12070 9460
rect 12150 9430 12180 9460
rect 12260 9430 12290 9460
rect 12370 9430 12400 9460
rect 12480 9430 12510 9460
rect 12590 9430 12620 9460
rect 12700 9430 12730 9460
rect 12810 9430 12840 9460
rect 12920 9430 12950 9460
rect 13610 9430 13640 9460
rect 13720 9430 13750 9460
rect 13830 9430 13860 9460
rect 13940 9430 13970 9460
rect 14050 9430 14080 9460
rect 14160 9430 14190 9460
rect 14270 9430 14300 9460
rect 14380 9430 14410 9460
rect 14490 9430 14520 9460
rect 14600 9430 14630 9460
rect 14710 9430 14740 9460
rect 14820 9430 14850 9460
rect 11630 9410 11740 9430
rect 11630 9370 11650 9410
rect 11690 9400 11740 9410
rect 12920 9410 13030 9430
rect 12920 9400 12970 9410
rect 11690 9370 11710 9400
rect 11630 9350 11710 9370
rect 12950 9370 12970 9400
rect 13010 9370 13030 9410
rect 12950 9350 13030 9370
rect 13530 9410 13640 9430
rect 13530 9370 13550 9410
rect 13590 9400 13640 9410
rect 14820 9410 14930 9430
rect 14820 9400 14870 9410
rect 13590 9370 13610 9400
rect 13530 9350 13610 9370
rect 14850 9370 14870 9400
rect 14910 9370 14930 9410
rect 14850 9350 14930 9370
<< polycont >>
rect 11340 13990 11380 14030
rect 11500 13990 11540 14030
rect 11660 13990 11700 14030
rect 11820 13990 11860 14030
rect 11980 13990 12020 14030
rect 12140 13990 12180 14030
rect 12300 13990 12340 14030
rect 12460 13990 12500 14030
rect 12620 13990 12660 14030
rect 12780 13990 12820 14030
rect 12940 13990 12980 14030
rect 13100 13990 13140 14030
rect 13420 13990 13460 14030
rect 13580 13990 13620 14030
rect 13740 13990 13780 14030
rect 13900 13990 13940 14030
rect 14060 13990 14100 14030
rect 14220 13990 14260 14030
rect 14380 13990 14420 14030
rect 14540 13990 14580 14030
rect 14700 13990 14740 14030
rect 14860 13990 14900 14030
rect 15020 13990 15060 14030
rect 15180 13990 15220 14030
rect 10940 13080 10980 13120
rect 11180 13080 11220 13120
rect 11420 13080 11460 13120
rect 11660 13080 11700 13120
rect 12300 13080 12340 13120
rect 12540 13080 12580 13120
rect 12780 13080 12820 13120
rect 13740 13080 13780 13120
rect 13980 13080 14020 13120
rect 14220 13080 14260 13120
rect 14860 13080 14900 13120
rect 15100 13080 15140 13120
rect 15340 13080 15380 13120
rect 15580 13080 15620 13120
rect 11443 12708 11477 12742
rect 11803 12708 11837 12742
rect 11923 12708 11957 12742
rect 12283 12708 12317 12742
rect 12403 12708 12437 12742
rect 11544 12478 11578 12512
rect 11702 12478 11736 12512
rect 12026 12478 12060 12512
rect 12180 12478 12214 12512
rect 12504 12478 12538 12512
rect 14123 12708 14157 12742
rect 14243 12708 14277 12742
rect 14603 12708 14637 12742
rect 14723 12708 14757 12742
rect 15083 12708 15117 12742
rect 14022 12478 14056 12512
rect 14346 12478 14380 12512
rect 14500 12478 14534 12512
rect 14824 12478 14858 12512
rect 14982 12478 15016 12512
rect 10720 11880 10760 11920
rect 10900 11870 10940 11910
rect 11380 11870 11420 11910
rect 11620 11870 11660 11910
rect 12100 11870 12140 11910
rect 12340 11870 12380 11910
rect 12760 11870 12800 11910
rect 13760 11870 13800 11910
rect 14180 11870 14220 11910
rect 14420 11870 14460 11910
rect 14900 11870 14940 11910
rect 15140 11870 15180 11910
rect 15620 11870 15660 11910
rect 15800 11880 15840 11920
rect 10540 11530 10580 11570
rect 12940 11530 12980 11570
rect 13580 11530 13620 11570
rect 15980 11530 16020 11570
rect 11910 10710 11950 10750
rect 12090 10710 12130 10750
rect 12270 10710 12310 10750
rect 12450 10710 12490 10750
rect 12630 10710 12670 10750
rect 12810 10710 12850 10750
rect 12990 10710 13030 10750
rect 13170 10710 13210 10750
rect 13350 10710 13390 10750
rect 13530 10710 13570 10750
rect 13710 10710 13750 10750
rect 13890 10710 13930 10750
rect 14070 10710 14110 10750
rect 14250 10710 14290 10750
rect 14430 10710 14470 10750
rect 14610 10710 14650 10750
rect 15730 10510 15770 10550
rect 15510 10170 15550 10210
rect 15950 10170 15990 10210
rect 11640 9970 11680 10010
rect 14880 9970 14920 10010
rect 11818 9708 11852 9742
rect 11928 9708 11962 9742
rect 12038 9708 12072 9742
rect 12148 9708 12182 9742
rect 12258 9708 12292 9742
rect 12368 9708 12402 9742
rect 12478 9708 12512 9742
rect 12588 9708 12622 9742
rect 12698 9708 12732 9742
rect 12808 9708 12842 9742
rect 13718 9708 13752 9742
rect 13828 9708 13862 9742
rect 13938 9708 13972 9742
rect 14048 9708 14082 9742
rect 14158 9708 14192 9742
rect 14268 9708 14302 9742
rect 14378 9708 14412 9742
rect 14488 9708 14522 9742
rect 14598 9708 14632 9742
rect 14708 9708 14742 9742
rect 11650 9370 11690 9410
rect 12970 9370 13010 9410
rect 13550 9370 13590 9410
rect 14870 9370 14910 9410
<< xpolycontact >>
rect 8454 18026 8524 18458
rect 8454 17216 8524 17648
rect 9241 18029 9311 18461
rect 9573 16817 9643 17249
rect 10686 18026 10756 18458
rect 10354 16286 10424 16718
rect 15674 18026 15744 18458
rect 16006 16286 16076 16718
rect 16787 18023 16857 18455
rect 16787 17423 16857 17855
rect 17574 18026 17644 18458
rect 17574 17216 17644 17648
rect 12632 14540 13072 14610
rect 13500 14540 13940 14610
<< ppolyres >>
rect 8454 17648 8524 18026
rect 17574 17648 17644 18026
<< xpolyres >>
rect 9241 17423 9311 18029
rect 9407 17855 9643 17925
rect 9407 17423 9477 17855
rect 9241 17353 9477 17423
rect 9573 17249 9643 17855
rect 10354 17852 10590 17922
rect 10354 16718 10424 17852
rect 10520 16892 10590 17852
rect 10686 16892 10756 18026
rect 10520 16822 10756 16892
rect 15674 16892 15744 18026
rect 15840 17852 16076 17922
rect 15840 16892 15910 17852
rect 15674 16822 15910 16892
rect 16006 16718 16076 17852
rect 16787 17855 16857 18023
rect 13072 14540 13500 14610
<< locali >>
rect 13240 19070 13320 19090
rect 13240 19030 13260 19070
rect 13300 19030 13320 19070
rect 13240 18990 13320 19030
rect 13240 18950 13260 18990
rect 13300 18950 13320 18990
rect 13240 18910 13320 18950
rect 13240 18870 13260 18910
rect 13300 18870 13320 18910
rect 12560 18784 12640 18790
rect 13240 18784 13320 18870
rect 13920 18784 14000 18790
rect 11276 18752 15284 18784
rect 11276 18718 11410 18752
rect 11444 18718 11500 18752
rect 11534 18718 11590 18752
rect 11624 18718 11680 18752
rect 11714 18718 11770 18752
rect 11804 18718 11860 18752
rect 11894 18718 11950 18752
rect 11984 18718 12040 18752
rect 12074 18718 12130 18752
rect 12164 18718 12220 18752
rect 12254 18718 12310 18752
rect 12344 18718 12400 18752
rect 12434 18718 12770 18752
rect 12804 18718 12860 18752
rect 12894 18718 12950 18752
rect 12984 18718 13040 18752
rect 13074 18718 13130 18752
rect 13164 18718 13220 18752
rect 13254 18718 13310 18752
rect 13344 18718 13400 18752
rect 13434 18718 13490 18752
rect 13524 18718 13580 18752
rect 13614 18718 13670 18752
rect 13704 18718 13760 18752
rect 13794 18718 14130 18752
rect 14164 18718 14220 18752
rect 14254 18718 14310 18752
rect 14344 18718 14400 18752
rect 14434 18718 14490 18752
rect 14524 18718 14580 18752
rect 14614 18718 14670 18752
rect 14704 18718 14760 18752
rect 14794 18718 14850 18752
rect 14884 18718 14940 18752
rect 14974 18718 15030 18752
rect 15064 18718 15120 18752
rect 15154 18718 15284 18752
rect 11276 18685 15284 18718
rect 11276 18668 11375 18685
rect 11276 18634 11309 18668
rect 11343 18634 11375 18668
rect 8450 18610 8530 18630
rect 8450 18597 8470 18610
rect 8510 18597 8530 18610
rect 9240 18610 9320 18630
rect 9240 18600 9260 18610
rect 9300 18600 9320 18610
rect 10680 18610 10760 18630
rect 8263 18563 8359 18597
rect 8619 18563 8715 18597
rect 8263 18501 8297 18563
rect 8450 18550 8530 18563
rect 8681 18501 8715 18563
rect 8263 17111 8297 17173
rect 8681 17111 8715 17173
rect 8263 17077 8359 17111
rect 8619 17077 8715 17111
rect 9050 18566 9146 18600
rect 9738 18566 9834 18600
rect 10680 18597 10700 18610
rect 10740 18597 10760 18610
rect 9050 18504 9084 18566
rect 9240 18550 9320 18566
rect 9800 18504 9834 18566
rect 9050 16712 9084 16774
rect 9800 16712 9834 16774
rect 9050 16678 9146 16712
rect 9738 16678 9834 16712
rect 10163 18563 10259 18597
rect 10851 18563 10947 18597
rect 10163 18501 10197 18563
rect 10680 18550 10760 18563
rect 10913 18501 10947 18563
rect 10163 16181 10197 16243
rect 11276 18578 11375 18634
rect 12465 18668 12735 18685
rect 12465 18634 12496 18668
rect 12530 18634 12669 18668
rect 12703 18634 12735 18668
rect 11276 18544 11309 18578
rect 11343 18544 11375 18578
rect 11276 18488 11375 18544
rect 11276 18454 11309 18488
rect 11343 18454 11375 18488
rect 11276 18398 11375 18454
rect 11276 18364 11309 18398
rect 11343 18364 11375 18398
rect 11276 18308 11375 18364
rect 11276 18274 11309 18308
rect 11343 18274 11375 18308
rect 11276 18218 11375 18274
rect 11276 18184 11309 18218
rect 11343 18184 11375 18218
rect 11276 18128 11375 18184
rect 11276 18094 11309 18128
rect 11343 18094 11375 18128
rect 11276 18038 11375 18094
rect 11276 18004 11309 18038
rect 11343 18004 11375 18038
rect 11276 17948 11375 18004
rect 11276 17914 11309 17948
rect 11343 17914 11375 17948
rect 11276 17858 11375 17914
rect 11276 17824 11309 17858
rect 11343 17824 11375 17858
rect 11276 17768 11375 17824
rect 11276 17740 11309 17768
rect 11270 17734 11309 17740
rect 11343 17740 11375 17768
rect 11439 18602 12401 18621
rect 11439 18568 11550 18602
rect 11584 18568 11640 18602
rect 11674 18568 11730 18602
rect 11764 18568 11820 18602
rect 11854 18568 11910 18602
rect 11944 18568 12000 18602
rect 12034 18568 12090 18602
rect 12124 18568 12180 18602
rect 12214 18568 12270 18602
rect 12304 18568 12401 18602
rect 11439 18549 12401 18568
rect 11439 18508 11511 18549
rect 11439 18474 11458 18508
rect 11492 18474 11511 18508
rect 12329 18489 12401 18549
rect 11439 18418 11511 18474
rect 11439 18384 11458 18418
rect 11492 18384 11511 18418
rect 11439 18328 11511 18384
rect 11439 18294 11458 18328
rect 11492 18294 11511 18328
rect 11439 18238 11511 18294
rect 11439 18204 11458 18238
rect 11492 18204 11511 18238
rect 11439 18148 11511 18204
rect 11439 18114 11458 18148
rect 11492 18114 11511 18148
rect 11439 18058 11511 18114
rect 11439 18024 11458 18058
rect 11492 18024 11511 18058
rect 11439 17968 11511 18024
rect 11439 17934 11458 17968
rect 11492 17934 11511 17968
rect 11439 17878 11511 17934
rect 11439 17844 11458 17878
rect 11492 17844 11511 17878
rect 11439 17788 11511 17844
rect 11573 18426 12267 18487
rect 11573 18392 11632 18426
rect 11666 18414 11722 18426
rect 11694 18392 11722 18414
rect 11756 18414 11812 18426
rect 11756 18392 11760 18414
rect 11573 18380 11660 18392
rect 11694 18380 11760 18392
rect 11794 18392 11812 18414
rect 11846 18414 11902 18426
rect 11846 18392 11860 18414
rect 11794 18380 11860 18392
rect 11894 18392 11902 18414
rect 11936 18414 11992 18426
rect 12026 18414 12082 18426
rect 12116 18414 12172 18426
rect 11936 18392 11960 18414
rect 12026 18392 12060 18414
rect 12116 18392 12160 18414
rect 12206 18392 12267 18426
rect 11894 18380 11960 18392
rect 11994 18380 12060 18392
rect 12094 18380 12160 18392
rect 12194 18380 12267 18392
rect 11573 18336 12267 18380
rect 11573 18302 11632 18336
rect 11666 18314 11722 18336
rect 11694 18302 11722 18314
rect 11756 18314 11812 18336
rect 11756 18302 11760 18314
rect 11573 18280 11660 18302
rect 11694 18280 11760 18302
rect 11794 18302 11812 18314
rect 11846 18314 11902 18336
rect 11846 18302 11860 18314
rect 11794 18280 11860 18302
rect 11894 18302 11902 18314
rect 11936 18314 11992 18336
rect 12026 18314 12082 18336
rect 12116 18314 12172 18336
rect 11936 18302 11960 18314
rect 12026 18302 12060 18314
rect 12116 18302 12160 18314
rect 12206 18302 12267 18336
rect 11894 18280 11960 18302
rect 11994 18280 12060 18302
rect 12094 18280 12160 18302
rect 12194 18280 12267 18302
rect 11573 18246 12267 18280
rect 11573 18212 11632 18246
rect 11666 18214 11722 18246
rect 11694 18212 11722 18214
rect 11756 18214 11812 18246
rect 11756 18212 11760 18214
rect 11573 18180 11660 18212
rect 11694 18180 11760 18212
rect 11794 18212 11812 18214
rect 11846 18214 11902 18246
rect 11846 18212 11860 18214
rect 11794 18180 11860 18212
rect 11894 18212 11902 18214
rect 11936 18214 11992 18246
rect 12026 18214 12082 18246
rect 12116 18214 12172 18246
rect 11936 18212 11960 18214
rect 12026 18212 12060 18214
rect 12116 18212 12160 18214
rect 12206 18212 12267 18246
rect 11894 18180 11960 18212
rect 11994 18180 12060 18212
rect 12094 18180 12160 18212
rect 12194 18180 12267 18212
rect 11573 18156 12267 18180
rect 11573 18122 11632 18156
rect 11666 18122 11722 18156
rect 11756 18122 11812 18156
rect 11846 18122 11902 18156
rect 11936 18122 11992 18156
rect 12026 18122 12082 18156
rect 12116 18122 12172 18156
rect 12206 18122 12267 18156
rect 11573 18114 12267 18122
rect 11573 18080 11660 18114
rect 11694 18080 11760 18114
rect 11794 18080 11860 18114
rect 11894 18080 11960 18114
rect 11994 18080 12060 18114
rect 12094 18080 12160 18114
rect 12194 18080 12267 18114
rect 11573 18066 12267 18080
rect 11573 18032 11632 18066
rect 11666 18032 11722 18066
rect 11756 18032 11812 18066
rect 11846 18032 11902 18066
rect 11936 18032 11992 18066
rect 12026 18032 12082 18066
rect 12116 18032 12172 18066
rect 12206 18032 12267 18066
rect 11573 18014 12267 18032
rect 11573 17980 11660 18014
rect 11694 17980 11760 18014
rect 11794 17980 11860 18014
rect 11894 17980 11960 18014
rect 11994 17980 12060 18014
rect 12094 17980 12160 18014
rect 12194 17980 12267 18014
rect 11573 17976 12267 17980
rect 11573 17942 11632 17976
rect 11666 17942 11722 17976
rect 11756 17942 11812 17976
rect 11846 17942 11902 17976
rect 11936 17942 11992 17976
rect 12026 17942 12082 17976
rect 12116 17942 12172 17976
rect 12206 17942 12267 17976
rect 11573 17914 12267 17942
rect 11573 17886 11660 17914
rect 11694 17886 11760 17914
rect 11573 17852 11632 17886
rect 11694 17880 11722 17886
rect 11666 17852 11722 17880
rect 11756 17880 11760 17886
rect 11794 17886 11860 17914
rect 11794 17880 11812 17886
rect 11756 17852 11812 17880
rect 11846 17880 11860 17886
rect 11894 17886 11960 17914
rect 11994 17886 12060 17914
rect 12094 17886 12160 17914
rect 12194 17886 12267 17914
rect 11894 17880 11902 17886
rect 11846 17852 11902 17880
rect 11936 17880 11960 17886
rect 12026 17880 12060 17886
rect 12116 17880 12160 17886
rect 11936 17852 11992 17880
rect 12026 17852 12082 17880
rect 12116 17852 12172 17880
rect 12206 17852 12267 17886
rect 11573 17793 12267 17852
rect 12329 18455 12348 18489
rect 12382 18455 12401 18489
rect 12329 18399 12401 18455
rect 12329 18365 12348 18399
rect 12382 18365 12401 18399
rect 12329 18309 12401 18365
rect 12329 18275 12348 18309
rect 12382 18275 12401 18309
rect 12329 18219 12401 18275
rect 12329 18185 12348 18219
rect 12382 18185 12401 18219
rect 12329 18129 12401 18185
rect 12329 18095 12348 18129
rect 12382 18095 12401 18129
rect 12329 18039 12401 18095
rect 12329 18005 12348 18039
rect 12382 18005 12401 18039
rect 12329 17949 12401 18005
rect 12329 17915 12348 17949
rect 12382 17915 12401 17949
rect 12329 17859 12401 17915
rect 12329 17825 12348 17859
rect 12382 17825 12401 17859
rect 11439 17754 11458 17788
rect 11492 17754 11511 17788
rect 11439 17740 11511 17754
rect 12329 17769 12401 17825
rect 12329 17740 12348 17769
rect 11343 17735 12348 17740
rect 12382 17740 12401 17769
rect 12465 18578 12735 18634
rect 13825 18668 14095 18685
rect 13825 18634 13856 18668
rect 13890 18634 14029 18668
rect 14063 18634 14095 18668
rect 12465 18544 12496 18578
rect 12530 18544 12669 18578
rect 12703 18544 12735 18578
rect 12465 18488 12735 18544
rect 12465 18454 12496 18488
rect 12530 18454 12669 18488
rect 12703 18454 12735 18488
rect 12465 18398 12735 18454
rect 12465 18364 12496 18398
rect 12530 18364 12669 18398
rect 12703 18364 12735 18398
rect 12465 18308 12735 18364
rect 12465 18274 12496 18308
rect 12530 18274 12669 18308
rect 12703 18274 12735 18308
rect 12465 18218 12735 18274
rect 12465 18184 12496 18218
rect 12530 18184 12669 18218
rect 12703 18184 12735 18218
rect 12465 18128 12735 18184
rect 12465 18094 12496 18128
rect 12530 18094 12669 18128
rect 12703 18094 12735 18128
rect 12465 18038 12735 18094
rect 12465 18004 12496 18038
rect 12530 18004 12669 18038
rect 12703 18004 12735 18038
rect 12465 17948 12735 18004
rect 12465 17914 12496 17948
rect 12530 17914 12669 17948
rect 12703 17914 12735 17948
rect 12465 17858 12735 17914
rect 12465 17824 12496 17858
rect 12530 17824 12669 17858
rect 12703 17824 12735 17858
rect 12465 17768 12735 17824
rect 12465 17740 12496 17768
rect 12382 17735 12496 17740
rect 11343 17734 12496 17735
rect 12530 17734 12669 17768
rect 12703 17740 12735 17768
rect 12799 18602 13761 18621
rect 12799 18568 12910 18602
rect 12944 18568 13000 18602
rect 13034 18568 13090 18602
rect 13124 18568 13180 18602
rect 13214 18568 13270 18602
rect 13304 18568 13360 18602
rect 13394 18568 13450 18602
rect 13484 18568 13540 18602
rect 13574 18568 13630 18602
rect 13664 18568 13761 18602
rect 12799 18549 13761 18568
rect 12799 18508 12871 18549
rect 12799 18474 12818 18508
rect 12852 18474 12871 18508
rect 13689 18489 13761 18549
rect 12799 18418 12871 18474
rect 12799 18384 12818 18418
rect 12852 18384 12871 18418
rect 12799 18328 12871 18384
rect 12799 18294 12818 18328
rect 12852 18294 12871 18328
rect 12799 18238 12871 18294
rect 12799 18204 12818 18238
rect 12852 18204 12871 18238
rect 12799 18148 12871 18204
rect 12799 18114 12818 18148
rect 12852 18114 12871 18148
rect 12799 18058 12871 18114
rect 12799 18024 12818 18058
rect 12852 18024 12871 18058
rect 12799 17968 12871 18024
rect 12799 17934 12818 17968
rect 12852 17934 12871 17968
rect 12799 17878 12871 17934
rect 12799 17844 12818 17878
rect 12852 17844 12871 17878
rect 12799 17788 12871 17844
rect 12933 18426 13627 18487
rect 12933 18392 12992 18426
rect 13026 18414 13082 18426
rect 13054 18392 13082 18414
rect 13116 18414 13172 18426
rect 13116 18392 13120 18414
rect 12933 18380 13020 18392
rect 13054 18380 13120 18392
rect 13154 18392 13172 18414
rect 13206 18414 13262 18426
rect 13206 18392 13220 18414
rect 13154 18380 13220 18392
rect 13254 18392 13262 18414
rect 13296 18414 13352 18426
rect 13386 18414 13442 18426
rect 13476 18414 13532 18426
rect 13296 18392 13320 18414
rect 13386 18392 13420 18414
rect 13476 18392 13520 18414
rect 13566 18392 13627 18426
rect 13254 18380 13320 18392
rect 13354 18380 13420 18392
rect 13454 18380 13520 18392
rect 13554 18380 13627 18392
rect 12933 18336 13627 18380
rect 12933 18302 12992 18336
rect 13026 18314 13082 18336
rect 13054 18302 13082 18314
rect 13116 18314 13172 18336
rect 13116 18302 13120 18314
rect 12933 18280 13020 18302
rect 13054 18280 13120 18302
rect 13154 18302 13172 18314
rect 13206 18314 13262 18336
rect 13206 18302 13220 18314
rect 13154 18280 13220 18302
rect 13254 18302 13262 18314
rect 13296 18314 13352 18336
rect 13386 18314 13442 18336
rect 13476 18314 13532 18336
rect 13296 18302 13320 18314
rect 13386 18302 13420 18314
rect 13476 18302 13520 18314
rect 13566 18302 13627 18336
rect 13254 18280 13320 18302
rect 13354 18280 13420 18302
rect 13454 18280 13520 18302
rect 13554 18280 13627 18302
rect 12933 18246 13627 18280
rect 12933 18212 12992 18246
rect 13026 18214 13082 18246
rect 13054 18212 13082 18214
rect 13116 18214 13172 18246
rect 13116 18212 13120 18214
rect 12933 18180 13020 18212
rect 13054 18180 13120 18212
rect 13154 18212 13172 18214
rect 13206 18214 13262 18246
rect 13206 18212 13220 18214
rect 13154 18180 13220 18212
rect 13254 18212 13262 18214
rect 13296 18214 13352 18246
rect 13386 18214 13442 18246
rect 13476 18214 13532 18246
rect 13296 18212 13320 18214
rect 13386 18212 13420 18214
rect 13476 18212 13520 18214
rect 13566 18212 13627 18246
rect 13254 18180 13320 18212
rect 13354 18180 13420 18212
rect 13454 18180 13520 18212
rect 13554 18180 13627 18212
rect 12933 18156 13627 18180
rect 12933 18122 12992 18156
rect 13026 18122 13082 18156
rect 13116 18122 13172 18156
rect 13206 18122 13262 18156
rect 13296 18122 13352 18156
rect 13386 18122 13442 18156
rect 13476 18122 13532 18156
rect 13566 18122 13627 18156
rect 12933 18114 13627 18122
rect 12933 18080 13020 18114
rect 13054 18080 13120 18114
rect 13154 18080 13220 18114
rect 13254 18080 13320 18114
rect 13354 18080 13420 18114
rect 13454 18080 13520 18114
rect 13554 18080 13627 18114
rect 12933 18066 13627 18080
rect 12933 18032 12992 18066
rect 13026 18032 13082 18066
rect 13116 18032 13172 18066
rect 13206 18032 13262 18066
rect 13296 18032 13352 18066
rect 13386 18032 13442 18066
rect 13476 18032 13532 18066
rect 13566 18032 13627 18066
rect 12933 18014 13627 18032
rect 12933 17980 13020 18014
rect 13054 17980 13120 18014
rect 13154 17980 13220 18014
rect 13254 17980 13320 18014
rect 13354 17980 13420 18014
rect 13454 17980 13520 18014
rect 13554 17980 13627 18014
rect 12933 17976 13627 17980
rect 12933 17942 12992 17976
rect 13026 17942 13082 17976
rect 13116 17942 13172 17976
rect 13206 17942 13262 17976
rect 13296 17942 13352 17976
rect 13386 17942 13442 17976
rect 13476 17942 13532 17976
rect 13566 17942 13627 17976
rect 12933 17914 13627 17942
rect 12933 17886 13020 17914
rect 13054 17886 13120 17914
rect 12933 17852 12992 17886
rect 13054 17880 13082 17886
rect 13026 17852 13082 17880
rect 13116 17880 13120 17886
rect 13154 17886 13220 17914
rect 13154 17880 13172 17886
rect 13116 17852 13172 17880
rect 13206 17880 13220 17886
rect 13254 17886 13320 17914
rect 13354 17886 13420 17914
rect 13454 17886 13520 17914
rect 13554 17886 13627 17914
rect 13254 17880 13262 17886
rect 13206 17852 13262 17880
rect 13296 17880 13320 17886
rect 13386 17880 13420 17886
rect 13476 17880 13520 17886
rect 13296 17852 13352 17880
rect 13386 17852 13442 17880
rect 13476 17852 13532 17880
rect 13566 17852 13627 17886
rect 12933 17793 13627 17852
rect 13689 18455 13708 18489
rect 13742 18455 13761 18489
rect 13689 18399 13761 18455
rect 13689 18365 13708 18399
rect 13742 18365 13761 18399
rect 13689 18309 13761 18365
rect 13689 18275 13708 18309
rect 13742 18275 13761 18309
rect 13689 18219 13761 18275
rect 13689 18185 13708 18219
rect 13742 18185 13761 18219
rect 13689 18129 13761 18185
rect 13689 18095 13708 18129
rect 13742 18095 13761 18129
rect 13689 18039 13761 18095
rect 13689 18005 13708 18039
rect 13742 18005 13761 18039
rect 13689 17949 13761 18005
rect 13689 17915 13708 17949
rect 13742 17915 13761 17949
rect 13689 17859 13761 17915
rect 13689 17825 13708 17859
rect 13742 17825 13761 17859
rect 12799 17754 12818 17788
rect 12852 17754 12871 17788
rect 12799 17740 12871 17754
rect 13689 17769 13761 17825
rect 13689 17740 13708 17769
rect 12703 17735 13708 17740
rect 13742 17740 13761 17769
rect 13825 18578 14095 18634
rect 15185 18668 15284 18685
rect 15185 18634 15216 18668
rect 15250 18634 15284 18668
rect 13825 18544 13856 18578
rect 13890 18544 14029 18578
rect 14063 18544 14095 18578
rect 13825 18488 14095 18544
rect 13825 18454 13856 18488
rect 13890 18454 14029 18488
rect 14063 18454 14095 18488
rect 13825 18398 14095 18454
rect 13825 18364 13856 18398
rect 13890 18364 14029 18398
rect 14063 18364 14095 18398
rect 13825 18308 14095 18364
rect 13825 18274 13856 18308
rect 13890 18274 14029 18308
rect 14063 18274 14095 18308
rect 13825 18218 14095 18274
rect 13825 18184 13856 18218
rect 13890 18184 14029 18218
rect 14063 18184 14095 18218
rect 13825 18128 14095 18184
rect 13825 18094 13856 18128
rect 13890 18094 14029 18128
rect 14063 18094 14095 18128
rect 13825 18038 14095 18094
rect 13825 18004 13856 18038
rect 13890 18004 14029 18038
rect 14063 18004 14095 18038
rect 13825 17948 14095 18004
rect 13825 17914 13856 17948
rect 13890 17914 14029 17948
rect 14063 17914 14095 17948
rect 13825 17858 14095 17914
rect 13825 17824 13856 17858
rect 13890 17824 14029 17858
rect 14063 17824 14095 17858
rect 13825 17768 14095 17824
rect 13825 17740 13856 17768
rect 13742 17735 13856 17740
rect 12703 17734 13856 17735
rect 13890 17734 14029 17768
rect 14063 17740 14095 17768
rect 14159 18602 15121 18621
rect 14159 18568 14270 18602
rect 14304 18568 14360 18602
rect 14394 18568 14450 18602
rect 14484 18568 14540 18602
rect 14574 18568 14630 18602
rect 14664 18568 14720 18602
rect 14754 18568 14810 18602
rect 14844 18568 14900 18602
rect 14934 18568 14990 18602
rect 15024 18568 15121 18602
rect 14159 18549 15121 18568
rect 14159 18508 14231 18549
rect 14159 18474 14178 18508
rect 14212 18474 14231 18508
rect 15049 18489 15121 18549
rect 14159 18418 14231 18474
rect 14159 18384 14178 18418
rect 14212 18384 14231 18418
rect 14159 18328 14231 18384
rect 14159 18294 14178 18328
rect 14212 18294 14231 18328
rect 14159 18238 14231 18294
rect 14159 18204 14178 18238
rect 14212 18204 14231 18238
rect 14159 18148 14231 18204
rect 14159 18114 14178 18148
rect 14212 18114 14231 18148
rect 14159 18058 14231 18114
rect 14159 18024 14178 18058
rect 14212 18024 14231 18058
rect 14159 17968 14231 18024
rect 14159 17934 14178 17968
rect 14212 17934 14231 17968
rect 14159 17878 14231 17934
rect 14159 17844 14178 17878
rect 14212 17844 14231 17878
rect 14159 17788 14231 17844
rect 14293 18426 14987 18487
rect 14293 18392 14352 18426
rect 14386 18414 14442 18426
rect 14414 18392 14442 18414
rect 14476 18414 14532 18426
rect 14476 18392 14480 18414
rect 14293 18380 14380 18392
rect 14414 18380 14480 18392
rect 14514 18392 14532 18414
rect 14566 18414 14622 18426
rect 14566 18392 14580 18414
rect 14514 18380 14580 18392
rect 14614 18392 14622 18414
rect 14656 18414 14712 18426
rect 14746 18414 14802 18426
rect 14836 18414 14892 18426
rect 14656 18392 14680 18414
rect 14746 18392 14780 18414
rect 14836 18392 14880 18414
rect 14926 18392 14987 18426
rect 14614 18380 14680 18392
rect 14714 18380 14780 18392
rect 14814 18380 14880 18392
rect 14914 18380 14987 18392
rect 14293 18336 14987 18380
rect 14293 18302 14352 18336
rect 14386 18314 14442 18336
rect 14414 18302 14442 18314
rect 14476 18314 14532 18336
rect 14476 18302 14480 18314
rect 14293 18280 14380 18302
rect 14414 18280 14480 18302
rect 14514 18302 14532 18314
rect 14566 18314 14622 18336
rect 14566 18302 14580 18314
rect 14514 18280 14580 18302
rect 14614 18302 14622 18314
rect 14656 18314 14712 18336
rect 14746 18314 14802 18336
rect 14836 18314 14892 18336
rect 14656 18302 14680 18314
rect 14746 18302 14780 18314
rect 14836 18302 14880 18314
rect 14926 18302 14987 18336
rect 14614 18280 14680 18302
rect 14714 18280 14780 18302
rect 14814 18280 14880 18302
rect 14914 18280 14987 18302
rect 14293 18246 14987 18280
rect 14293 18212 14352 18246
rect 14386 18214 14442 18246
rect 14414 18212 14442 18214
rect 14476 18214 14532 18246
rect 14476 18212 14480 18214
rect 14293 18180 14380 18212
rect 14414 18180 14480 18212
rect 14514 18212 14532 18214
rect 14566 18214 14622 18246
rect 14566 18212 14580 18214
rect 14514 18180 14580 18212
rect 14614 18212 14622 18214
rect 14656 18214 14712 18246
rect 14746 18214 14802 18246
rect 14836 18214 14892 18246
rect 14656 18212 14680 18214
rect 14746 18212 14780 18214
rect 14836 18212 14880 18214
rect 14926 18212 14987 18246
rect 14614 18180 14680 18212
rect 14714 18180 14780 18212
rect 14814 18180 14880 18212
rect 14914 18180 14987 18212
rect 14293 18156 14987 18180
rect 14293 18122 14352 18156
rect 14386 18122 14442 18156
rect 14476 18122 14532 18156
rect 14566 18122 14622 18156
rect 14656 18122 14712 18156
rect 14746 18122 14802 18156
rect 14836 18122 14892 18156
rect 14926 18122 14987 18156
rect 14293 18114 14987 18122
rect 14293 18080 14380 18114
rect 14414 18080 14480 18114
rect 14514 18080 14580 18114
rect 14614 18080 14680 18114
rect 14714 18080 14780 18114
rect 14814 18080 14880 18114
rect 14914 18080 14987 18114
rect 14293 18066 14987 18080
rect 14293 18032 14352 18066
rect 14386 18032 14442 18066
rect 14476 18032 14532 18066
rect 14566 18032 14622 18066
rect 14656 18032 14712 18066
rect 14746 18032 14802 18066
rect 14836 18032 14892 18066
rect 14926 18032 14987 18066
rect 14293 18014 14987 18032
rect 14293 17980 14380 18014
rect 14414 17980 14480 18014
rect 14514 17980 14580 18014
rect 14614 17980 14680 18014
rect 14714 17980 14780 18014
rect 14814 17980 14880 18014
rect 14914 17980 14987 18014
rect 14293 17976 14987 17980
rect 14293 17942 14352 17976
rect 14386 17942 14442 17976
rect 14476 17942 14532 17976
rect 14566 17942 14622 17976
rect 14656 17942 14712 17976
rect 14746 17942 14802 17976
rect 14836 17942 14892 17976
rect 14926 17942 14987 17976
rect 14293 17914 14987 17942
rect 14293 17886 14380 17914
rect 14414 17886 14480 17914
rect 14293 17852 14352 17886
rect 14414 17880 14442 17886
rect 14386 17852 14442 17880
rect 14476 17880 14480 17886
rect 14514 17886 14580 17914
rect 14514 17880 14532 17886
rect 14476 17852 14532 17880
rect 14566 17880 14580 17886
rect 14614 17886 14680 17914
rect 14714 17886 14780 17914
rect 14814 17886 14880 17914
rect 14914 17886 14987 17914
rect 14614 17880 14622 17886
rect 14566 17852 14622 17880
rect 14656 17880 14680 17886
rect 14746 17880 14780 17886
rect 14836 17880 14880 17886
rect 14656 17852 14712 17880
rect 14746 17852 14802 17880
rect 14836 17852 14892 17880
rect 14926 17852 14987 17886
rect 14293 17793 14987 17852
rect 15049 18455 15068 18489
rect 15102 18455 15121 18489
rect 15049 18399 15121 18455
rect 15049 18365 15068 18399
rect 15102 18365 15121 18399
rect 15049 18309 15121 18365
rect 15049 18275 15068 18309
rect 15102 18275 15121 18309
rect 15049 18219 15121 18275
rect 15049 18185 15068 18219
rect 15102 18185 15121 18219
rect 15049 18129 15121 18185
rect 15049 18095 15068 18129
rect 15102 18095 15121 18129
rect 15049 18039 15121 18095
rect 15049 18005 15068 18039
rect 15102 18005 15121 18039
rect 15049 17949 15121 18005
rect 15049 17915 15068 17949
rect 15102 17915 15121 17949
rect 15049 17859 15121 17915
rect 15049 17825 15068 17859
rect 15102 17825 15121 17859
rect 14159 17754 14178 17788
rect 14212 17754 14231 17788
rect 14159 17740 14231 17754
rect 15049 17769 15121 17825
rect 15049 17740 15068 17769
rect 14063 17735 15068 17740
rect 15102 17740 15121 17769
rect 15185 18578 15284 18634
rect 15670 18610 15750 18630
rect 15670 18597 15690 18610
rect 15730 18597 15750 18610
rect 16780 18610 16860 18630
rect 15185 18544 15216 18578
rect 15250 18544 15284 18578
rect 15185 18488 15284 18544
rect 15185 18454 15216 18488
rect 15250 18454 15284 18488
rect 15185 18398 15284 18454
rect 15185 18364 15216 18398
rect 15250 18364 15284 18398
rect 15185 18308 15284 18364
rect 15185 18274 15216 18308
rect 15250 18274 15284 18308
rect 15185 18218 15284 18274
rect 15185 18184 15216 18218
rect 15250 18184 15284 18218
rect 15185 18128 15284 18184
rect 15185 18094 15216 18128
rect 15250 18094 15284 18128
rect 15185 18038 15284 18094
rect 15185 18004 15216 18038
rect 15250 18004 15284 18038
rect 15185 17948 15284 18004
rect 15185 17914 15216 17948
rect 15250 17914 15284 17948
rect 15185 17858 15284 17914
rect 15185 17824 15216 17858
rect 15250 17824 15284 17858
rect 15185 17768 15284 17824
rect 15185 17740 15216 17768
rect 15102 17735 15216 17740
rect 14063 17734 15216 17735
rect 15250 17740 15284 17768
rect 15483 18563 15579 18597
rect 16171 18563 16267 18597
rect 16780 18594 16800 18610
rect 16840 18594 16860 18610
rect 17570 18610 17650 18630
rect 17570 18597 17590 18610
rect 17630 18597 17650 18610
rect 15483 18501 15517 18563
rect 15670 18550 15750 18563
rect 15250 17734 15290 17740
rect 11270 17712 15290 17734
rect 11270 17678 11516 17712
rect 11550 17678 11606 17712
rect 11640 17678 11696 17712
rect 11730 17678 11786 17712
rect 11820 17678 11876 17712
rect 11910 17678 11966 17712
rect 12000 17678 12056 17712
rect 12090 17678 12146 17712
rect 12180 17678 12236 17712
rect 12270 17678 12876 17712
rect 12910 17678 12966 17712
rect 13000 17678 13056 17712
rect 13090 17678 13146 17712
rect 13180 17678 13236 17712
rect 13270 17678 13326 17712
rect 13360 17678 13416 17712
rect 13450 17678 13506 17712
rect 13540 17678 13596 17712
rect 13630 17678 14236 17712
rect 14270 17678 14326 17712
rect 14360 17678 14416 17712
rect 14450 17678 14506 17712
rect 14540 17678 14596 17712
rect 14630 17678 14686 17712
rect 14720 17678 14776 17712
rect 14810 17678 14866 17712
rect 14900 17678 14956 17712
rect 14990 17678 15290 17712
rect 11270 17644 11309 17678
rect 11343 17644 12496 17678
rect 12530 17644 12669 17678
rect 12703 17644 13856 17678
rect 13890 17644 14029 17678
rect 14063 17644 15216 17678
rect 15250 17644 15290 17678
rect 11270 17588 15290 17644
rect 11270 17554 11309 17588
rect 11343 17565 12496 17588
rect 11343 17554 11410 17565
rect 11270 17531 11410 17554
rect 11444 17531 11500 17565
rect 11534 17531 11590 17565
rect 11624 17531 11680 17565
rect 11714 17531 11770 17565
rect 11804 17531 11860 17565
rect 11894 17531 11950 17565
rect 11984 17531 12040 17565
rect 12074 17531 12130 17565
rect 12164 17531 12220 17565
rect 12254 17531 12310 17565
rect 12344 17531 12400 17565
rect 12434 17554 12496 17565
rect 12530 17554 12669 17588
rect 12703 17565 13856 17588
rect 12703 17554 12770 17565
rect 12434 17531 12770 17554
rect 12804 17531 12860 17565
rect 12894 17531 12950 17565
rect 12984 17531 13040 17565
rect 13074 17531 13130 17565
rect 13164 17531 13220 17565
rect 13254 17531 13310 17565
rect 13344 17531 13400 17565
rect 13434 17531 13490 17565
rect 13524 17531 13580 17565
rect 13614 17531 13670 17565
rect 13704 17531 13760 17565
rect 13794 17554 13856 17565
rect 13890 17554 14029 17588
rect 14063 17565 15216 17588
rect 14063 17554 14130 17565
rect 13794 17531 14130 17554
rect 14164 17531 14220 17565
rect 14254 17531 14310 17565
rect 14344 17531 14400 17565
rect 14434 17531 14490 17565
rect 14524 17531 14580 17565
rect 14614 17531 14670 17565
rect 14704 17531 14760 17565
rect 14794 17531 14850 17565
rect 14884 17531 14940 17565
rect 14974 17531 15030 17565
rect 15064 17531 15120 17565
rect 15154 17554 15216 17565
rect 15250 17554 15290 17588
rect 15154 17531 15290 17554
rect 11270 17490 15290 17531
rect 12560 17424 12640 17490
rect 13920 17424 14000 17490
rect 11276 17392 15284 17424
rect 11276 17358 11410 17392
rect 11444 17358 11500 17392
rect 11534 17358 11590 17392
rect 11624 17358 11680 17392
rect 11714 17358 11770 17392
rect 11804 17358 11860 17392
rect 11894 17358 11950 17392
rect 11984 17358 12040 17392
rect 12074 17358 12130 17392
rect 12164 17358 12220 17392
rect 12254 17358 12310 17392
rect 12344 17358 12400 17392
rect 12434 17358 12770 17392
rect 12804 17358 12860 17392
rect 12894 17358 12950 17392
rect 12984 17358 13040 17392
rect 13074 17358 13130 17392
rect 13164 17358 13220 17392
rect 13254 17358 13310 17392
rect 13344 17358 13400 17392
rect 13434 17358 13490 17392
rect 13524 17358 13580 17392
rect 13614 17358 13670 17392
rect 13704 17358 13760 17392
rect 13794 17358 14130 17392
rect 14164 17358 14220 17392
rect 14254 17358 14310 17392
rect 14344 17358 14400 17392
rect 14434 17358 14490 17392
rect 14524 17358 14580 17392
rect 14614 17358 14670 17392
rect 14704 17358 14760 17392
rect 14794 17358 14850 17392
rect 14884 17358 14940 17392
rect 14974 17358 15030 17392
rect 15064 17358 15120 17392
rect 15154 17358 15284 17392
rect 11276 17325 15284 17358
rect 11276 17308 11375 17325
rect 11276 17274 11309 17308
rect 11343 17274 11375 17308
rect 11276 17218 11375 17274
rect 12465 17308 12735 17325
rect 12465 17274 12496 17308
rect 12530 17274 12669 17308
rect 12703 17274 12735 17308
rect 11276 17184 11309 17218
rect 11343 17184 11375 17218
rect 11276 17128 11375 17184
rect 11276 17094 11309 17128
rect 11343 17094 11375 17128
rect 11276 17038 11375 17094
rect 11276 17004 11309 17038
rect 11343 17004 11375 17038
rect 11276 16948 11375 17004
rect 11276 16914 11309 16948
rect 11343 16914 11375 16948
rect 11276 16858 11375 16914
rect 11276 16824 11309 16858
rect 11343 16824 11375 16858
rect 11276 16768 11375 16824
rect 11276 16734 11309 16768
rect 11343 16734 11375 16768
rect 11276 16678 11375 16734
rect 11276 16644 11309 16678
rect 11343 16644 11375 16678
rect 11276 16588 11375 16644
rect 11276 16554 11309 16588
rect 11343 16554 11375 16588
rect 11276 16498 11375 16554
rect 11276 16464 11309 16498
rect 11343 16464 11375 16498
rect 11276 16408 11375 16464
rect 11276 16380 11309 16408
rect 10913 16181 10947 16243
rect 10163 16147 10259 16181
rect 10851 16147 10947 16181
rect 11270 16374 11309 16380
rect 11343 16380 11375 16408
rect 11439 17242 12401 17261
rect 11439 17208 11550 17242
rect 11584 17208 11640 17242
rect 11674 17208 11730 17242
rect 11764 17208 11820 17242
rect 11854 17208 11910 17242
rect 11944 17208 12000 17242
rect 12034 17208 12090 17242
rect 12124 17208 12180 17242
rect 12214 17208 12270 17242
rect 12304 17208 12401 17242
rect 11439 17189 12401 17208
rect 11439 17148 11511 17189
rect 11439 17114 11458 17148
rect 11492 17114 11511 17148
rect 12329 17129 12401 17189
rect 11439 17058 11511 17114
rect 11439 17024 11458 17058
rect 11492 17024 11511 17058
rect 11439 16968 11511 17024
rect 11439 16934 11458 16968
rect 11492 16934 11511 16968
rect 11439 16878 11511 16934
rect 11439 16844 11458 16878
rect 11492 16844 11511 16878
rect 11439 16788 11511 16844
rect 11439 16754 11458 16788
rect 11492 16754 11511 16788
rect 11439 16698 11511 16754
rect 11439 16664 11458 16698
rect 11492 16664 11511 16698
rect 11439 16608 11511 16664
rect 11439 16574 11458 16608
rect 11492 16574 11511 16608
rect 11439 16518 11511 16574
rect 11439 16484 11458 16518
rect 11492 16484 11511 16518
rect 11439 16428 11511 16484
rect 11573 17066 12267 17127
rect 11573 17032 11632 17066
rect 11666 17054 11722 17066
rect 11694 17032 11722 17054
rect 11756 17054 11812 17066
rect 11756 17032 11760 17054
rect 11573 17020 11660 17032
rect 11694 17020 11760 17032
rect 11794 17032 11812 17054
rect 11846 17054 11902 17066
rect 11846 17032 11860 17054
rect 11794 17020 11860 17032
rect 11894 17032 11902 17054
rect 11936 17054 11992 17066
rect 12026 17054 12082 17066
rect 12116 17054 12172 17066
rect 11936 17032 11960 17054
rect 12026 17032 12060 17054
rect 12116 17032 12160 17054
rect 12206 17032 12267 17066
rect 11894 17020 11960 17032
rect 11994 17020 12060 17032
rect 12094 17020 12160 17032
rect 12194 17020 12267 17032
rect 11573 16976 12267 17020
rect 11573 16942 11632 16976
rect 11666 16954 11722 16976
rect 11694 16942 11722 16954
rect 11756 16954 11812 16976
rect 11756 16942 11760 16954
rect 11573 16920 11660 16942
rect 11694 16920 11760 16942
rect 11794 16942 11812 16954
rect 11846 16954 11902 16976
rect 11846 16942 11860 16954
rect 11794 16920 11860 16942
rect 11894 16942 11902 16954
rect 11936 16954 11992 16976
rect 12026 16954 12082 16976
rect 12116 16954 12172 16976
rect 11936 16942 11960 16954
rect 12026 16942 12060 16954
rect 12116 16942 12160 16954
rect 12206 16942 12267 16976
rect 11894 16920 11960 16942
rect 11994 16920 12060 16942
rect 12094 16920 12160 16942
rect 12194 16920 12267 16942
rect 11573 16886 12267 16920
rect 11573 16852 11632 16886
rect 11666 16854 11722 16886
rect 11694 16852 11722 16854
rect 11756 16854 11812 16886
rect 11756 16852 11760 16854
rect 11573 16820 11660 16852
rect 11694 16820 11760 16852
rect 11794 16852 11812 16854
rect 11846 16854 11902 16886
rect 11846 16852 11860 16854
rect 11794 16820 11860 16852
rect 11894 16852 11902 16854
rect 11936 16854 11992 16886
rect 12026 16854 12082 16886
rect 12116 16854 12172 16886
rect 11936 16852 11960 16854
rect 12026 16852 12060 16854
rect 12116 16852 12160 16854
rect 12206 16852 12267 16886
rect 11894 16820 11960 16852
rect 11994 16820 12060 16852
rect 12094 16820 12160 16852
rect 12194 16820 12267 16852
rect 11573 16796 12267 16820
rect 11573 16762 11632 16796
rect 11666 16762 11722 16796
rect 11756 16762 11812 16796
rect 11846 16762 11902 16796
rect 11936 16762 11992 16796
rect 12026 16762 12082 16796
rect 12116 16762 12172 16796
rect 12206 16762 12267 16796
rect 11573 16754 12267 16762
rect 11573 16720 11660 16754
rect 11694 16720 11760 16754
rect 11794 16720 11860 16754
rect 11894 16720 11960 16754
rect 11994 16720 12060 16754
rect 12094 16720 12160 16754
rect 12194 16720 12267 16754
rect 11573 16706 12267 16720
rect 11573 16672 11632 16706
rect 11666 16672 11722 16706
rect 11756 16672 11812 16706
rect 11846 16672 11902 16706
rect 11936 16672 11992 16706
rect 12026 16672 12082 16706
rect 12116 16672 12172 16706
rect 12206 16672 12267 16706
rect 11573 16654 12267 16672
rect 11573 16620 11660 16654
rect 11694 16620 11760 16654
rect 11794 16620 11860 16654
rect 11894 16620 11960 16654
rect 11994 16620 12060 16654
rect 12094 16620 12160 16654
rect 12194 16620 12267 16654
rect 11573 16616 12267 16620
rect 11573 16582 11632 16616
rect 11666 16582 11722 16616
rect 11756 16582 11812 16616
rect 11846 16582 11902 16616
rect 11936 16582 11992 16616
rect 12026 16582 12082 16616
rect 12116 16582 12172 16616
rect 12206 16582 12267 16616
rect 11573 16554 12267 16582
rect 11573 16526 11660 16554
rect 11694 16526 11760 16554
rect 11573 16492 11632 16526
rect 11694 16520 11722 16526
rect 11666 16492 11722 16520
rect 11756 16520 11760 16526
rect 11794 16526 11860 16554
rect 11794 16520 11812 16526
rect 11756 16492 11812 16520
rect 11846 16520 11860 16526
rect 11894 16526 11960 16554
rect 11994 16526 12060 16554
rect 12094 16526 12160 16554
rect 12194 16526 12267 16554
rect 11894 16520 11902 16526
rect 11846 16492 11902 16520
rect 11936 16520 11960 16526
rect 12026 16520 12060 16526
rect 12116 16520 12160 16526
rect 11936 16492 11992 16520
rect 12026 16492 12082 16520
rect 12116 16492 12172 16520
rect 12206 16492 12267 16526
rect 11573 16433 12267 16492
rect 12329 17095 12348 17129
rect 12382 17095 12401 17129
rect 12329 17039 12401 17095
rect 12329 17005 12348 17039
rect 12382 17005 12401 17039
rect 12329 16949 12401 17005
rect 12329 16915 12348 16949
rect 12382 16915 12401 16949
rect 12329 16859 12401 16915
rect 12329 16825 12348 16859
rect 12382 16825 12401 16859
rect 12329 16769 12401 16825
rect 12329 16735 12348 16769
rect 12382 16735 12401 16769
rect 12329 16679 12401 16735
rect 12329 16645 12348 16679
rect 12382 16645 12401 16679
rect 12329 16589 12401 16645
rect 12329 16555 12348 16589
rect 12382 16555 12401 16589
rect 12329 16499 12401 16555
rect 12329 16465 12348 16499
rect 12382 16465 12401 16499
rect 11439 16394 11458 16428
rect 11492 16394 11511 16428
rect 11439 16380 11511 16394
rect 12329 16409 12401 16465
rect 12329 16380 12348 16409
rect 11343 16375 12348 16380
rect 12382 16380 12401 16409
rect 12465 17218 12735 17274
rect 13825 17308 14095 17325
rect 13825 17274 13856 17308
rect 13890 17274 14029 17308
rect 14063 17274 14095 17308
rect 12465 17184 12496 17218
rect 12530 17184 12669 17218
rect 12703 17184 12735 17218
rect 12465 17128 12735 17184
rect 12465 17094 12496 17128
rect 12530 17094 12669 17128
rect 12703 17094 12735 17128
rect 12465 17038 12735 17094
rect 12465 17004 12496 17038
rect 12530 17004 12669 17038
rect 12703 17004 12735 17038
rect 12465 16948 12735 17004
rect 12465 16914 12496 16948
rect 12530 16914 12669 16948
rect 12703 16914 12735 16948
rect 12465 16858 12735 16914
rect 12465 16824 12496 16858
rect 12530 16824 12669 16858
rect 12703 16824 12735 16858
rect 12465 16768 12735 16824
rect 12465 16734 12496 16768
rect 12530 16734 12669 16768
rect 12703 16734 12735 16768
rect 12465 16678 12735 16734
rect 12465 16644 12496 16678
rect 12530 16644 12669 16678
rect 12703 16644 12735 16678
rect 12465 16588 12735 16644
rect 12465 16554 12496 16588
rect 12530 16554 12669 16588
rect 12703 16554 12735 16588
rect 12465 16498 12735 16554
rect 12465 16464 12496 16498
rect 12530 16464 12669 16498
rect 12703 16464 12735 16498
rect 12465 16408 12735 16464
rect 12465 16380 12496 16408
rect 12382 16375 12496 16380
rect 11343 16374 12496 16375
rect 12530 16374 12669 16408
rect 12703 16380 12735 16408
rect 12799 17242 13761 17261
rect 12799 17208 12910 17242
rect 12944 17208 13000 17242
rect 13034 17208 13090 17242
rect 13124 17208 13180 17242
rect 13214 17208 13270 17242
rect 13304 17208 13360 17242
rect 13394 17208 13450 17242
rect 13484 17208 13540 17242
rect 13574 17208 13630 17242
rect 13664 17208 13761 17242
rect 12799 17189 13761 17208
rect 12799 17148 12871 17189
rect 12799 17114 12818 17148
rect 12852 17114 12871 17148
rect 13689 17129 13761 17189
rect 12799 17058 12871 17114
rect 12799 17024 12818 17058
rect 12852 17024 12871 17058
rect 12799 16968 12871 17024
rect 12799 16934 12818 16968
rect 12852 16934 12871 16968
rect 12799 16878 12871 16934
rect 12799 16844 12818 16878
rect 12852 16844 12871 16878
rect 12799 16788 12871 16844
rect 12799 16754 12818 16788
rect 12852 16754 12871 16788
rect 12799 16698 12871 16754
rect 12799 16664 12818 16698
rect 12852 16664 12871 16698
rect 12799 16608 12871 16664
rect 12799 16574 12818 16608
rect 12852 16574 12871 16608
rect 12799 16518 12871 16574
rect 12799 16484 12818 16518
rect 12852 16484 12871 16518
rect 12799 16428 12871 16484
rect 12933 17066 13627 17127
rect 12933 17032 12992 17066
rect 13026 17054 13082 17066
rect 13054 17032 13082 17054
rect 13116 17054 13172 17066
rect 13116 17032 13120 17054
rect 12933 17020 13020 17032
rect 13054 17020 13120 17032
rect 13154 17032 13172 17054
rect 13206 17054 13262 17066
rect 13206 17032 13220 17054
rect 13154 17020 13220 17032
rect 13254 17032 13262 17054
rect 13296 17054 13352 17066
rect 13386 17054 13442 17066
rect 13476 17054 13532 17066
rect 13296 17032 13320 17054
rect 13386 17032 13420 17054
rect 13476 17032 13520 17054
rect 13566 17032 13627 17066
rect 13254 17020 13320 17032
rect 13354 17020 13420 17032
rect 13454 17020 13520 17032
rect 13554 17020 13627 17032
rect 12933 16976 13627 17020
rect 12933 16942 12992 16976
rect 13026 16954 13082 16976
rect 13054 16942 13082 16954
rect 13116 16954 13172 16976
rect 13116 16942 13120 16954
rect 12933 16920 13020 16942
rect 13054 16920 13120 16942
rect 13154 16942 13172 16954
rect 13206 16954 13262 16976
rect 13206 16942 13220 16954
rect 13154 16920 13220 16942
rect 13254 16942 13262 16954
rect 13296 16954 13352 16976
rect 13386 16954 13442 16976
rect 13476 16954 13532 16976
rect 13296 16942 13320 16954
rect 13386 16942 13420 16954
rect 13476 16942 13520 16954
rect 13566 16942 13627 16976
rect 13254 16920 13320 16942
rect 13354 16920 13420 16942
rect 13454 16920 13520 16942
rect 13554 16920 13627 16942
rect 12933 16886 13627 16920
rect 12933 16852 12992 16886
rect 13026 16854 13082 16886
rect 13054 16852 13082 16854
rect 13116 16854 13172 16886
rect 13116 16852 13120 16854
rect 12933 16820 13020 16852
rect 13054 16820 13120 16852
rect 13154 16852 13172 16854
rect 13206 16854 13262 16886
rect 13206 16852 13220 16854
rect 13154 16820 13220 16852
rect 13254 16852 13262 16854
rect 13296 16854 13352 16886
rect 13386 16854 13442 16886
rect 13476 16854 13532 16886
rect 13296 16852 13320 16854
rect 13386 16852 13420 16854
rect 13476 16852 13520 16854
rect 13566 16852 13627 16886
rect 13254 16820 13320 16852
rect 13354 16820 13420 16852
rect 13454 16820 13520 16852
rect 13554 16820 13627 16852
rect 12933 16796 13627 16820
rect 12933 16762 12992 16796
rect 13026 16762 13082 16796
rect 13116 16762 13172 16796
rect 13206 16762 13262 16796
rect 13296 16762 13352 16796
rect 13386 16762 13442 16796
rect 13476 16762 13532 16796
rect 13566 16762 13627 16796
rect 12933 16754 13627 16762
rect 12933 16720 13020 16754
rect 13054 16720 13120 16754
rect 13154 16720 13220 16754
rect 13254 16720 13320 16754
rect 13354 16720 13420 16754
rect 13454 16720 13520 16754
rect 13554 16720 13627 16754
rect 12933 16706 13627 16720
rect 12933 16672 12992 16706
rect 13026 16672 13082 16706
rect 13116 16672 13172 16706
rect 13206 16672 13262 16706
rect 13296 16672 13352 16706
rect 13386 16672 13442 16706
rect 13476 16672 13532 16706
rect 13566 16672 13627 16706
rect 12933 16654 13627 16672
rect 12933 16620 13020 16654
rect 13054 16620 13120 16654
rect 13154 16620 13220 16654
rect 13254 16620 13320 16654
rect 13354 16620 13420 16654
rect 13454 16620 13520 16654
rect 13554 16620 13627 16654
rect 12933 16616 13627 16620
rect 12933 16582 12992 16616
rect 13026 16582 13082 16616
rect 13116 16582 13172 16616
rect 13206 16582 13262 16616
rect 13296 16582 13352 16616
rect 13386 16582 13442 16616
rect 13476 16582 13532 16616
rect 13566 16582 13627 16616
rect 12933 16554 13627 16582
rect 12933 16526 13020 16554
rect 13054 16526 13120 16554
rect 12933 16492 12992 16526
rect 13054 16520 13082 16526
rect 13026 16492 13082 16520
rect 13116 16520 13120 16526
rect 13154 16526 13220 16554
rect 13154 16520 13172 16526
rect 13116 16492 13172 16520
rect 13206 16520 13220 16526
rect 13254 16526 13320 16554
rect 13354 16526 13420 16554
rect 13454 16526 13520 16554
rect 13554 16526 13627 16554
rect 13254 16520 13262 16526
rect 13206 16492 13262 16520
rect 13296 16520 13320 16526
rect 13386 16520 13420 16526
rect 13476 16520 13520 16526
rect 13296 16492 13352 16520
rect 13386 16492 13442 16520
rect 13476 16492 13532 16520
rect 13566 16492 13627 16526
rect 12933 16433 13627 16492
rect 13689 17095 13708 17129
rect 13742 17095 13761 17129
rect 13689 17039 13761 17095
rect 13689 17005 13708 17039
rect 13742 17005 13761 17039
rect 13689 16949 13761 17005
rect 13689 16915 13708 16949
rect 13742 16915 13761 16949
rect 13689 16859 13761 16915
rect 13689 16825 13708 16859
rect 13742 16825 13761 16859
rect 13689 16769 13761 16825
rect 13689 16735 13708 16769
rect 13742 16735 13761 16769
rect 13689 16679 13761 16735
rect 13689 16645 13708 16679
rect 13742 16645 13761 16679
rect 13689 16589 13761 16645
rect 13689 16555 13708 16589
rect 13742 16555 13761 16589
rect 13689 16499 13761 16555
rect 13689 16465 13708 16499
rect 13742 16465 13761 16499
rect 12799 16394 12818 16428
rect 12852 16394 12871 16428
rect 12799 16380 12871 16394
rect 13689 16409 13761 16465
rect 13689 16380 13708 16409
rect 12703 16375 13708 16380
rect 13742 16380 13761 16409
rect 13825 17218 14095 17274
rect 15185 17308 15284 17325
rect 15185 17274 15216 17308
rect 15250 17274 15284 17308
rect 13825 17184 13856 17218
rect 13890 17184 14029 17218
rect 14063 17184 14095 17218
rect 13825 17128 14095 17184
rect 13825 17094 13856 17128
rect 13890 17094 14029 17128
rect 14063 17094 14095 17128
rect 13825 17038 14095 17094
rect 13825 17004 13856 17038
rect 13890 17004 14029 17038
rect 14063 17004 14095 17038
rect 13825 16948 14095 17004
rect 13825 16914 13856 16948
rect 13890 16914 14029 16948
rect 14063 16914 14095 16948
rect 13825 16858 14095 16914
rect 13825 16824 13856 16858
rect 13890 16824 14029 16858
rect 14063 16824 14095 16858
rect 13825 16768 14095 16824
rect 13825 16734 13856 16768
rect 13890 16734 14029 16768
rect 14063 16734 14095 16768
rect 13825 16678 14095 16734
rect 13825 16644 13856 16678
rect 13890 16644 14029 16678
rect 14063 16644 14095 16678
rect 13825 16588 14095 16644
rect 13825 16554 13856 16588
rect 13890 16554 14029 16588
rect 14063 16554 14095 16588
rect 13825 16498 14095 16554
rect 13825 16464 13856 16498
rect 13890 16464 14029 16498
rect 14063 16464 14095 16498
rect 13825 16408 14095 16464
rect 13825 16380 13856 16408
rect 13742 16375 13856 16380
rect 12703 16374 13856 16375
rect 13890 16374 14029 16408
rect 14063 16380 14095 16408
rect 14159 17242 15121 17261
rect 14159 17208 14270 17242
rect 14304 17208 14360 17242
rect 14394 17208 14450 17242
rect 14484 17208 14540 17242
rect 14574 17208 14630 17242
rect 14664 17208 14720 17242
rect 14754 17208 14810 17242
rect 14844 17208 14900 17242
rect 14934 17208 14990 17242
rect 15024 17208 15121 17242
rect 14159 17189 15121 17208
rect 14159 17148 14231 17189
rect 14159 17114 14178 17148
rect 14212 17114 14231 17148
rect 15049 17129 15121 17189
rect 14159 17058 14231 17114
rect 14159 17024 14178 17058
rect 14212 17024 14231 17058
rect 14159 16968 14231 17024
rect 14159 16934 14178 16968
rect 14212 16934 14231 16968
rect 14159 16878 14231 16934
rect 14159 16844 14178 16878
rect 14212 16844 14231 16878
rect 14159 16788 14231 16844
rect 14159 16754 14178 16788
rect 14212 16754 14231 16788
rect 14159 16698 14231 16754
rect 14159 16664 14178 16698
rect 14212 16664 14231 16698
rect 14159 16608 14231 16664
rect 14159 16574 14178 16608
rect 14212 16574 14231 16608
rect 14159 16518 14231 16574
rect 14159 16484 14178 16518
rect 14212 16484 14231 16518
rect 14159 16428 14231 16484
rect 14293 17066 14987 17127
rect 14293 17032 14352 17066
rect 14386 17054 14442 17066
rect 14414 17032 14442 17054
rect 14476 17054 14532 17066
rect 14476 17032 14480 17054
rect 14293 17020 14380 17032
rect 14414 17020 14480 17032
rect 14514 17032 14532 17054
rect 14566 17054 14622 17066
rect 14566 17032 14580 17054
rect 14514 17020 14580 17032
rect 14614 17032 14622 17054
rect 14656 17054 14712 17066
rect 14746 17054 14802 17066
rect 14836 17054 14892 17066
rect 14656 17032 14680 17054
rect 14746 17032 14780 17054
rect 14836 17032 14880 17054
rect 14926 17032 14987 17066
rect 14614 17020 14680 17032
rect 14714 17020 14780 17032
rect 14814 17020 14880 17032
rect 14914 17020 14987 17032
rect 14293 16976 14987 17020
rect 14293 16942 14352 16976
rect 14386 16954 14442 16976
rect 14414 16942 14442 16954
rect 14476 16954 14532 16976
rect 14476 16942 14480 16954
rect 14293 16920 14380 16942
rect 14414 16920 14480 16942
rect 14514 16942 14532 16954
rect 14566 16954 14622 16976
rect 14566 16942 14580 16954
rect 14514 16920 14580 16942
rect 14614 16942 14622 16954
rect 14656 16954 14712 16976
rect 14746 16954 14802 16976
rect 14836 16954 14892 16976
rect 14656 16942 14680 16954
rect 14746 16942 14780 16954
rect 14836 16942 14880 16954
rect 14926 16942 14987 16976
rect 14614 16920 14680 16942
rect 14714 16920 14780 16942
rect 14814 16920 14880 16942
rect 14914 16920 14987 16942
rect 14293 16886 14987 16920
rect 14293 16852 14352 16886
rect 14386 16854 14442 16886
rect 14414 16852 14442 16854
rect 14476 16854 14532 16886
rect 14476 16852 14480 16854
rect 14293 16820 14380 16852
rect 14414 16820 14480 16852
rect 14514 16852 14532 16854
rect 14566 16854 14622 16886
rect 14566 16852 14580 16854
rect 14514 16820 14580 16852
rect 14614 16852 14622 16854
rect 14656 16854 14712 16886
rect 14746 16854 14802 16886
rect 14836 16854 14892 16886
rect 14656 16852 14680 16854
rect 14746 16852 14780 16854
rect 14836 16852 14880 16854
rect 14926 16852 14987 16886
rect 14614 16820 14680 16852
rect 14714 16820 14780 16852
rect 14814 16820 14880 16852
rect 14914 16820 14987 16852
rect 14293 16796 14987 16820
rect 14293 16762 14352 16796
rect 14386 16762 14442 16796
rect 14476 16762 14532 16796
rect 14566 16762 14622 16796
rect 14656 16762 14712 16796
rect 14746 16762 14802 16796
rect 14836 16762 14892 16796
rect 14926 16762 14987 16796
rect 14293 16754 14987 16762
rect 14293 16720 14380 16754
rect 14414 16720 14480 16754
rect 14514 16720 14580 16754
rect 14614 16720 14680 16754
rect 14714 16720 14780 16754
rect 14814 16720 14880 16754
rect 14914 16720 14987 16754
rect 14293 16706 14987 16720
rect 14293 16672 14352 16706
rect 14386 16672 14442 16706
rect 14476 16672 14532 16706
rect 14566 16672 14622 16706
rect 14656 16672 14712 16706
rect 14746 16672 14802 16706
rect 14836 16672 14892 16706
rect 14926 16672 14987 16706
rect 14293 16654 14987 16672
rect 14293 16620 14380 16654
rect 14414 16620 14480 16654
rect 14514 16620 14580 16654
rect 14614 16620 14680 16654
rect 14714 16620 14780 16654
rect 14814 16620 14880 16654
rect 14914 16620 14987 16654
rect 14293 16616 14987 16620
rect 14293 16582 14352 16616
rect 14386 16582 14442 16616
rect 14476 16582 14532 16616
rect 14566 16582 14622 16616
rect 14656 16582 14712 16616
rect 14746 16582 14802 16616
rect 14836 16582 14892 16616
rect 14926 16582 14987 16616
rect 14293 16554 14987 16582
rect 14293 16526 14380 16554
rect 14414 16526 14480 16554
rect 14293 16492 14352 16526
rect 14414 16520 14442 16526
rect 14386 16492 14442 16520
rect 14476 16520 14480 16526
rect 14514 16526 14580 16554
rect 14514 16520 14532 16526
rect 14476 16492 14532 16520
rect 14566 16520 14580 16526
rect 14614 16526 14680 16554
rect 14714 16526 14780 16554
rect 14814 16526 14880 16554
rect 14914 16526 14987 16554
rect 14614 16520 14622 16526
rect 14566 16492 14622 16520
rect 14656 16520 14680 16526
rect 14746 16520 14780 16526
rect 14836 16520 14880 16526
rect 14656 16492 14712 16520
rect 14746 16492 14802 16520
rect 14836 16492 14892 16520
rect 14926 16492 14987 16526
rect 14293 16433 14987 16492
rect 15049 17095 15068 17129
rect 15102 17095 15121 17129
rect 15049 17039 15121 17095
rect 15049 17005 15068 17039
rect 15102 17005 15121 17039
rect 15049 16949 15121 17005
rect 15049 16915 15068 16949
rect 15102 16915 15121 16949
rect 15049 16859 15121 16915
rect 15049 16825 15068 16859
rect 15102 16825 15121 16859
rect 15049 16769 15121 16825
rect 15049 16735 15068 16769
rect 15102 16735 15121 16769
rect 15049 16679 15121 16735
rect 15049 16645 15068 16679
rect 15102 16645 15121 16679
rect 15049 16589 15121 16645
rect 15049 16555 15068 16589
rect 15102 16555 15121 16589
rect 15049 16499 15121 16555
rect 15049 16465 15068 16499
rect 15102 16465 15121 16499
rect 14159 16394 14178 16428
rect 14212 16394 14231 16428
rect 14159 16380 14231 16394
rect 15049 16409 15121 16465
rect 15049 16380 15068 16409
rect 14063 16375 15068 16380
rect 15102 16380 15121 16409
rect 15185 17218 15284 17274
rect 15185 17184 15216 17218
rect 15250 17184 15284 17218
rect 15185 17128 15284 17184
rect 15185 17094 15216 17128
rect 15250 17094 15284 17128
rect 15185 17038 15284 17094
rect 15185 17004 15216 17038
rect 15250 17004 15284 17038
rect 15185 16948 15284 17004
rect 15185 16914 15216 16948
rect 15250 16914 15284 16948
rect 15185 16858 15284 16914
rect 15185 16824 15216 16858
rect 15250 16824 15284 16858
rect 15185 16768 15284 16824
rect 15185 16734 15216 16768
rect 15250 16734 15284 16768
rect 15185 16678 15284 16734
rect 15185 16644 15216 16678
rect 15250 16644 15284 16678
rect 15185 16588 15284 16644
rect 15185 16554 15216 16588
rect 15250 16554 15284 16588
rect 15185 16498 15284 16554
rect 15185 16464 15216 16498
rect 15250 16464 15284 16498
rect 15185 16408 15284 16464
rect 15185 16380 15216 16408
rect 15102 16375 15216 16380
rect 14063 16374 15216 16375
rect 15250 16380 15284 16408
rect 15250 16374 15290 16380
rect 11270 16352 15290 16374
rect 11270 16318 11516 16352
rect 11550 16318 11606 16352
rect 11640 16318 11696 16352
rect 11730 16318 11786 16352
rect 11820 16318 11876 16352
rect 11910 16318 11966 16352
rect 12000 16318 12056 16352
rect 12090 16318 12146 16352
rect 12180 16318 12236 16352
rect 12270 16318 12876 16352
rect 12910 16318 12966 16352
rect 13000 16318 13056 16352
rect 13090 16318 13146 16352
rect 13180 16318 13236 16352
rect 13270 16318 13326 16352
rect 13360 16318 13416 16352
rect 13450 16318 13506 16352
rect 13540 16318 13596 16352
rect 13630 16318 14236 16352
rect 14270 16318 14326 16352
rect 14360 16318 14416 16352
rect 14450 16318 14506 16352
rect 14540 16318 14596 16352
rect 14630 16318 14686 16352
rect 14720 16318 14776 16352
rect 14810 16318 14866 16352
rect 14900 16318 14956 16352
rect 14990 16318 15290 16352
rect 11270 16284 11309 16318
rect 11343 16284 12496 16318
rect 12530 16284 12669 16318
rect 12703 16284 13856 16318
rect 13890 16284 14029 16318
rect 14063 16284 15216 16318
rect 15250 16284 15290 16318
rect 11270 16228 15290 16284
rect 11270 16194 11309 16228
rect 11343 16205 12496 16228
rect 11343 16194 11410 16205
rect 11270 16171 11410 16194
rect 11444 16171 11500 16205
rect 11534 16171 11590 16205
rect 11624 16171 11680 16205
rect 11714 16171 11770 16205
rect 11804 16171 11860 16205
rect 11894 16171 11950 16205
rect 11984 16171 12040 16205
rect 12074 16171 12130 16205
rect 12164 16171 12220 16205
rect 12254 16171 12310 16205
rect 12344 16171 12400 16205
rect 12434 16194 12496 16205
rect 12530 16194 12669 16228
rect 12703 16205 13856 16228
rect 12703 16194 12770 16205
rect 12434 16171 12770 16194
rect 12804 16171 12860 16205
rect 12894 16171 12950 16205
rect 12984 16171 13040 16205
rect 13074 16171 13130 16205
rect 13164 16171 13220 16205
rect 13254 16171 13310 16205
rect 13344 16171 13400 16205
rect 13434 16171 13490 16205
rect 13524 16171 13580 16205
rect 13614 16171 13670 16205
rect 13704 16171 13760 16205
rect 13794 16194 13856 16205
rect 13890 16194 14029 16228
rect 14063 16205 15216 16228
rect 14063 16194 14130 16205
rect 13794 16171 14130 16194
rect 14164 16171 14220 16205
rect 14254 16171 14310 16205
rect 14344 16171 14400 16205
rect 14434 16171 14490 16205
rect 14524 16171 14580 16205
rect 14614 16171 14670 16205
rect 14704 16171 14760 16205
rect 14794 16171 14850 16205
rect 14884 16171 14940 16205
rect 14974 16171 15030 16205
rect 15064 16171 15120 16205
rect 15154 16194 15216 16205
rect 15250 16194 15290 16228
rect 15154 16171 15290 16194
rect 11270 16130 15290 16171
rect 16233 18501 16267 18563
rect 15483 16181 15517 16243
rect 16596 18560 16692 18594
rect 16952 18560 17048 18594
rect 16596 18498 16630 18560
rect 16780 18550 16860 18560
rect 17014 18498 17048 18560
rect 16596 17318 16630 17380
rect 17014 17318 17048 17380
rect 16596 17284 16692 17318
rect 16952 17284 17048 17318
rect 17383 18563 17479 18597
rect 17739 18563 17835 18597
rect 17383 18501 17417 18563
rect 17570 18550 17650 18563
rect 17801 18501 17835 18563
rect 17383 17111 17417 17173
rect 17801 17111 17835 17173
rect 17383 17077 17479 17111
rect 17739 17077 17835 17111
rect 16233 16181 16267 16243
rect 15483 16147 15579 16181
rect 16171 16147 16267 16181
rect 12560 16064 12640 16130
rect 13920 16064 14000 16130
rect 11276 16032 15284 16064
rect 11276 15998 11410 16032
rect 11444 15998 11500 16032
rect 11534 15998 11590 16032
rect 11624 15998 11680 16032
rect 11714 15998 11770 16032
rect 11804 15998 11860 16032
rect 11894 15998 11950 16032
rect 11984 15998 12040 16032
rect 12074 15998 12130 16032
rect 12164 15998 12220 16032
rect 12254 15998 12310 16032
rect 12344 15998 12400 16032
rect 12434 15998 12770 16032
rect 12804 15998 12860 16032
rect 12894 15998 12950 16032
rect 12984 15998 13040 16032
rect 13074 15998 13130 16032
rect 13164 15998 13220 16032
rect 13254 15998 13310 16032
rect 13344 15998 13400 16032
rect 13434 15998 13490 16032
rect 13524 15998 13580 16032
rect 13614 15998 13670 16032
rect 13704 15998 13760 16032
rect 13794 15998 14130 16032
rect 14164 15998 14220 16032
rect 14254 15998 14310 16032
rect 14344 15998 14400 16032
rect 14434 15998 14490 16032
rect 14524 15998 14580 16032
rect 14614 15998 14670 16032
rect 14704 15998 14760 16032
rect 14794 15998 14850 16032
rect 14884 15998 14940 16032
rect 14974 15998 15030 16032
rect 15064 15998 15120 16032
rect 15154 15998 15284 16032
rect 11276 15965 15284 15998
rect 11276 15948 11375 15965
rect 11276 15914 11309 15948
rect 11343 15914 11375 15948
rect 11276 15858 11375 15914
rect 12465 15948 12735 15965
rect 12465 15914 12496 15948
rect 12530 15914 12669 15948
rect 12703 15914 12735 15948
rect 11276 15824 11309 15858
rect 11343 15824 11375 15858
rect 11276 15768 11375 15824
rect 11276 15734 11309 15768
rect 11343 15734 11375 15768
rect 11276 15678 11375 15734
rect 11276 15644 11309 15678
rect 11343 15644 11375 15678
rect 11276 15588 11375 15644
rect 11276 15554 11309 15588
rect 11343 15554 11375 15588
rect 11276 15498 11375 15554
rect 11276 15464 11309 15498
rect 11343 15464 11375 15498
rect 11276 15408 11375 15464
rect 11276 15374 11309 15408
rect 11343 15374 11375 15408
rect 11276 15318 11375 15374
rect 11276 15284 11309 15318
rect 11343 15284 11375 15318
rect 11276 15228 11375 15284
rect 11276 15194 11309 15228
rect 11343 15194 11375 15228
rect 11276 15138 11375 15194
rect 11276 15104 11309 15138
rect 11343 15104 11375 15138
rect 11276 15048 11375 15104
rect 11276 15020 11309 15048
rect 11270 15014 11309 15020
rect 11343 15020 11375 15048
rect 11439 15882 12401 15901
rect 11439 15848 11550 15882
rect 11584 15848 11640 15882
rect 11674 15848 11730 15882
rect 11764 15848 11820 15882
rect 11854 15848 11910 15882
rect 11944 15848 12000 15882
rect 12034 15848 12090 15882
rect 12124 15848 12180 15882
rect 12214 15848 12270 15882
rect 12304 15848 12401 15882
rect 11439 15829 12401 15848
rect 11439 15788 11511 15829
rect 11439 15754 11458 15788
rect 11492 15754 11511 15788
rect 12329 15769 12401 15829
rect 11439 15698 11511 15754
rect 11439 15664 11458 15698
rect 11492 15664 11511 15698
rect 11439 15608 11511 15664
rect 11439 15574 11458 15608
rect 11492 15574 11511 15608
rect 11439 15518 11511 15574
rect 11439 15484 11458 15518
rect 11492 15484 11511 15518
rect 11439 15428 11511 15484
rect 11439 15394 11458 15428
rect 11492 15394 11511 15428
rect 11439 15338 11511 15394
rect 11439 15304 11458 15338
rect 11492 15304 11511 15338
rect 11439 15248 11511 15304
rect 11439 15214 11458 15248
rect 11492 15214 11511 15248
rect 11439 15158 11511 15214
rect 11439 15124 11458 15158
rect 11492 15124 11511 15158
rect 11439 15068 11511 15124
rect 11573 15706 12267 15767
rect 11573 15672 11632 15706
rect 11666 15694 11722 15706
rect 11694 15672 11722 15694
rect 11756 15694 11812 15706
rect 11756 15672 11760 15694
rect 11573 15660 11660 15672
rect 11694 15660 11760 15672
rect 11794 15672 11812 15694
rect 11846 15694 11902 15706
rect 11846 15672 11860 15694
rect 11794 15660 11860 15672
rect 11894 15672 11902 15694
rect 11936 15694 11992 15706
rect 12026 15694 12082 15706
rect 12116 15694 12172 15706
rect 11936 15672 11960 15694
rect 12026 15672 12060 15694
rect 12116 15672 12160 15694
rect 12206 15672 12267 15706
rect 11894 15660 11960 15672
rect 11994 15660 12060 15672
rect 12094 15660 12160 15672
rect 12194 15660 12267 15672
rect 11573 15616 12267 15660
rect 11573 15582 11632 15616
rect 11666 15594 11722 15616
rect 11694 15582 11722 15594
rect 11756 15594 11812 15616
rect 11756 15582 11760 15594
rect 11573 15560 11660 15582
rect 11694 15560 11760 15582
rect 11794 15582 11812 15594
rect 11846 15594 11902 15616
rect 11846 15582 11860 15594
rect 11794 15560 11860 15582
rect 11894 15582 11902 15594
rect 11936 15594 11992 15616
rect 12026 15594 12082 15616
rect 12116 15594 12172 15616
rect 11936 15582 11960 15594
rect 12026 15582 12060 15594
rect 12116 15582 12160 15594
rect 12206 15582 12267 15616
rect 11894 15560 11960 15582
rect 11994 15560 12060 15582
rect 12094 15560 12160 15582
rect 12194 15560 12267 15582
rect 11573 15526 12267 15560
rect 11573 15492 11632 15526
rect 11666 15494 11722 15526
rect 11694 15492 11722 15494
rect 11756 15494 11812 15526
rect 11756 15492 11760 15494
rect 11573 15460 11660 15492
rect 11694 15460 11760 15492
rect 11794 15492 11812 15494
rect 11846 15494 11902 15526
rect 11846 15492 11860 15494
rect 11794 15460 11860 15492
rect 11894 15492 11902 15494
rect 11936 15494 11992 15526
rect 12026 15494 12082 15526
rect 12116 15494 12172 15526
rect 11936 15492 11960 15494
rect 12026 15492 12060 15494
rect 12116 15492 12160 15494
rect 12206 15492 12267 15526
rect 11894 15460 11960 15492
rect 11994 15460 12060 15492
rect 12094 15460 12160 15492
rect 12194 15460 12267 15492
rect 11573 15436 12267 15460
rect 11573 15402 11632 15436
rect 11666 15402 11722 15436
rect 11756 15402 11812 15436
rect 11846 15402 11902 15436
rect 11936 15402 11992 15436
rect 12026 15402 12082 15436
rect 12116 15402 12172 15436
rect 12206 15402 12267 15436
rect 11573 15394 12267 15402
rect 11573 15360 11660 15394
rect 11694 15360 11760 15394
rect 11794 15360 11860 15394
rect 11894 15360 11960 15394
rect 11994 15360 12060 15394
rect 12094 15360 12160 15394
rect 12194 15360 12267 15394
rect 11573 15346 12267 15360
rect 11573 15312 11632 15346
rect 11666 15312 11722 15346
rect 11756 15312 11812 15346
rect 11846 15312 11902 15346
rect 11936 15312 11992 15346
rect 12026 15312 12082 15346
rect 12116 15312 12172 15346
rect 12206 15312 12267 15346
rect 11573 15294 12267 15312
rect 11573 15260 11660 15294
rect 11694 15260 11760 15294
rect 11794 15260 11860 15294
rect 11894 15260 11960 15294
rect 11994 15260 12060 15294
rect 12094 15260 12160 15294
rect 12194 15260 12267 15294
rect 11573 15256 12267 15260
rect 11573 15222 11632 15256
rect 11666 15222 11722 15256
rect 11756 15222 11812 15256
rect 11846 15222 11902 15256
rect 11936 15222 11992 15256
rect 12026 15222 12082 15256
rect 12116 15222 12172 15256
rect 12206 15222 12267 15256
rect 11573 15194 12267 15222
rect 11573 15166 11660 15194
rect 11694 15166 11760 15194
rect 11573 15132 11632 15166
rect 11694 15160 11722 15166
rect 11666 15132 11722 15160
rect 11756 15160 11760 15166
rect 11794 15166 11860 15194
rect 11794 15160 11812 15166
rect 11756 15132 11812 15160
rect 11846 15160 11860 15166
rect 11894 15166 11960 15194
rect 11994 15166 12060 15194
rect 12094 15166 12160 15194
rect 12194 15166 12267 15194
rect 11894 15160 11902 15166
rect 11846 15132 11902 15160
rect 11936 15160 11960 15166
rect 12026 15160 12060 15166
rect 12116 15160 12160 15166
rect 11936 15132 11992 15160
rect 12026 15132 12082 15160
rect 12116 15132 12172 15160
rect 12206 15132 12267 15166
rect 11573 15073 12267 15132
rect 12329 15735 12348 15769
rect 12382 15735 12401 15769
rect 12329 15679 12401 15735
rect 12329 15645 12348 15679
rect 12382 15645 12401 15679
rect 12329 15589 12401 15645
rect 12329 15555 12348 15589
rect 12382 15555 12401 15589
rect 12329 15499 12401 15555
rect 12329 15465 12348 15499
rect 12382 15465 12401 15499
rect 12329 15409 12401 15465
rect 12329 15375 12348 15409
rect 12382 15375 12401 15409
rect 12329 15319 12401 15375
rect 12329 15285 12348 15319
rect 12382 15285 12401 15319
rect 12329 15229 12401 15285
rect 12329 15195 12348 15229
rect 12382 15195 12401 15229
rect 12329 15139 12401 15195
rect 12329 15105 12348 15139
rect 12382 15105 12401 15139
rect 11439 15034 11458 15068
rect 11492 15034 11511 15068
rect 11439 15020 11511 15034
rect 12329 15049 12401 15105
rect 12329 15020 12348 15049
rect 11343 15015 12348 15020
rect 12382 15020 12401 15049
rect 12465 15858 12735 15914
rect 13825 15948 14095 15965
rect 13825 15914 13856 15948
rect 13890 15914 14029 15948
rect 14063 15914 14095 15948
rect 12465 15824 12496 15858
rect 12530 15824 12669 15858
rect 12703 15824 12735 15858
rect 12465 15768 12735 15824
rect 12465 15734 12496 15768
rect 12530 15734 12669 15768
rect 12703 15734 12735 15768
rect 12465 15678 12735 15734
rect 12465 15644 12496 15678
rect 12530 15644 12669 15678
rect 12703 15644 12735 15678
rect 12465 15588 12735 15644
rect 12465 15554 12496 15588
rect 12530 15554 12669 15588
rect 12703 15554 12735 15588
rect 12465 15498 12735 15554
rect 12465 15464 12496 15498
rect 12530 15464 12669 15498
rect 12703 15464 12735 15498
rect 12465 15408 12735 15464
rect 12465 15374 12496 15408
rect 12530 15374 12669 15408
rect 12703 15374 12735 15408
rect 12465 15318 12735 15374
rect 12465 15284 12496 15318
rect 12530 15284 12669 15318
rect 12703 15284 12735 15318
rect 12465 15228 12735 15284
rect 12465 15194 12496 15228
rect 12530 15194 12669 15228
rect 12703 15194 12735 15228
rect 12465 15138 12735 15194
rect 12465 15104 12496 15138
rect 12530 15104 12669 15138
rect 12703 15104 12735 15138
rect 12465 15048 12735 15104
rect 12465 15020 12496 15048
rect 12382 15015 12496 15020
rect 11343 15014 12496 15015
rect 12530 15014 12669 15048
rect 12703 15020 12735 15048
rect 12799 15882 13761 15901
rect 12799 15848 12910 15882
rect 12944 15848 13000 15882
rect 13034 15848 13090 15882
rect 13124 15848 13180 15882
rect 13214 15848 13270 15882
rect 13304 15848 13360 15882
rect 13394 15848 13450 15882
rect 13484 15848 13540 15882
rect 13574 15848 13630 15882
rect 13664 15848 13761 15882
rect 12799 15829 13761 15848
rect 12799 15788 12871 15829
rect 12799 15754 12818 15788
rect 12852 15754 12871 15788
rect 13689 15769 13761 15829
rect 12799 15698 12871 15754
rect 12799 15664 12818 15698
rect 12852 15664 12871 15698
rect 12799 15608 12871 15664
rect 12799 15574 12818 15608
rect 12852 15574 12871 15608
rect 12799 15518 12871 15574
rect 12799 15484 12818 15518
rect 12852 15484 12871 15518
rect 12799 15428 12871 15484
rect 12799 15394 12818 15428
rect 12852 15394 12871 15428
rect 12799 15338 12871 15394
rect 12799 15304 12818 15338
rect 12852 15304 12871 15338
rect 12799 15248 12871 15304
rect 12799 15214 12818 15248
rect 12852 15214 12871 15248
rect 12799 15158 12871 15214
rect 12799 15124 12818 15158
rect 12852 15124 12871 15158
rect 12799 15068 12871 15124
rect 12933 15706 13627 15767
rect 12933 15672 12992 15706
rect 13026 15694 13082 15706
rect 13054 15672 13082 15694
rect 13116 15694 13172 15706
rect 13116 15672 13120 15694
rect 12933 15660 13020 15672
rect 13054 15660 13120 15672
rect 13154 15672 13172 15694
rect 13206 15694 13262 15706
rect 13206 15672 13220 15694
rect 13154 15660 13220 15672
rect 13254 15672 13262 15694
rect 13296 15694 13352 15706
rect 13386 15694 13442 15706
rect 13476 15694 13532 15706
rect 13296 15672 13320 15694
rect 13386 15672 13420 15694
rect 13476 15672 13520 15694
rect 13566 15672 13627 15706
rect 13254 15660 13320 15672
rect 13354 15660 13420 15672
rect 13454 15660 13520 15672
rect 13554 15660 13627 15672
rect 12933 15616 13627 15660
rect 12933 15582 12992 15616
rect 13026 15594 13082 15616
rect 13054 15582 13082 15594
rect 13116 15594 13172 15616
rect 13116 15582 13120 15594
rect 12933 15560 13020 15582
rect 13054 15560 13120 15582
rect 13154 15582 13172 15594
rect 13206 15594 13262 15616
rect 13206 15582 13220 15594
rect 13154 15560 13220 15582
rect 13254 15582 13262 15594
rect 13296 15594 13352 15616
rect 13386 15594 13442 15616
rect 13476 15594 13532 15616
rect 13296 15582 13320 15594
rect 13386 15582 13420 15594
rect 13476 15582 13520 15594
rect 13566 15582 13627 15616
rect 13254 15560 13320 15582
rect 13354 15560 13420 15582
rect 13454 15560 13520 15582
rect 13554 15560 13627 15582
rect 12933 15526 13627 15560
rect 12933 15492 12992 15526
rect 13026 15494 13082 15526
rect 13054 15492 13082 15494
rect 13116 15494 13172 15526
rect 13116 15492 13120 15494
rect 12933 15460 13020 15492
rect 13054 15460 13120 15492
rect 13154 15492 13172 15494
rect 13206 15494 13262 15526
rect 13206 15492 13220 15494
rect 13154 15460 13220 15492
rect 13254 15492 13262 15494
rect 13296 15494 13352 15526
rect 13386 15494 13442 15526
rect 13476 15494 13532 15526
rect 13296 15492 13320 15494
rect 13386 15492 13420 15494
rect 13476 15492 13520 15494
rect 13566 15492 13627 15526
rect 13254 15460 13320 15492
rect 13354 15460 13420 15492
rect 13454 15460 13520 15492
rect 13554 15460 13627 15492
rect 12933 15436 13627 15460
rect 12933 15402 12992 15436
rect 13026 15402 13082 15436
rect 13116 15402 13172 15436
rect 13206 15402 13262 15436
rect 13296 15402 13352 15436
rect 13386 15402 13442 15436
rect 13476 15402 13532 15436
rect 13566 15402 13627 15436
rect 12933 15394 13627 15402
rect 12933 15360 13020 15394
rect 13054 15360 13120 15394
rect 13154 15360 13220 15394
rect 13254 15360 13320 15394
rect 13354 15360 13420 15394
rect 13454 15360 13520 15394
rect 13554 15360 13627 15394
rect 12933 15346 13627 15360
rect 12933 15312 12992 15346
rect 13026 15312 13082 15346
rect 13116 15312 13172 15346
rect 13206 15312 13262 15346
rect 13296 15312 13352 15346
rect 13386 15312 13442 15346
rect 13476 15312 13532 15346
rect 13566 15312 13627 15346
rect 12933 15294 13627 15312
rect 12933 15260 13020 15294
rect 13054 15260 13120 15294
rect 13154 15260 13220 15294
rect 13254 15260 13320 15294
rect 13354 15260 13420 15294
rect 13454 15260 13520 15294
rect 13554 15260 13627 15294
rect 12933 15256 13627 15260
rect 12933 15222 12992 15256
rect 13026 15222 13082 15256
rect 13116 15222 13172 15256
rect 13206 15222 13262 15256
rect 13296 15222 13352 15256
rect 13386 15222 13442 15256
rect 13476 15222 13532 15256
rect 13566 15222 13627 15256
rect 12933 15194 13627 15222
rect 12933 15166 13020 15194
rect 13054 15166 13120 15194
rect 12933 15132 12992 15166
rect 13054 15160 13082 15166
rect 13026 15132 13082 15160
rect 13116 15160 13120 15166
rect 13154 15166 13220 15194
rect 13154 15160 13172 15166
rect 13116 15132 13172 15160
rect 13206 15160 13220 15166
rect 13254 15166 13320 15194
rect 13354 15166 13420 15194
rect 13454 15166 13520 15194
rect 13554 15166 13627 15194
rect 13254 15160 13262 15166
rect 13206 15132 13262 15160
rect 13296 15160 13320 15166
rect 13386 15160 13420 15166
rect 13476 15160 13520 15166
rect 13296 15132 13352 15160
rect 13386 15132 13442 15160
rect 13476 15132 13532 15160
rect 13566 15132 13627 15166
rect 12933 15073 13627 15132
rect 13689 15735 13708 15769
rect 13742 15735 13761 15769
rect 13689 15679 13761 15735
rect 13689 15645 13708 15679
rect 13742 15645 13761 15679
rect 13689 15589 13761 15645
rect 13689 15555 13708 15589
rect 13742 15555 13761 15589
rect 13689 15499 13761 15555
rect 13689 15465 13708 15499
rect 13742 15465 13761 15499
rect 13689 15409 13761 15465
rect 13689 15375 13708 15409
rect 13742 15375 13761 15409
rect 13689 15319 13761 15375
rect 13689 15285 13708 15319
rect 13742 15285 13761 15319
rect 13689 15229 13761 15285
rect 13689 15195 13708 15229
rect 13742 15195 13761 15229
rect 13689 15139 13761 15195
rect 13689 15105 13708 15139
rect 13742 15105 13761 15139
rect 12799 15034 12818 15068
rect 12852 15034 12871 15068
rect 12799 15020 12871 15034
rect 13689 15049 13761 15105
rect 13689 15020 13708 15049
rect 12703 15015 13708 15020
rect 13742 15020 13761 15049
rect 13825 15858 14095 15914
rect 15185 15948 15284 15965
rect 15185 15914 15216 15948
rect 15250 15914 15284 15948
rect 13825 15824 13856 15858
rect 13890 15824 14029 15858
rect 14063 15824 14095 15858
rect 13825 15768 14095 15824
rect 13825 15734 13856 15768
rect 13890 15734 14029 15768
rect 14063 15734 14095 15768
rect 13825 15678 14095 15734
rect 13825 15644 13856 15678
rect 13890 15644 14029 15678
rect 14063 15644 14095 15678
rect 13825 15588 14095 15644
rect 13825 15554 13856 15588
rect 13890 15554 14029 15588
rect 14063 15554 14095 15588
rect 13825 15498 14095 15554
rect 13825 15464 13856 15498
rect 13890 15464 14029 15498
rect 14063 15464 14095 15498
rect 13825 15408 14095 15464
rect 13825 15374 13856 15408
rect 13890 15374 14029 15408
rect 14063 15374 14095 15408
rect 13825 15318 14095 15374
rect 13825 15284 13856 15318
rect 13890 15284 14029 15318
rect 14063 15284 14095 15318
rect 13825 15228 14095 15284
rect 13825 15194 13856 15228
rect 13890 15194 14029 15228
rect 14063 15194 14095 15228
rect 13825 15138 14095 15194
rect 13825 15104 13856 15138
rect 13890 15104 14029 15138
rect 14063 15104 14095 15138
rect 13825 15048 14095 15104
rect 13825 15020 13856 15048
rect 13742 15015 13856 15020
rect 12703 15014 13856 15015
rect 13890 15014 14029 15048
rect 14063 15020 14095 15048
rect 14159 15882 15121 15901
rect 14159 15848 14270 15882
rect 14304 15848 14360 15882
rect 14394 15848 14450 15882
rect 14484 15848 14540 15882
rect 14574 15848 14630 15882
rect 14664 15848 14720 15882
rect 14754 15848 14810 15882
rect 14844 15848 14900 15882
rect 14934 15848 14990 15882
rect 15024 15848 15121 15882
rect 14159 15829 15121 15848
rect 14159 15788 14231 15829
rect 14159 15754 14178 15788
rect 14212 15754 14231 15788
rect 15049 15769 15121 15829
rect 14159 15698 14231 15754
rect 14159 15664 14178 15698
rect 14212 15664 14231 15698
rect 14159 15608 14231 15664
rect 14159 15574 14178 15608
rect 14212 15574 14231 15608
rect 14159 15518 14231 15574
rect 14159 15484 14178 15518
rect 14212 15484 14231 15518
rect 14159 15428 14231 15484
rect 14159 15394 14178 15428
rect 14212 15394 14231 15428
rect 14159 15338 14231 15394
rect 14159 15304 14178 15338
rect 14212 15304 14231 15338
rect 14159 15248 14231 15304
rect 14159 15214 14178 15248
rect 14212 15214 14231 15248
rect 14159 15158 14231 15214
rect 14159 15124 14178 15158
rect 14212 15124 14231 15158
rect 14159 15068 14231 15124
rect 14293 15706 14987 15767
rect 14293 15672 14352 15706
rect 14386 15694 14442 15706
rect 14414 15672 14442 15694
rect 14476 15694 14532 15706
rect 14476 15672 14480 15694
rect 14293 15660 14380 15672
rect 14414 15660 14480 15672
rect 14514 15672 14532 15694
rect 14566 15694 14622 15706
rect 14566 15672 14580 15694
rect 14514 15660 14580 15672
rect 14614 15672 14622 15694
rect 14656 15694 14712 15706
rect 14746 15694 14802 15706
rect 14836 15694 14892 15706
rect 14656 15672 14680 15694
rect 14746 15672 14780 15694
rect 14836 15672 14880 15694
rect 14926 15672 14987 15706
rect 14614 15660 14680 15672
rect 14714 15660 14780 15672
rect 14814 15660 14880 15672
rect 14914 15660 14987 15672
rect 14293 15616 14987 15660
rect 14293 15582 14352 15616
rect 14386 15594 14442 15616
rect 14414 15582 14442 15594
rect 14476 15594 14532 15616
rect 14476 15582 14480 15594
rect 14293 15560 14380 15582
rect 14414 15560 14480 15582
rect 14514 15582 14532 15594
rect 14566 15594 14622 15616
rect 14566 15582 14580 15594
rect 14514 15560 14580 15582
rect 14614 15582 14622 15594
rect 14656 15594 14712 15616
rect 14746 15594 14802 15616
rect 14836 15594 14892 15616
rect 14656 15582 14680 15594
rect 14746 15582 14780 15594
rect 14836 15582 14880 15594
rect 14926 15582 14987 15616
rect 14614 15560 14680 15582
rect 14714 15560 14780 15582
rect 14814 15560 14880 15582
rect 14914 15560 14987 15582
rect 14293 15526 14987 15560
rect 14293 15492 14352 15526
rect 14386 15494 14442 15526
rect 14414 15492 14442 15494
rect 14476 15494 14532 15526
rect 14476 15492 14480 15494
rect 14293 15460 14380 15492
rect 14414 15460 14480 15492
rect 14514 15492 14532 15494
rect 14566 15494 14622 15526
rect 14566 15492 14580 15494
rect 14514 15460 14580 15492
rect 14614 15492 14622 15494
rect 14656 15494 14712 15526
rect 14746 15494 14802 15526
rect 14836 15494 14892 15526
rect 14656 15492 14680 15494
rect 14746 15492 14780 15494
rect 14836 15492 14880 15494
rect 14926 15492 14987 15526
rect 14614 15460 14680 15492
rect 14714 15460 14780 15492
rect 14814 15460 14880 15492
rect 14914 15460 14987 15492
rect 14293 15436 14987 15460
rect 14293 15402 14352 15436
rect 14386 15402 14442 15436
rect 14476 15402 14532 15436
rect 14566 15402 14622 15436
rect 14656 15402 14712 15436
rect 14746 15402 14802 15436
rect 14836 15402 14892 15436
rect 14926 15402 14987 15436
rect 14293 15394 14987 15402
rect 14293 15360 14380 15394
rect 14414 15360 14480 15394
rect 14514 15360 14580 15394
rect 14614 15360 14680 15394
rect 14714 15360 14780 15394
rect 14814 15360 14880 15394
rect 14914 15360 14987 15394
rect 14293 15346 14987 15360
rect 14293 15312 14352 15346
rect 14386 15312 14442 15346
rect 14476 15312 14532 15346
rect 14566 15312 14622 15346
rect 14656 15312 14712 15346
rect 14746 15312 14802 15346
rect 14836 15312 14892 15346
rect 14926 15312 14987 15346
rect 14293 15294 14987 15312
rect 14293 15260 14380 15294
rect 14414 15260 14480 15294
rect 14514 15260 14580 15294
rect 14614 15260 14680 15294
rect 14714 15260 14780 15294
rect 14814 15260 14880 15294
rect 14914 15260 14987 15294
rect 14293 15256 14987 15260
rect 14293 15222 14352 15256
rect 14386 15222 14442 15256
rect 14476 15222 14532 15256
rect 14566 15222 14622 15256
rect 14656 15222 14712 15256
rect 14746 15222 14802 15256
rect 14836 15222 14892 15256
rect 14926 15222 14987 15256
rect 14293 15194 14987 15222
rect 14293 15166 14380 15194
rect 14414 15166 14480 15194
rect 14293 15132 14352 15166
rect 14414 15160 14442 15166
rect 14386 15132 14442 15160
rect 14476 15160 14480 15166
rect 14514 15166 14580 15194
rect 14514 15160 14532 15166
rect 14476 15132 14532 15160
rect 14566 15160 14580 15166
rect 14614 15166 14680 15194
rect 14714 15166 14780 15194
rect 14814 15166 14880 15194
rect 14914 15166 14987 15194
rect 14614 15160 14622 15166
rect 14566 15132 14622 15160
rect 14656 15160 14680 15166
rect 14746 15160 14780 15166
rect 14836 15160 14880 15166
rect 14656 15132 14712 15160
rect 14746 15132 14802 15160
rect 14836 15132 14892 15160
rect 14926 15132 14987 15166
rect 14293 15073 14987 15132
rect 15049 15735 15068 15769
rect 15102 15735 15121 15769
rect 15049 15679 15121 15735
rect 15049 15645 15068 15679
rect 15102 15645 15121 15679
rect 15049 15589 15121 15645
rect 15049 15555 15068 15589
rect 15102 15555 15121 15589
rect 15049 15499 15121 15555
rect 15049 15465 15068 15499
rect 15102 15465 15121 15499
rect 15049 15409 15121 15465
rect 15049 15375 15068 15409
rect 15102 15375 15121 15409
rect 15049 15319 15121 15375
rect 15049 15285 15068 15319
rect 15102 15285 15121 15319
rect 15049 15229 15121 15285
rect 15049 15195 15068 15229
rect 15102 15195 15121 15229
rect 15049 15139 15121 15195
rect 15049 15105 15068 15139
rect 15102 15105 15121 15139
rect 14159 15034 14178 15068
rect 14212 15034 14231 15068
rect 14159 15020 14231 15034
rect 15049 15049 15121 15105
rect 15049 15020 15068 15049
rect 14063 15015 15068 15020
rect 15102 15020 15121 15049
rect 15185 15858 15284 15914
rect 15185 15824 15216 15858
rect 15250 15824 15284 15858
rect 15185 15768 15284 15824
rect 15185 15734 15216 15768
rect 15250 15734 15284 15768
rect 15185 15678 15284 15734
rect 15185 15644 15216 15678
rect 15250 15644 15284 15678
rect 15185 15588 15284 15644
rect 15185 15554 15216 15588
rect 15250 15554 15284 15588
rect 15185 15498 15284 15554
rect 15185 15464 15216 15498
rect 15250 15464 15284 15498
rect 15185 15408 15284 15464
rect 15185 15374 15216 15408
rect 15250 15374 15284 15408
rect 15185 15318 15284 15374
rect 15185 15284 15216 15318
rect 15250 15284 15284 15318
rect 15185 15228 15284 15284
rect 15185 15194 15216 15228
rect 15250 15194 15284 15228
rect 15185 15138 15284 15194
rect 15185 15104 15216 15138
rect 15250 15104 15284 15138
rect 15185 15048 15284 15104
rect 15185 15020 15216 15048
rect 15102 15015 15216 15020
rect 14063 15014 15216 15015
rect 15250 15020 15284 15048
rect 15250 15014 15290 15020
rect 11270 14992 15290 15014
rect 11270 14958 11516 14992
rect 11550 14958 11606 14992
rect 11640 14958 11696 14992
rect 11730 14958 11786 14992
rect 11820 14958 11876 14992
rect 11910 14958 11966 14992
rect 12000 14958 12056 14992
rect 12090 14958 12146 14992
rect 12180 14958 12236 14992
rect 12270 14958 12876 14992
rect 12910 14958 12966 14992
rect 13000 14958 13056 14992
rect 13090 14958 13146 14992
rect 13180 14958 13236 14992
rect 13270 14958 13326 14992
rect 13360 14958 13416 14992
rect 13450 14958 13506 14992
rect 13540 14958 13596 14992
rect 13630 14958 14236 14992
rect 14270 14958 14326 14992
rect 14360 14958 14416 14992
rect 14450 14958 14506 14992
rect 14540 14958 14596 14992
rect 14630 14958 14686 14992
rect 14720 14958 14776 14992
rect 14810 14958 14866 14992
rect 14900 14958 14956 14992
rect 14990 14958 15290 14992
rect 11270 14924 11309 14958
rect 11343 14924 12496 14958
rect 12530 14924 12669 14958
rect 12703 14924 13856 14958
rect 13890 14924 14029 14958
rect 14063 14924 15216 14958
rect 15250 14924 15290 14958
rect 11270 14868 15290 14924
rect 11270 14834 11309 14868
rect 11343 14845 12496 14868
rect 11343 14834 11410 14845
rect 11270 14811 11410 14834
rect 11444 14811 11500 14845
rect 11534 14811 11590 14845
rect 11624 14811 11680 14845
rect 11714 14811 11770 14845
rect 11804 14811 11860 14845
rect 11894 14811 11950 14845
rect 11984 14811 12040 14845
rect 12074 14811 12130 14845
rect 12164 14811 12220 14845
rect 12254 14811 12310 14845
rect 12344 14811 12400 14845
rect 12434 14834 12496 14845
rect 12530 14834 12669 14868
rect 12703 14845 13856 14868
rect 12703 14834 12770 14845
rect 12434 14811 12770 14834
rect 12804 14811 12860 14845
rect 12894 14811 12950 14845
rect 12984 14811 13040 14845
rect 13074 14811 13130 14845
rect 13164 14811 13220 14845
rect 13254 14811 13310 14845
rect 13344 14811 13400 14845
rect 13434 14811 13490 14845
rect 13524 14811 13580 14845
rect 13614 14811 13670 14845
rect 13704 14811 13760 14845
rect 13794 14834 13856 14845
rect 13890 14834 14029 14868
rect 14063 14845 15216 14868
rect 14063 14834 14130 14845
rect 13794 14811 14130 14834
rect 14164 14811 14220 14845
rect 14254 14811 14310 14845
rect 14344 14811 14400 14845
rect 14434 14811 14490 14845
rect 14524 14811 14580 14845
rect 14614 14811 14670 14845
rect 14704 14811 14760 14845
rect 14794 14811 14850 14845
rect 14884 14811 14940 14845
rect 14974 14811 15030 14845
rect 15064 14811 15120 14845
rect 15154 14834 15216 14845
rect 15250 14834 15290 14868
rect 15154 14811 15290 14834
rect 11270 14770 15290 14811
rect 12542 14600 12632 14610
rect 12542 14550 12562 14600
rect 12612 14550 12632 14600
rect 12542 14540 12632 14550
rect 13940 14600 14030 14610
rect 13940 14550 13960 14600
rect 14010 14550 14030 14600
rect 13940 14540 14030 14550
rect 11170 14250 11230 14270
rect 11170 14220 11180 14250
rect 11080 14210 11180 14220
rect 11220 14210 11230 14250
rect 11080 14200 11230 14210
rect 11080 14160 11100 14200
rect 11140 14160 11230 14200
rect 11080 14150 11230 14160
rect 11080 14140 11180 14150
rect 11170 14110 11180 14140
rect 11220 14110 11230 14150
rect 11170 14090 11230 14110
rect 13250 14250 13310 14270
rect 13250 14210 13260 14250
rect 13300 14210 13310 14250
rect 13250 14150 13310 14210
rect 13250 14110 13260 14150
rect 13300 14110 13310 14150
rect 13250 14090 13310 14110
rect 15330 14260 15470 14270
rect 15330 14250 15550 14260
rect 15330 14210 15340 14250
rect 15380 14210 15420 14250
rect 15460 14240 15550 14250
rect 15460 14210 15490 14240
rect 15330 14200 15490 14210
rect 15530 14200 15550 14240
rect 15330 14160 15550 14200
rect 15330 14150 15490 14160
rect 15330 14110 15340 14150
rect 15380 14110 15420 14150
rect 15460 14120 15490 14150
rect 15530 14120 15550 14160
rect 15460 14110 15550 14120
rect 15330 14100 15550 14110
rect 15330 14090 15470 14100
rect 11180 14050 11220 14090
rect 13260 14050 13300 14090
rect 11160 14030 11240 14050
rect 11160 13990 11180 14030
rect 11220 13990 11240 14030
rect 11160 13970 11240 13990
rect 11320 14030 11400 14050
rect 11320 13990 11340 14030
rect 11380 13990 11400 14030
rect 11320 13970 11400 13990
rect 11480 14030 11560 14050
rect 11480 13990 11500 14030
rect 11540 13990 11560 14030
rect 11480 13970 11560 13990
rect 11640 14030 11720 14050
rect 11640 13990 11660 14030
rect 11700 13990 11720 14030
rect 11640 13970 11720 13990
rect 11800 14030 11880 14050
rect 11800 13990 11820 14030
rect 11860 13990 11880 14030
rect 11800 13970 11880 13990
rect 11960 14030 12040 14050
rect 11960 13990 11980 14030
rect 12020 13990 12040 14030
rect 11960 13970 12040 13990
rect 12120 14030 12200 14050
rect 12120 13990 12140 14030
rect 12180 13990 12200 14030
rect 12120 13970 12200 13990
rect 12280 14030 12360 14050
rect 12280 13990 12300 14030
rect 12340 13990 12360 14030
rect 12280 13970 12360 13990
rect 12440 14030 12520 14050
rect 12440 13990 12460 14030
rect 12500 13990 12520 14030
rect 12440 13970 12520 13990
rect 12600 14030 12680 14050
rect 12600 13990 12620 14030
rect 12660 13990 12680 14030
rect 12600 13970 12680 13990
rect 12760 14030 12840 14050
rect 12760 13990 12780 14030
rect 12820 13990 12840 14030
rect 12760 13970 12840 13990
rect 12920 14030 13000 14050
rect 12920 13990 12940 14030
rect 12980 13990 13000 14030
rect 12920 13970 13000 13990
rect 13080 14030 13160 14050
rect 13080 13990 13100 14030
rect 13140 13990 13160 14030
rect 13080 13970 13160 13990
rect 13240 14030 13320 14050
rect 13240 13990 13260 14030
rect 13300 13990 13320 14030
rect 13240 13970 13320 13990
rect 13400 14030 13480 14050
rect 13400 13990 13420 14030
rect 13460 13990 13480 14030
rect 13400 13970 13480 13990
rect 13560 14030 13640 14050
rect 13560 13990 13580 14030
rect 13620 13990 13640 14030
rect 13560 13970 13640 13990
rect 13720 14030 13800 14050
rect 13720 13990 13740 14030
rect 13780 13990 13800 14030
rect 13720 13970 13800 13990
rect 13880 14030 13960 14050
rect 13880 13990 13900 14030
rect 13940 13990 13960 14030
rect 13880 13970 13960 13990
rect 14040 14030 14120 14050
rect 14040 13990 14060 14030
rect 14100 13990 14120 14030
rect 14040 13970 14120 13990
rect 14200 14030 14280 14050
rect 14200 13990 14220 14030
rect 14260 13990 14280 14030
rect 14200 13970 14280 13990
rect 14360 14030 14440 14050
rect 14360 13990 14380 14030
rect 14420 13990 14440 14030
rect 14360 13970 14440 13990
rect 14520 14030 14600 14050
rect 14520 13990 14540 14030
rect 14580 13990 14600 14030
rect 14520 13970 14600 13990
rect 14680 14030 14760 14050
rect 14680 13990 14700 14030
rect 14740 13990 14760 14030
rect 14680 13970 14760 13990
rect 14840 14030 14920 14050
rect 14840 13990 14860 14030
rect 14900 13990 14920 14030
rect 14840 13970 14920 13990
rect 15000 14030 15080 14050
rect 15000 13990 15020 14030
rect 15060 13990 15080 14030
rect 15000 13970 15080 13990
rect 15160 14030 15240 14050
rect 15160 13990 15180 14030
rect 15220 13990 15240 14030
rect 15160 13970 15240 13990
rect 11900 13760 11980 13780
rect 11900 13720 11920 13760
rect 11960 13720 11980 13760
rect 11900 13660 11980 13720
rect 14580 13760 14660 13780
rect 14580 13720 14600 13760
rect 14640 13720 14660 13760
rect 14580 13660 14660 13720
rect 10750 13640 10810 13660
rect 10750 13600 10760 13640
rect 10800 13600 10810 13640
rect 10750 13540 10810 13600
rect 10750 13500 10760 13540
rect 10800 13500 10810 13540
rect 10750 13440 10810 13500
rect 10750 13400 10760 13440
rect 10800 13400 10810 13440
rect 10750 13340 10810 13400
rect 10750 13300 10760 13340
rect 10800 13300 10810 13340
rect 10750 13240 10810 13300
rect 10750 13200 10760 13240
rect 10800 13200 10810 13240
rect 10750 13180 10810 13200
rect 11830 13640 12050 13660
rect 11830 13600 11840 13640
rect 11880 13600 11920 13640
rect 11960 13600 12000 13640
rect 12040 13600 12050 13640
rect 11830 13540 12050 13600
rect 11830 13500 11840 13540
rect 11880 13500 11920 13540
rect 11960 13500 12000 13540
rect 12040 13500 12050 13540
rect 11830 13440 12050 13500
rect 11830 13400 11840 13440
rect 11880 13400 11920 13440
rect 11960 13400 12000 13440
rect 12040 13400 12050 13440
rect 11830 13340 12050 13400
rect 11830 13300 11840 13340
rect 11880 13300 11920 13340
rect 11960 13300 12000 13340
rect 12040 13300 12050 13340
rect 11830 13240 12050 13300
rect 11830 13200 11840 13240
rect 11880 13200 11920 13240
rect 11960 13200 12000 13240
rect 12040 13200 12050 13240
rect 11830 13180 12050 13200
rect 13070 13640 13130 13660
rect 13070 13600 13080 13640
rect 13120 13600 13130 13640
rect 13070 13540 13130 13600
rect 13070 13500 13080 13540
rect 13120 13500 13130 13540
rect 13070 13440 13130 13500
rect 13070 13400 13080 13440
rect 13120 13400 13130 13440
rect 13070 13340 13130 13400
rect 13070 13300 13080 13340
rect 13120 13300 13130 13340
rect 13070 13240 13130 13300
rect 13070 13200 13080 13240
rect 13120 13200 13130 13240
rect 10740 13160 10820 13180
rect 10740 13120 10760 13160
rect 10800 13120 10820 13160
rect 13070 13150 13130 13200
rect 10740 13100 10820 13120
rect 10920 13120 11000 13140
rect 10920 13080 10940 13120
rect 10980 13080 11000 13120
rect 10920 13060 11000 13080
rect 11160 13120 11240 13140
rect 11160 13080 11180 13120
rect 11220 13080 11240 13120
rect 11160 13060 11240 13080
rect 11400 13120 11480 13140
rect 11400 13080 11420 13120
rect 11460 13080 11480 13120
rect 11400 13060 11480 13080
rect 11640 13120 11720 13140
rect 11640 13080 11660 13120
rect 11700 13080 11720 13120
rect 11640 13060 11720 13080
rect 12280 13120 12360 13140
rect 12280 13080 12300 13120
rect 12340 13080 12360 13120
rect 12280 13060 12360 13080
rect 12520 13120 12600 13140
rect 12520 13080 12540 13120
rect 12580 13080 12600 13120
rect 12520 13060 12600 13080
rect 12760 13120 12840 13140
rect 12760 13080 12780 13120
rect 12820 13080 12840 13120
rect 13070 13110 13080 13150
rect 13120 13110 13130 13150
rect 13070 13090 13130 13110
rect 13430 13640 13490 13660
rect 13430 13600 13440 13640
rect 13480 13600 13490 13640
rect 13430 13540 13490 13600
rect 13430 13500 13440 13540
rect 13480 13500 13490 13540
rect 13430 13440 13490 13500
rect 13430 13400 13440 13440
rect 13480 13400 13490 13440
rect 13430 13340 13490 13400
rect 13430 13300 13440 13340
rect 13480 13300 13490 13340
rect 13430 13240 13490 13300
rect 13430 13200 13440 13240
rect 13480 13200 13490 13240
rect 13430 13150 13490 13200
rect 14510 13640 14730 13660
rect 14510 13600 14520 13640
rect 14560 13600 14600 13640
rect 14640 13600 14680 13640
rect 14720 13600 14730 13640
rect 14510 13540 14730 13600
rect 14510 13500 14520 13540
rect 14560 13500 14600 13540
rect 14640 13500 14680 13540
rect 14720 13500 14730 13540
rect 14510 13440 14730 13500
rect 14510 13400 14520 13440
rect 14560 13400 14600 13440
rect 14640 13400 14680 13440
rect 14720 13400 14730 13440
rect 14510 13340 14730 13400
rect 14510 13300 14520 13340
rect 14560 13300 14600 13340
rect 14640 13300 14680 13340
rect 14720 13300 14730 13340
rect 14510 13240 14730 13300
rect 14510 13200 14520 13240
rect 14560 13200 14600 13240
rect 14640 13200 14680 13240
rect 14720 13200 14730 13240
rect 14510 13180 14730 13200
rect 15750 13640 15810 13660
rect 15750 13600 15760 13640
rect 15800 13600 15810 13640
rect 15750 13540 15810 13600
rect 15750 13500 15760 13540
rect 15800 13500 15810 13540
rect 15750 13440 15810 13500
rect 15750 13400 15760 13440
rect 15800 13400 15810 13440
rect 15750 13340 15810 13400
rect 15750 13300 15760 13340
rect 15800 13300 15810 13340
rect 15750 13240 15810 13300
rect 15750 13200 15760 13240
rect 15800 13200 15810 13240
rect 15750 13180 15810 13200
rect 13430 13110 13440 13150
rect 13480 13110 13490 13150
rect 13430 13090 13490 13110
rect 13720 13120 13800 13140
rect 12760 13060 12840 13080
rect 13720 13080 13740 13120
rect 13780 13080 13800 13120
rect 13720 13060 13800 13080
rect 13960 13120 14040 13140
rect 13960 13080 13980 13120
rect 14020 13080 14040 13120
rect 13960 13060 14040 13080
rect 14200 13120 14280 13140
rect 14200 13080 14220 13120
rect 14260 13080 14280 13120
rect 14200 13060 14280 13080
rect 14840 13120 14920 13140
rect 14840 13080 14860 13120
rect 14900 13080 14920 13120
rect 14840 13060 14920 13080
rect 15080 13120 15160 13140
rect 15080 13080 15100 13120
rect 15140 13080 15160 13120
rect 15080 13060 15160 13080
rect 15320 13120 15400 13140
rect 15320 13080 15340 13120
rect 15380 13080 15400 13120
rect 15320 13060 15400 13080
rect 15560 13120 15640 13140
rect 15560 13080 15580 13120
rect 15620 13080 15640 13120
rect 15560 13060 15640 13080
rect 11431 12742 11489 12760
rect 11431 12708 11443 12742
rect 11477 12708 11489 12742
rect 11431 12690 11489 12708
rect 11791 12742 11849 12760
rect 11791 12708 11803 12742
rect 11837 12708 11849 12742
rect 11791 12690 11849 12708
rect 11911 12742 11969 12760
rect 11911 12708 11923 12742
rect 11957 12708 11969 12742
rect 11911 12690 11969 12708
rect 12271 12742 12329 12760
rect 12271 12708 12283 12742
rect 12317 12708 12329 12742
rect 12271 12690 12329 12708
rect 12391 12742 12449 12760
rect 12391 12708 12403 12742
rect 12437 12708 12449 12742
rect 14111 12742 14169 12760
rect 12391 12690 12449 12708
rect 12800 12720 12880 12740
rect 12800 12680 12820 12720
rect 12860 12680 12880 12720
rect 11370 12630 11430 12650
rect 11370 12590 11380 12630
rect 11420 12590 11430 12630
rect 11370 12570 11430 12590
rect 11490 12630 11550 12650
rect 11490 12590 11500 12630
rect 11540 12590 11550 12630
rect 11490 12570 11550 12590
rect 11610 12630 11670 12650
rect 11610 12590 11620 12630
rect 11660 12590 11670 12630
rect 11610 12570 11670 12590
rect 11730 12630 11790 12650
rect 11730 12590 11740 12630
rect 11780 12590 11790 12630
rect 11730 12570 11790 12590
rect 11850 12630 11910 12650
rect 11850 12590 11860 12630
rect 11900 12590 11910 12630
rect 11850 12570 11910 12590
rect 11970 12630 12030 12650
rect 11970 12590 11980 12630
rect 12020 12590 12030 12630
rect 11970 12570 12030 12590
rect 12090 12630 12150 12650
rect 12090 12590 12100 12630
rect 12140 12590 12150 12630
rect 12090 12570 12150 12590
rect 12210 12630 12270 12650
rect 12210 12590 12220 12630
rect 12260 12590 12270 12630
rect 12210 12570 12270 12590
rect 12330 12630 12390 12650
rect 12330 12590 12340 12630
rect 12380 12590 12390 12630
rect 12330 12570 12390 12590
rect 12450 12630 12510 12650
rect 12450 12590 12460 12630
rect 12500 12590 12510 12630
rect 12450 12570 12510 12590
rect 12570 12630 12630 12650
rect 12570 12590 12580 12630
rect 12620 12590 12630 12630
rect 12570 12570 12630 12590
rect 12800 12640 12880 12680
rect 12800 12600 12820 12640
rect 12860 12600 12880 12640
rect 12800 12560 12880 12600
rect 11532 12512 11590 12530
rect 11532 12478 11544 12512
rect 11578 12478 11590 12512
rect 11532 12460 11590 12478
rect 11690 12512 11748 12530
rect 11690 12478 11702 12512
rect 11736 12478 11748 12512
rect 11690 12460 11748 12478
rect 12014 12512 12072 12530
rect 12014 12478 12026 12512
rect 12060 12478 12072 12512
rect 12014 12460 12072 12478
rect 12168 12512 12226 12530
rect 12168 12478 12180 12512
rect 12214 12478 12226 12512
rect 12168 12460 12226 12478
rect 12492 12512 12550 12530
rect 12492 12478 12504 12512
rect 12538 12478 12550 12512
rect 12800 12520 12820 12560
rect 12860 12520 12880 12560
rect 12800 12500 12880 12520
rect 13680 12720 13760 12740
rect 13680 12680 13700 12720
rect 13740 12680 13760 12720
rect 14111 12708 14123 12742
rect 14157 12708 14169 12742
rect 14111 12690 14169 12708
rect 14231 12742 14289 12760
rect 14231 12708 14243 12742
rect 14277 12708 14289 12742
rect 14231 12690 14289 12708
rect 14591 12742 14649 12760
rect 14591 12708 14603 12742
rect 14637 12708 14649 12742
rect 14591 12690 14649 12708
rect 14711 12742 14769 12760
rect 14711 12708 14723 12742
rect 14757 12708 14769 12742
rect 14711 12690 14769 12708
rect 15071 12742 15129 12760
rect 15071 12708 15083 12742
rect 15117 12708 15129 12742
rect 15071 12690 15129 12708
rect 13680 12640 13760 12680
rect 13680 12600 13700 12640
rect 13740 12600 13760 12640
rect 13680 12560 13760 12600
rect 13930 12630 13990 12650
rect 13930 12590 13940 12630
rect 13980 12590 13990 12630
rect 13930 12570 13990 12590
rect 14050 12630 14110 12650
rect 14050 12590 14060 12630
rect 14100 12590 14110 12630
rect 14050 12570 14110 12590
rect 14170 12630 14230 12650
rect 14170 12590 14180 12630
rect 14220 12590 14230 12630
rect 14170 12570 14230 12590
rect 14290 12630 14350 12650
rect 14290 12590 14300 12630
rect 14340 12590 14350 12630
rect 14290 12570 14350 12590
rect 14410 12630 14470 12650
rect 14410 12590 14420 12630
rect 14460 12590 14470 12630
rect 14410 12570 14470 12590
rect 14530 12630 14590 12650
rect 14530 12590 14540 12630
rect 14580 12590 14590 12630
rect 14530 12570 14590 12590
rect 14650 12630 14710 12650
rect 14650 12590 14660 12630
rect 14700 12590 14710 12630
rect 14650 12570 14710 12590
rect 14770 12630 14830 12650
rect 14770 12590 14780 12630
rect 14820 12590 14830 12630
rect 14770 12570 14830 12590
rect 14890 12630 14950 12650
rect 14890 12590 14900 12630
rect 14940 12590 14950 12630
rect 14890 12570 14950 12590
rect 15010 12630 15070 12650
rect 15010 12590 15020 12630
rect 15060 12590 15070 12630
rect 15010 12570 15070 12590
rect 15130 12630 15190 12650
rect 15130 12590 15140 12630
rect 15180 12590 15190 12630
rect 15130 12570 15190 12590
rect 13680 12520 13700 12560
rect 13740 12520 13760 12560
rect 13680 12500 13760 12520
rect 14010 12512 14068 12530
rect 12492 12460 12550 12478
rect 14010 12478 14022 12512
rect 14056 12478 14068 12512
rect 14010 12460 14068 12478
rect 14334 12512 14392 12530
rect 14334 12478 14346 12512
rect 14380 12478 14392 12512
rect 14334 12460 14392 12478
rect 14488 12512 14546 12530
rect 14488 12478 14500 12512
rect 14534 12478 14546 12512
rect 14488 12460 14546 12478
rect 14812 12512 14870 12530
rect 14812 12478 14824 12512
rect 14858 12478 14870 12512
rect 14812 12460 14870 12478
rect 14970 12512 15028 12530
rect 14970 12478 14982 12512
rect 15016 12478 15028 12512
rect 14970 12460 15028 12478
rect 10710 11920 10770 11940
rect 10710 11880 10720 11920
rect 10760 11880 10770 11920
rect 10710 11860 10770 11880
rect 10880 11910 10960 11930
rect 10880 11870 10900 11910
rect 10940 11870 10960 11910
rect 10880 11850 10960 11870
rect 11370 11910 11430 11930
rect 11370 11870 11380 11910
rect 11420 11870 11430 11910
rect 11370 11850 11430 11870
rect 11600 11910 11680 11930
rect 11600 11870 11620 11910
rect 11660 11870 11680 11910
rect 11600 11850 11680 11870
rect 12090 11910 12150 11930
rect 12090 11870 12100 11910
rect 12140 11870 12150 11910
rect 12090 11850 12150 11870
rect 12320 11910 12400 11930
rect 12320 11870 12340 11910
rect 12380 11870 12400 11910
rect 12320 11850 12400 11870
rect 12750 11910 12810 11930
rect 12750 11870 12760 11910
rect 12800 11870 12810 11910
rect 12750 11850 12810 11870
rect 13750 11910 13810 11930
rect 13750 11870 13760 11910
rect 13800 11870 13810 11910
rect 13750 11850 13810 11870
rect 14160 11910 14240 11930
rect 14160 11870 14180 11910
rect 14220 11870 14240 11910
rect 14160 11850 14240 11870
rect 14410 11910 14470 11930
rect 14410 11870 14420 11910
rect 14460 11870 14470 11910
rect 14410 11850 14470 11870
rect 14880 11910 14960 11930
rect 14880 11870 14900 11910
rect 14940 11870 14960 11910
rect 14880 11850 14960 11870
rect 15130 11910 15190 11930
rect 15130 11870 15140 11910
rect 15180 11870 15190 11910
rect 15130 11850 15190 11870
rect 15600 11910 15680 11930
rect 15600 11870 15620 11910
rect 15660 11870 15680 11910
rect 15600 11850 15680 11870
rect 15790 11920 15850 11940
rect 15790 11880 15800 11920
rect 15840 11880 15850 11920
rect 15790 11860 15850 11880
rect 10450 11790 10590 11810
rect 10450 11750 10460 11790
rect 10500 11750 10540 11790
rect 10580 11750 10590 11790
rect 10450 11690 10590 11750
rect 10450 11650 10460 11690
rect 10500 11650 10540 11690
rect 10580 11650 10590 11690
rect 10450 11630 10590 11650
rect 10650 11790 10710 11810
rect 10650 11750 10660 11790
rect 10700 11750 10710 11790
rect 10650 11690 10710 11750
rect 10650 11650 10660 11690
rect 10700 11650 10710 11690
rect 10650 11630 10710 11650
rect 10770 11790 10830 11810
rect 10770 11750 10780 11790
rect 10820 11750 10830 11790
rect 10770 11690 10830 11750
rect 10770 11650 10780 11690
rect 10820 11650 10830 11690
rect 10770 11630 10830 11650
rect 10890 11790 10950 11810
rect 10890 11750 10900 11790
rect 10940 11750 10950 11790
rect 10890 11690 10950 11750
rect 10890 11650 10900 11690
rect 10940 11650 10950 11690
rect 10890 11630 10950 11650
rect 11010 11790 11070 11810
rect 11010 11750 11020 11790
rect 11060 11750 11070 11790
rect 11010 11690 11070 11750
rect 11010 11650 11020 11690
rect 11060 11650 11070 11690
rect 11010 11630 11070 11650
rect 11130 11790 11190 11810
rect 11130 11750 11140 11790
rect 11180 11750 11190 11790
rect 11130 11690 11190 11750
rect 11130 11650 11140 11690
rect 11180 11650 11190 11690
rect 11130 11630 11190 11650
rect 11250 11790 11310 11810
rect 11250 11750 11260 11790
rect 11300 11750 11310 11790
rect 11250 11690 11310 11750
rect 11250 11650 11260 11690
rect 11300 11650 11310 11690
rect 11250 11630 11310 11650
rect 11370 11790 11430 11810
rect 11370 11750 11380 11790
rect 11420 11750 11430 11790
rect 11370 11690 11430 11750
rect 11370 11650 11380 11690
rect 11420 11650 11430 11690
rect 11370 11630 11430 11650
rect 11490 11790 11550 11810
rect 11490 11750 11500 11790
rect 11540 11750 11550 11790
rect 11490 11690 11550 11750
rect 11490 11650 11500 11690
rect 11540 11650 11550 11690
rect 11490 11630 11550 11650
rect 11610 11790 11670 11810
rect 11610 11750 11620 11790
rect 11660 11750 11670 11790
rect 11610 11690 11670 11750
rect 11610 11650 11620 11690
rect 11660 11650 11670 11690
rect 11610 11630 11670 11650
rect 11730 11790 11790 11810
rect 11730 11750 11740 11790
rect 11780 11750 11790 11790
rect 11730 11690 11790 11750
rect 11730 11650 11740 11690
rect 11780 11650 11790 11690
rect 11730 11630 11790 11650
rect 11850 11790 11910 11810
rect 11850 11750 11860 11790
rect 11900 11750 11910 11790
rect 11850 11690 11910 11750
rect 11850 11650 11860 11690
rect 11900 11650 11910 11690
rect 11850 11630 11910 11650
rect 11970 11790 12030 11810
rect 11970 11750 11980 11790
rect 12020 11750 12030 11790
rect 11970 11690 12030 11750
rect 11970 11650 11980 11690
rect 12020 11650 12030 11690
rect 11970 11630 12030 11650
rect 12090 11790 12150 11810
rect 12090 11750 12100 11790
rect 12140 11750 12150 11790
rect 12090 11690 12150 11750
rect 12090 11650 12100 11690
rect 12140 11650 12150 11690
rect 12090 11630 12150 11650
rect 12210 11790 12270 11810
rect 12210 11750 12220 11790
rect 12260 11750 12270 11790
rect 12210 11690 12270 11750
rect 12210 11650 12220 11690
rect 12260 11650 12270 11690
rect 12210 11630 12270 11650
rect 12330 11790 12390 11810
rect 12330 11750 12340 11790
rect 12380 11750 12390 11790
rect 12330 11690 12390 11750
rect 12330 11650 12340 11690
rect 12380 11650 12390 11690
rect 12330 11630 12390 11650
rect 12450 11790 12510 11810
rect 12450 11750 12460 11790
rect 12500 11750 12510 11790
rect 12450 11690 12510 11750
rect 12450 11650 12460 11690
rect 12500 11650 12510 11690
rect 12450 11630 12510 11650
rect 12570 11790 12630 11810
rect 12570 11750 12580 11790
rect 12620 11750 12630 11790
rect 12570 11690 12630 11750
rect 12570 11650 12580 11690
rect 12620 11650 12630 11690
rect 12570 11630 12630 11650
rect 12690 11790 12750 11810
rect 12690 11750 12700 11790
rect 12740 11750 12750 11790
rect 12690 11690 12750 11750
rect 12690 11650 12700 11690
rect 12740 11650 12750 11690
rect 12690 11630 12750 11650
rect 12810 11790 12870 11810
rect 12810 11750 12820 11790
rect 12860 11750 12870 11790
rect 12810 11690 12870 11750
rect 12810 11650 12820 11690
rect 12860 11650 12870 11690
rect 12810 11630 12870 11650
rect 12930 11790 13070 11810
rect 12930 11750 12940 11790
rect 12980 11750 13020 11790
rect 13060 11750 13070 11790
rect 12930 11690 13070 11750
rect 12930 11650 12940 11690
rect 12980 11650 13020 11690
rect 13060 11650 13070 11690
rect 12930 11630 13070 11650
rect 13490 11790 13630 11810
rect 13490 11750 13500 11790
rect 13540 11750 13580 11790
rect 13620 11750 13630 11790
rect 13490 11690 13630 11750
rect 13490 11650 13500 11690
rect 13540 11650 13580 11690
rect 13620 11650 13630 11690
rect 13490 11630 13630 11650
rect 13690 11790 13750 11810
rect 13690 11750 13700 11790
rect 13740 11750 13750 11790
rect 13690 11690 13750 11750
rect 13690 11650 13700 11690
rect 13740 11650 13750 11690
rect 13690 11630 13750 11650
rect 13810 11790 13870 11810
rect 13810 11750 13820 11790
rect 13860 11750 13870 11790
rect 13810 11690 13870 11750
rect 13810 11650 13820 11690
rect 13860 11650 13870 11690
rect 13810 11630 13870 11650
rect 13930 11790 13990 11810
rect 13930 11750 13940 11790
rect 13980 11750 13990 11790
rect 13930 11690 13990 11750
rect 13930 11650 13940 11690
rect 13980 11650 13990 11690
rect 13930 11630 13990 11650
rect 14050 11790 14110 11810
rect 14050 11750 14060 11790
rect 14100 11750 14110 11790
rect 14050 11690 14110 11750
rect 14050 11650 14060 11690
rect 14100 11650 14110 11690
rect 14050 11630 14110 11650
rect 14170 11790 14230 11810
rect 14170 11750 14180 11790
rect 14220 11750 14230 11790
rect 14170 11690 14230 11750
rect 14170 11650 14180 11690
rect 14220 11650 14230 11690
rect 14170 11630 14230 11650
rect 14290 11790 14350 11810
rect 14290 11750 14300 11790
rect 14340 11750 14350 11790
rect 14290 11690 14350 11750
rect 14290 11650 14300 11690
rect 14340 11650 14350 11690
rect 14290 11630 14350 11650
rect 14410 11790 14470 11810
rect 14410 11750 14420 11790
rect 14460 11750 14470 11790
rect 14410 11690 14470 11750
rect 14410 11650 14420 11690
rect 14460 11650 14470 11690
rect 14410 11630 14470 11650
rect 14530 11790 14590 11810
rect 14530 11750 14540 11790
rect 14580 11750 14590 11790
rect 14530 11690 14590 11750
rect 14530 11650 14540 11690
rect 14580 11650 14590 11690
rect 14530 11630 14590 11650
rect 14650 11790 14710 11810
rect 14650 11750 14660 11790
rect 14700 11750 14710 11790
rect 14650 11690 14710 11750
rect 14650 11650 14660 11690
rect 14700 11650 14710 11690
rect 14650 11630 14710 11650
rect 14770 11790 14830 11810
rect 14770 11750 14780 11790
rect 14820 11750 14830 11790
rect 14770 11690 14830 11750
rect 14770 11650 14780 11690
rect 14820 11650 14830 11690
rect 14770 11630 14830 11650
rect 14890 11790 14950 11810
rect 14890 11750 14900 11790
rect 14940 11750 14950 11790
rect 14890 11690 14950 11750
rect 14890 11650 14900 11690
rect 14940 11650 14950 11690
rect 14890 11630 14950 11650
rect 15010 11790 15070 11810
rect 15010 11750 15020 11790
rect 15060 11750 15070 11790
rect 15010 11690 15070 11750
rect 15010 11650 15020 11690
rect 15060 11650 15070 11690
rect 15010 11630 15070 11650
rect 15130 11790 15190 11810
rect 15130 11750 15140 11790
rect 15180 11750 15190 11790
rect 15130 11690 15190 11750
rect 15130 11650 15140 11690
rect 15180 11650 15190 11690
rect 15130 11630 15190 11650
rect 15250 11790 15310 11810
rect 15250 11750 15260 11790
rect 15300 11750 15310 11790
rect 15250 11690 15310 11750
rect 15250 11650 15260 11690
rect 15300 11650 15310 11690
rect 15250 11630 15310 11650
rect 15370 11790 15430 11810
rect 15370 11750 15380 11790
rect 15420 11750 15430 11790
rect 15370 11690 15430 11750
rect 15370 11650 15380 11690
rect 15420 11650 15430 11690
rect 15370 11630 15430 11650
rect 15490 11790 15550 11810
rect 15490 11750 15500 11790
rect 15540 11750 15550 11790
rect 15490 11690 15550 11750
rect 15490 11650 15500 11690
rect 15540 11650 15550 11690
rect 15490 11630 15550 11650
rect 15610 11790 15670 11810
rect 15610 11750 15620 11790
rect 15660 11750 15670 11790
rect 15610 11690 15670 11750
rect 15610 11650 15620 11690
rect 15660 11650 15670 11690
rect 15610 11630 15670 11650
rect 15730 11790 15790 11810
rect 15730 11750 15740 11790
rect 15780 11750 15790 11790
rect 15730 11690 15790 11750
rect 15730 11650 15740 11690
rect 15780 11650 15790 11690
rect 15730 11630 15790 11650
rect 15850 11790 15910 11810
rect 15850 11750 15860 11790
rect 15900 11750 15910 11790
rect 15850 11690 15910 11750
rect 15850 11650 15860 11690
rect 15900 11650 15910 11690
rect 15850 11630 15910 11650
rect 15970 11790 16110 11810
rect 15970 11750 15980 11790
rect 16020 11750 16060 11790
rect 16100 11750 16110 11790
rect 15970 11690 16110 11750
rect 15970 11650 15980 11690
rect 16020 11650 16060 11690
rect 16100 11650 16110 11690
rect 15970 11630 16110 11650
rect 10530 11570 10590 11590
rect 10530 11530 10540 11570
rect 10580 11530 10590 11570
rect 10530 11510 10590 11530
rect 12930 11570 12990 11590
rect 12930 11530 12940 11570
rect 12980 11530 12990 11570
rect 12930 11510 12990 11530
rect 13570 11570 13630 11590
rect 13570 11530 13580 11570
rect 13620 11530 13630 11570
rect 13570 11510 13630 11530
rect 15970 11570 16030 11590
rect 15970 11530 15980 11570
rect 16020 11530 16030 11570
rect 15970 11510 16030 11530
rect 11900 10750 11970 10770
rect 11900 10710 11910 10750
rect 11950 10710 11970 10750
rect 11900 10690 11970 10710
rect 12070 10750 12150 10770
rect 12070 10710 12090 10750
rect 12130 10710 12150 10750
rect 12070 10690 12150 10710
rect 12250 10750 12330 10770
rect 12250 10710 12270 10750
rect 12310 10710 12330 10750
rect 12250 10690 12330 10710
rect 12430 10750 12510 10770
rect 12430 10710 12450 10750
rect 12490 10710 12510 10750
rect 12430 10690 12510 10710
rect 12610 10750 12690 10770
rect 12610 10710 12630 10750
rect 12670 10710 12690 10750
rect 12610 10690 12690 10710
rect 12790 10750 12870 10770
rect 12790 10710 12810 10750
rect 12850 10710 12870 10750
rect 12790 10690 12870 10710
rect 12970 10750 13050 10770
rect 12970 10710 12990 10750
rect 13030 10710 13050 10750
rect 12970 10690 13050 10710
rect 13150 10750 13220 10770
rect 13150 10710 13170 10750
rect 13210 10710 13220 10750
rect 13150 10690 13220 10710
rect 13340 10750 13410 10770
rect 13340 10710 13350 10750
rect 13390 10710 13410 10750
rect 13340 10690 13410 10710
rect 13510 10750 13590 10770
rect 13510 10710 13530 10750
rect 13570 10710 13590 10750
rect 13510 10690 13590 10710
rect 13690 10750 13770 10770
rect 13690 10710 13710 10750
rect 13750 10710 13770 10750
rect 13690 10690 13770 10710
rect 13870 10750 13950 10770
rect 13870 10710 13890 10750
rect 13930 10710 13950 10750
rect 13870 10690 13950 10710
rect 14050 10750 14130 10770
rect 14050 10710 14070 10750
rect 14110 10710 14130 10750
rect 14050 10690 14130 10710
rect 14230 10750 14310 10770
rect 14230 10710 14250 10750
rect 14290 10710 14310 10750
rect 14230 10690 14310 10710
rect 14410 10750 14490 10770
rect 14410 10710 14430 10750
rect 14470 10710 14490 10750
rect 14410 10690 14490 10710
rect 14590 10750 14660 10770
rect 14590 10710 14610 10750
rect 14650 10710 14660 10750
rect 14590 10690 14660 10710
rect 11550 10630 11690 10650
rect 11550 10590 11560 10630
rect 11600 10590 11640 10630
rect 11680 10590 11690 10630
rect 11550 10530 11690 10590
rect 11550 10490 11560 10530
rect 11600 10490 11640 10530
rect 11680 10490 11690 10530
rect 11550 10430 11690 10490
rect 11550 10390 11560 10430
rect 11600 10390 11640 10430
rect 11680 10390 11690 10430
rect 11550 10330 11690 10390
rect 11550 10290 11560 10330
rect 11600 10290 11640 10330
rect 11680 10290 11690 10330
rect 11550 10230 11690 10290
rect 11550 10190 11560 10230
rect 11600 10190 11640 10230
rect 11680 10190 11690 10230
rect 11550 10130 11690 10190
rect 11550 10090 11560 10130
rect 11600 10090 11640 10130
rect 11680 10090 11690 10130
rect 11550 10070 11690 10090
rect 11810 10630 11870 10650
rect 11810 10590 11820 10630
rect 11860 10590 11870 10630
rect 11810 10530 11870 10590
rect 11810 10490 11820 10530
rect 11860 10490 11870 10530
rect 11810 10430 11870 10490
rect 11810 10390 11820 10430
rect 11860 10390 11870 10430
rect 11810 10330 11870 10390
rect 11810 10290 11820 10330
rect 11860 10290 11870 10330
rect 11810 10230 11870 10290
rect 11810 10190 11820 10230
rect 11860 10190 11870 10230
rect 11810 10130 11870 10190
rect 11810 10090 11820 10130
rect 11860 10090 11870 10130
rect 11810 10070 11870 10090
rect 11990 10630 12050 10650
rect 11990 10590 12000 10630
rect 12040 10590 12050 10630
rect 11990 10530 12050 10590
rect 11990 10490 12000 10530
rect 12040 10490 12050 10530
rect 11990 10430 12050 10490
rect 11990 10390 12000 10430
rect 12040 10390 12050 10430
rect 11990 10330 12050 10390
rect 11990 10290 12000 10330
rect 12040 10290 12050 10330
rect 11990 10230 12050 10290
rect 11990 10190 12000 10230
rect 12040 10190 12050 10230
rect 11990 10130 12050 10190
rect 11990 10090 12000 10130
rect 12040 10090 12050 10130
rect 11990 10070 12050 10090
rect 12170 10630 12230 10650
rect 12170 10590 12180 10630
rect 12220 10590 12230 10630
rect 12170 10530 12230 10590
rect 12170 10490 12180 10530
rect 12220 10490 12230 10530
rect 12170 10430 12230 10490
rect 12170 10390 12180 10430
rect 12220 10390 12230 10430
rect 12170 10330 12230 10390
rect 12170 10290 12180 10330
rect 12220 10290 12230 10330
rect 12170 10230 12230 10290
rect 12170 10190 12180 10230
rect 12220 10190 12230 10230
rect 12170 10130 12230 10190
rect 12170 10090 12180 10130
rect 12220 10090 12230 10130
rect 12170 10070 12230 10090
rect 12350 10630 12410 10650
rect 12350 10590 12360 10630
rect 12400 10590 12410 10630
rect 12350 10530 12410 10590
rect 12350 10490 12360 10530
rect 12400 10490 12410 10530
rect 12350 10430 12410 10490
rect 12350 10390 12360 10430
rect 12400 10390 12410 10430
rect 12350 10330 12410 10390
rect 12350 10290 12360 10330
rect 12400 10290 12410 10330
rect 12350 10230 12410 10290
rect 12350 10190 12360 10230
rect 12400 10190 12410 10230
rect 12350 10130 12410 10190
rect 12350 10090 12360 10130
rect 12400 10090 12410 10130
rect 12350 10070 12410 10090
rect 12530 10630 12590 10650
rect 12530 10590 12540 10630
rect 12580 10590 12590 10630
rect 12530 10530 12590 10590
rect 12530 10490 12540 10530
rect 12580 10490 12590 10530
rect 12530 10430 12590 10490
rect 12530 10390 12540 10430
rect 12580 10390 12590 10430
rect 12530 10330 12590 10390
rect 12530 10290 12540 10330
rect 12580 10290 12590 10330
rect 12530 10230 12590 10290
rect 12530 10190 12540 10230
rect 12580 10190 12590 10230
rect 12530 10130 12590 10190
rect 12530 10090 12540 10130
rect 12580 10090 12590 10130
rect 12530 10070 12590 10090
rect 12710 10630 12770 10650
rect 12710 10590 12720 10630
rect 12760 10590 12770 10630
rect 12710 10530 12770 10590
rect 12710 10490 12720 10530
rect 12760 10490 12770 10530
rect 12710 10430 12770 10490
rect 12710 10390 12720 10430
rect 12760 10390 12770 10430
rect 12710 10330 12770 10390
rect 12710 10290 12720 10330
rect 12760 10290 12770 10330
rect 12710 10230 12770 10290
rect 12710 10190 12720 10230
rect 12760 10190 12770 10230
rect 12710 10130 12770 10190
rect 12710 10090 12720 10130
rect 12760 10090 12770 10130
rect 12710 10070 12770 10090
rect 12890 10630 12950 10650
rect 12890 10590 12900 10630
rect 12940 10590 12950 10630
rect 12890 10530 12950 10590
rect 12890 10490 12900 10530
rect 12940 10490 12950 10530
rect 12890 10430 12950 10490
rect 12890 10390 12900 10430
rect 12940 10390 12950 10430
rect 12890 10330 12950 10390
rect 12890 10290 12900 10330
rect 12940 10290 12950 10330
rect 12890 10230 12950 10290
rect 12890 10190 12900 10230
rect 12940 10190 12950 10230
rect 12890 10130 12950 10190
rect 12890 10090 12900 10130
rect 12940 10090 12950 10130
rect 12890 10070 12950 10090
rect 13070 10630 13130 10650
rect 13070 10590 13080 10630
rect 13120 10590 13130 10630
rect 13070 10530 13130 10590
rect 13070 10490 13080 10530
rect 13120 10490 13130 10530
rect 13070 10430 13130 10490
rect 13070 10390 13080 10430
rect 13120 10390 13130 10430
rect 13070 10330 13130 10390
rect 13070 10290 13080 10330
rect 13120 10290 13130 10330
rect 13070 10230 13130 10290
rect 13070 10190 13080 10230
rect 13120 10190 13130 10230
rect 13070 10130 13130 10190
rect 13070 10090 13080 10130
rect 13120 10090 13130 10130
rect 13070 10070 13130 10090
rect 13250 10630 13310 10650
rect 13250 10590 13260 10630
rect 13300 10590 13310 10630
rect 13250 10530 13310 10590
rect 13250 10490 13260 10530
rect 13300 10490 13310 10530
rect 13250 10430 13310 10490
rect 13250 10390 13260 10430
rect 13300 10390 13310 10430
rect 13250 10330 13310 10390
rect 13250 10290 13260 10330
rect 13300 10290 13310 10330
rect 13250 10230 13310 10290
rect 13250 10190 13260 10230
rect 13300 10190 13310 10230
rect 13250 10130 13310 10190
rect 13250 10090 13260 10130
rect 13300 10090 13310 10130
rect 13250 10070 13310 10090
rect 13430 10630 13490 10650
rect 13430 10590 13440 10630
rect 13480 10590 13490 10630
rect 13430 10530 13490 10590
rect 13430 10490 13440 10530
rect 13480 10490 13490 10530
rect 13430 10430 13490 10490
rect 13430 10390 13440 10430
rect 13480 10390 13490 10430
rect 13430 10330 13490 10390
rect 13430 10290 13440 10330
rect 13480 10290 13490 10330
rect 13430 10230 13490 10290
rect 13430 10190 13440 10230
rect 13480 10190 13490 10230
rect 13430 10130 13490 10190
rect 13430 10090 13440 10130
rect 13480 10090 13490 10130
rect 13430 10070 13490 10090
rect 13610 10630 13670 10650
rect 13610 10590 13620 10630
rect 13660 10590 13670 10630
rect 13610 10530 13670 10590
rect 13610 10490 13620 10530
rect 13660 10490 13670 10530
rect 13610 10430 13670 10490
rect 13610 10390 13620 10430
rect 13660 10390 13670 10430
rect 13610 10330 13670 10390
rect 13610 10290 13620 10330
rect 13660 10290 13670 10330
rect 13610 10230 13670 10290
rect 13610 10190 13620 10230
rect 13660 10190 13670 10230
rect 13610 10130 13670 10190
rect 13610 10090 13620 10130
rect 13660 10090 13670 10130
rect 13610 10070 13670 10090
rect 13790 10630 13850 10650
rect 13790 10590 13800 10630
rect 13840 10590 13850 10630
rect 13790 10530 13850 10590
rect 13790 10490 13800 10530
rect 13840 10490 13850 10530
rect 13790 10430 13850 10490
rect 13790 10390 13800 10430
rect 13840 10390 13850 10430
rect 13790 10330 13850 10390
rect 13790 10290 13800 10330
rect 13840 10290 13850 10330
rect 13790 10230 13850 10290
rect 13790 10190 13800 10230
rect 13840 10190 13850 10230
rect 13790 10130 13850 10190
rect 13790 10090 13800 10130
rect 13840 10090 13850 10130
rect 13790 10070 13850 10090
rect 13970 10630 14030 10650
rect 13970 10590 13980 10630
rect 14020 10590 14030 10630
rect 13970 10530 14030 10590
rect 13970 10490 13980 10530
rect 14020 10490 14030 10530
rect 13970 10430 14030 10490
rect 13970 10390 13980 10430
rect 14020 10390 14030 10430
rect 13970 10330 14030 10390
rect 13970 10290 13980 10330
rect 14020 10290 14030 10330
rect 13970 10230 14030 10290
rect 13970 10190 13980 10230
rect 14020 10190 14030 10230
rect 13970 10130 14030 10190
rect 13970 10090 13980 10130
rect 14020 10090 14030 10130
rect 13970 10070 14030 10090
rect 14150 10630 14210 10650
rect 14150 10590 14160 10630
rect 14200 10590 14210 10630
rect 14150 10530 14210 10590
rect 14150 10490 14160 10530
rect 14200 10490 14210 10530
rect 14150 10430 14210 10490
rect 14150 10390 14160 10430
rect 14200 10390 14210 10430
rect 14150 10330 14210 10390
rect 14150 10290 14160 10330
rect 14200 10290 14210 10330
rect 14150 10230 14210 10290
rect 14150 10190 14160 10230
rect 14200 10190 14210 10230
rect 14150 10130 14210 10190
rect 14150 10090 14160 10130
rect 14200 10090 14210 10130
rect 14150 10070 14210 10090
rect 14330 10630 14390 10650
rect 14330 10590 14340 10630
rect 14380 10590 14390 10630
rect 14330 10530 14390 10590
rect 14330 10490 14340 10530
rect 14380 10490 14390 10530
rect 14330 10430 14390 10490
rect 14330 10390 14340 10430
rect 14380 10390 14390 10430
rect 14330 10330 14390 10390
rect 14330 10290 14340 10330
rect 14380 10290 14390 10330
rect 14330 10230 14390 10290
rect 14330 10190 14340 10230
rect 14380 10190 14390 10230
rect 14330 10130 14390 10190
rect 14330 10090 14340 10130
rect 14380 10090 14390 10130
rect 14330 10070 14390 10090
rect 14510 10630 14570 10650
rect 14510 10590 14520 10630
rect 14560 10590 14570 10630
rect 14510 10530 14570 10590
rect 14510 10490 14520 10530
rect 14560 10490 14570 10530
rect 14510 10430 14570 10490
rect 14510 10390 14520 10430
rect 14560 10390 14570 10430
rect 14510 10330 14570 10390
rect 14510 10290 14520 10330
rect 14560 10290 14570 10330
rect 14510 10230 14570 10290
rect 14510 10190 14520 10230
rect 14560 10190 14570 10230
rect 14510 10130 14570 10190
rect 14510 10090 14520 10130
rect 14560 10090 14570 10130
rect 14510 10070 14570 10090
rect 14690 10630 14750 10650
rect 14690 10590 14700 10630
rect 14740 10590 14750 10630
rect 14690 10530 14750 10590
rect 14690 10490 14700 10530
rect 14740 10490 14750 10530
rect 14690 10430 14750 10490
rect 14690 10390 14700 10430
rect 14740 10390 14750 10430
rect 14690 10330 14750 10390
rect 14690 10290 14700 10330
rect 14740 10290 14750 10330
rect 14690 10230 14750 10290
rect 14690 10190 14700 10230
rect 14740 10190 14750 10230
rect 14690 10130 14750 10190
rect 14690 10090 14700 10130
rect 14740 10090 14750 10130
rect 14690 10070 14750 10090
rect 14870 10630 15010 10650
rect 14870 10590 14880 10630
rect 14920 10590 14960 10630
rect 15000 10590 15010 10630
rect 14870 10530 15010 10590
rect 14870 10490 14880 10530
rect 14920 10490 14960 10530
rect 15000 10490 15010 10530
rect 15590 10550 15670 10570
rect 15590 10510 15610 10550
rect 15650 10510 15670 10550
rect 15590 10490 15670 10510
rect 15710 10550 15790 10570
rect 15710 10510 15730 10550
rect 15770 10510 15790 10550
rect 15710 10490 15790 10510
rect 15830 10550 15910 10570
rect 15830 10510 15850 10550
rect 15890 10510 15910 10550
rect 15830 10490 15910 10510
rect 14870 10430 15010 10490
rect 14870 10390 14880 10430
rect 14920 10390 14960 10430
rect 15000 10390 15010 10430
rect 14870 10330 15010 10390
rect 14870 10290 14880 10330
rect 14920 10290 14960 10330
rect 15000 10290 15010 10330
rect 14870 10230 15010 10290
rect 15410 10430 15560 10450
rect 15410 10390 15420 10430
rect 15460 10390 15510 10430
rect 15550 10390 15560 10430
rect 15410 10330 15560 10390
rect 15410 10290 15420 10330
rect 15460 10290 15510 10330
rect 15550 10290 15560 10330
rect 15410 10270 15560 10290
rect 15610 10430 15670 10450
rect 15610 10390 15620 10430
rect 15660 10390 15670 10430
rect 15610 10330 15670 10390
rect 15610 10290 15620 10330
rect 15660 10290 15670 10330
rect 15610 10270 15670 10290
rect 15720 10430 15780 10450
rect 15720 10390 15730 10430
rect 15770 10390 15780 10430
rect 15720 10330 15780 10390
rect 15720 10290 15730 10330
rect 15770 10290 15780 10330
rect 15720 10270 15780 10290
rect 15830 10430 15890 10450
rect 15830 10390 15840 10430
rect 15880 10390 15890 10430
rect 15830 10330 15890 10390
rect 15830 10290 15840 10330
rect 15880 10290 15890 10330
rect 15830 10270 15890 10290
rect 15940 10430 16080 10450
rect 15940 10390 15950 10430
rect 15990 10390 16030 10430
rect 16070 10390 16080 10430
rect 15940 10330 16080 10390
rect 15940 10290 15950 10330
rect 15990 10290 16030 10330
rect 16070 10290 16080 10330
rect 15940 10270 16080 10290
rect 14870 10190 14880 10230
rect 14920 10190 14960 10230
rect 15000 10190 15010 10230
rect 14870 10130 15010 10190
rect 15490 10210 15570 10230
rect 15490 10170 15510 10210
rect 15550 10170 15570 10210
rect 15490 10150 15570 10170
rect 15710 10210 15790 10230
rect 15710 10170 15730 10210
rect 15770 10170 15790 10210
rect 15710 10150 15790 10170
rect 15940 10210 16000 10230
rect 15940 10170 15950 10210
rect 15990 10170 16000 10210
rect 15940 10150 16000 10170
rect 14870 10090 14880 10130
rect 14920 10090 14960 10130
rect 15000 10090 15010 10130
rect 14870 10070 15010 10090
rect 11640 10030 11680 10070
rect 12000 10030 12040 10070
rect 12360 10030 12400 10070
rect 12720 10030 12760 10070
rect 13080 10030 13120 10070
rect 13440 10030 13480 10070
rect 13800 10030 13840 10070
rect 14160 10030 14200 10070
rect 14520 10030 14560 10070
rect 14880 10030 14920 10070
rect 11620 10010 11700 10030
rect 11620 9970 11640 10010
rect 11680 9970 11700 10010
rect 11620 9950 11700 9970
rect 11980 10010 12060 10030
rect 11980 9970 12000 10010
rect 12040 9970 12060 10010
rect 11980 9950 12060 9970
rect 12340 10010 12420 10030
rect 12340 9970 12360 10010
rect 12400 9970 12420 10010
rect 12340 9950 12420 9970
rect 12700 10010 12780 10030
rect 12700 9970 12720 10010
rect 12760 9970 12780 10010
rect 12700 9950 12780 9970
rect 13060 10010 13140 10030
rect 13060 9970 13080 10010
rect 13120 9970 13140 10010
rect 13060 9950 13140 9970
rect 13420 10010 13500 10030
rect 13420 9970 13440 10010
rect 13480 9970 13500 10010
rect 13420 9950 13500 9970
rect 13780 10010 13860 10030
rect 13780 9970 13800 10010
rect 13840 9970 13860 10010
rect 13780 9950 13860 9970
rect 14140 10010 14220 10030
rect 14140 9970 14160 10010
rect 14200 9970 14220 10010
rect 14140 9950 14220 9970
rect 14500 10010 14580 10030
rect 14500 9970 14520 10010
rect 14560 9970 14580 10010
rect 14500 9950 14580 9970
rect 14860 10010 14940 10030
rect 14860 9970 14880 10010
rect 14920 9970 14940 10010
rect 14860 9950 14940 9970
rect 11806 9742 11864 9760
rect 11806 9708 11818 9742
rect 11852 9708 11864 9742
rect 11806 9690 11864 9708
rect 11916 9742 11974 9760
rect 11916 9708 11928 9742
rect 11962 9708 11974 9742
rect 11916 9690 11974 9708
rect 12026 9742 12084 9760
rect 12026 9708 12038 9742
rect 12072 9708 12084 9742
rect 12026 9690 12084 9708
rect 12136 9742 12194 9760
rect 12136 9708 12148 9742
rect 12182 9708 12194 9742
rect 12136 9690 12194 9708
rect 12246 9742 12304 9760
rect 12246 9708 12258 9742
rect 12292 9708 12304 9742
rect 12246 9690 12304 9708
rect 12356 9742 12414 9760
rect 12356 9708 12368 9742
rect 12402 9708 12414 9742
rect 12356 9690 12414 9708
rect 12466 9742 12524 9760
rect 12466 9708 12478 9742
rect 12512 9708 12524 9742
rect 12466 9690 12524 9708
rect 12576 9742 12634 9760
rect 12576 9708 12588 9742
rect 12622 9708 12634 9742
rect 12576 9690 12634 9708
rect 12686 9742 12744 9760
rect 12686 9708 12698 9742
rect 12732 9708 12744 9742
rect 12686 9690 12744 9708
rect 12796 9742 12854 9760
rect 12796 9708 12808 9742
rect 12842 9708 12854 9742
rect 12796 9690 12854 9708
rect 13706 9742 13764 9760
rect 13706 9708 13718 9742
rect 13752 9708 13764 9742
rect 13706 9690 13764 9708
rect 13816 9742 13874 9760
rect 13816 9708 13828 9742
rect 13862 9708 13874 9742
rect 13816 9690 13874 9708
rect 13926 9742 13984 9760
rect 13926 9708 13938 9742
rect 13972 9708 13984 9742
rect 13926 9690 13984 9708
rect 14036 9742 14094 9760
rect 14036 9708 14048 9742
rect 14082 9708 14094 9742
rect 14036 9690 14094 9708
rect 14146 9742 14204 9760
rect 14146 9708 14158 9742
rect 14192 9708 14204 9742
rect 14146 9690 14204 9708
rect 14256 9742 14314 9760
rect 14256 9708 14268 9742
rect 14302 9708 14314 9742
rect 14256 9690 14314 9708
rect 14366 9742 14424 9760
rect 14366 9708 14378 9742
rect 14412 9708 14424 9742
rect 14366 9690 14424 9708
rect 14476 9742 14534 9760
rect 14476 9708 14488 9742
rect 14522 9708 14534 9742
rect 14476 9690 14534 9708
rect 14586 9742 14644 9760
rect 14586 9708 14598 9742
rect 14632 9708 14644 9742
rect 14586 9690 14644 9708
rect 14696 9742 14754 9760
rect 14696 9708 14708 9742
rect 14742 9708 14754 9742
rect 14696 9690 14754 9708
rect 11560 9630 11700 9650
rect 11560 9590 11570 9630
rect 11610 9590 11650 9630
rect 11690 9590 11700 9630
rect 11560 9530 11700 9590
rect 11560 9490 11570 9530
rect 11610 9490 11650 9530
rect 11690 9490 11700 9530
rect 11560 9470 11700 9490
rect 11750 9630 11810 9650
rect 11750 9590 11760 9630
rect 11800 9590 11810 9630
rect 11750 9530 11810 9590
rect 11750 9490 11760 9530
rect 11800 9490 11810 9530
rect 11750 9470 11810 9490
rect 11860 9630 11920 9650
rect 11860 9590 11870 9630
rect 11910 9590 11920 9630
rect 11860 9530 11920 9590
rect 11860 9490 11870 9530
rect 11910 9490 11920 9530
rect 11860 9470 11920 9490
rect 11970 9630 12030 9650
rect 11970 9590 11980 9630
rect 12020 9590 12030 9630
rect 11970 9530 12030 9590
rect 11970 9490 11980 9530
rect 12020 9490 12030 9530
rect 11970 9470 12030 9490
rect 12080 9630 12140 9650
rect 12080 9590 12090 9630
rect 12130 9590 12140 9630
rect 12080 9530 12140 9590
rect 12080 9490 12090 9530
rect 12130 9490 12140 9530
rect 12080 9470 12140 9490
rect 12190 9630 12250 9650
rect 12190 9590 12200 9630
rect 12240 9590 12250 9630
rect 12190 9530 12250 9590
rect 12190 9490 12200 9530
rect 12240 9490 12250 9530
rect 12190 9470 12250 9490
rect 12300 9630 12360 9650
rect 12300 9590 12310 9630
rect 12350 9590 12360 9630
rect 12300 9530 12360 9590
rect 12300 9490 12310 9530
rect 12350 9490 12360 9530
rect 12300 9470 12360 9490
rect 12410 9630 12470 9650
rect 12410 9590 12420 9630
rect 12460 9590 12470 9630
rect 12410 9530 12470 9590
rect 12410 9490 12420 9530
rect 12460 9490 12470 9530
rect 12410 9470 12470 9490
rect 12520 9630 12580 9650
rect 12520 9590 12530 9630
rect 12570 9590 12580 9630
rect 12520 9530 12580 9590
rect 12520 9490 12530 9530
rect 12570 9490 12580 9530
rect 12520 9470 12580 9490
rect 12630 9630 12690 9650
rect 12630 9590 12640 9630
rect 12680 9590 12690 9630
rect 12630 9530 12690 9590
rect 12630 9490 12640 9530
rect 12680 9490 12690 9530
rect 12630 9470 12690 9490
rect 12740 9630 12800 9650
rect 12740 9590 12750 9630
rect 12790 9590 12800 9630
rect 12740 9530 12800 9590
rect 12740 9490 12750 9530
rect 12790 9490 12800 9530
rect 12740 9470 12800 9490
rect 12850 9630 12910 9650
rect 12850 9590 12860 9630
rect 12900 9590 12910 9630
rect 12850 9530 12910 9590
rect 12850 9490 12860 9530
rect 12900 9490 12910 9530
rect 12850 9470 12910 9490
rect 12960 9630 13100 9650
rect 12960 9590 12970 9630
rect 13010 9590 13050 9630
rect 13090 9590 13100 9630
rect 12960 9530 13100 9590
rect 12960 9490 12970 9530
rect 13010 9490 13050 9530
rect 13090 9490 13100 9530
rect 12960 9470 13100 9490
rect 13460 9630 13600 9650
rect 13460 9590 13470 9630
rect 13510 9590 13550 9630
rect 13590 9590 13600 9630
rect 13460 9530 13600 9590
rect 13460 9490 13470 9530
rect 13510 9490 13550 9530
rect 13590 9490 13600 9530
rect 13460 9470 13600 9490
rect 13650 9630 13710 9650
rect 13650 9590 13660 9630
rect 13700 9590 13710 9630
rect 13650 9530 13710 9590
rect 13650 9490 13660 9530
rect 13700 9490 13710 9530
rect 13650 9470 13710 9490
rect 13760 9630 13820 9650
rect 13760 9590 13770 9630
rect 13810 9590 13820 9630
rect 13760 9530 13820 9590
rect 13760 9490 13770 9530
rect 13810 9490 13820 9530
rect 13760 9470 13820 9490
rect 13870 9630 13930 9650
rect 13870 9590 13880 9630
rect 13920 9590 13930 9630
rect 13870 9530 13930 9590
rect 13870 9490 13880 9530
rect 13920 9490 13930 9530
rect 13870 9470 13930 9490
rect 13980 9630 14040 9650
rect 13980 9590 13990 9630
rect 14030 9590 14040 9630
rect 13980 9530 14040 9590
rect 13980 9490 13990 9530
rect 14030 9490 14040 9530
rect 13980 9470 14040 9490
rect 14090 9630 14150 9650
rect 14090 9590 14100 9630
rect 14140 9590 14150 9630
rect 14090 9530 14150 9590
rect 14090 9490 14100 9530
rect 14140 9490 14150 9530
rect 14090 9470 14150 9490
rect 14200 9630 14260 9650
rect 14200 9590 14210 9630
rect 14250 9590 14260 9630
rect 14200 9530 14260 9590
rect 14200 9490 14210 9530
rect 14250 9490 14260 9530
rect 14200 9470 14260 9490
rect 14310 9630 14370 9650
rect 14310 9590 14320 9630
rect 14360 9590 14370 9630
rect 14310 9530 14370 9590
rect 14310 9490 14320 9530
rect 14360 9490 14370 9530
rect 14310 9470 14370 9490
rect 14420 9630 14480 9650
rect 14420 9590 14430 9630
rect 14470 9590 14480 9630
rect 14420 9530 14480 9590
rect 14420 9490 14430 9530
rect 14470 9490 14480 9530
rect 14420 9470 14480 9490
rect 14530 9630 14590 9650
rect 14530 9590 14540 9630
rect 14580 9590 14590 9630
rect 14530 9530 14590 9590
rect 14530 9490 14540 9530
rect 14580 9490 14590 9530
rect 14530 9470 14590 9490
rect 14640 9630 14700 9650
rect 14640 9590 14650 9630
rect 14690 9590 14700 9630
rect 14640 9530 14700 9590
rect 14640 9490 14650 9530
rect 14690 9490 14700 9530
rect 14640 9470 14700 9490
rect 14750 9630 14810 9650
rect 14750 9590 14760 9630
rect 14800 9590 14810 9630
rect 14750 9530 14810 9590
rect 14750 9490 14760 9530
rect 14800 9490 14810 9530
rect 14750 9470 14810 9490
rect 14860 9630 15000 9650
rect 14860 9590 14870 9630
rect 14910 9590 14950 9630
rect 14990 9590 15000 9630
rect 14860 9530 15000 9590
rect 14860 9490 14870 9530
rect 14910 9490 14950 9530
rect 14990 9490 15000 9530
rect 14860 9470 15000 9490
rect 11630 9410 11710 9430
rect 11630 9370 11650 9410
rect 11690 9370 11710 9410
rect 11630 9350 11710 9370
rect 12950 9410 13030 9430
rect 12950 9370 12970 9410
rect 13010 9370 13030 9410
rect 12950 9350 13030 9370
rect 13530 9410 13610 9430
rect 13530 9370 13550 9410
rect 13590 9370 13610 9410
rect 13530 9350 13610 9370
rect 14850 9410 14930 9430
rect 14850 9370 14870 9410
rect 14910 9370 14930 9410
rect 14850 9350 14930 9370
<< viali >>
rect 13260 19030 13300 19070
rect 13260 18950 13300 18990
rect 13260 18870 13300 18910
rect 8470 18597 8510 18610
rect 9260 18600 9300 18610
rect 8470 18570 8510 18597
rect 8470 18043 8508 18440
rect 8470 17234 8508 17631
rect 9260 18570 9300 18600
rect 10700 18597 10740 18610
rect 9250 18060 9290 18450
rect 9590 16836 9630 17226
rect 10700 18570 10740 18597
rect 10700 18050 10740 18440
rect 10370 16310 10410 16700
rect 11660 18392 11666 18414
rect 11666 18392 11694 18414
rect 11660 18380 11694 18392
rect 11760 18380 11794 18414
rect 11860 18380 11894 18414
rect 11960 18392 11992 18414
rect 11992 18392 11994 18414
rect 12060 18392 12082 18414
rect 12082 18392 12094 18414
rect 12160 18392 12172 18414
rect 12172 18392 12194 18414
rect 11960 18380 11994 18392
rect 12060 18380 12094 18392
rect 12160 18380 12194 18392
rect 11660 18302 11666 18314
rect 11666 18302 11694 18314
rect 11660 18280 11694 18302
rect 11760 18280 11794 18314
rect 11860 18280 11894 18314
rect 11960 18302 11992 18314
rect 11992 18302 11994 18314
rect 12060 18302 12082 18314
rect 12082 18302 12094 18314
rect 12160 18302 12172 18314
rect 12172 18302 12194 18314
rect 11960 18280 11994 18302
rect 12060 18280 12094 18302
rect 12160 18280 12194 18302
rect 11660 18212 11666 18214
rect 11666 18212 11694 18214
rect 11660 18180 11694 18212
rect 11760 18180 11794 18214
rect 11860 18180 11894 18214
rect 11960 18212 11992 18214
rect 11992 18212 11994 18214
rect 12060 18212 12082 18214
rect 12082 18212 12094 18214
rect 12160 18212 12172 18214
rect 12172 18212 12194 18214
rect 11960 18180 11994 18212
rect 12060 18180 12094 18212
rect 12160 18180 12194 18212
rect 11660 18080 11694 18114
rect 11760 18080 11794 18114
rect 11860 18080 11894 18114
rect 11960 18080 11994 18114
rect 12060 18080 12094 18114
rect 12160 18080 12194 18114
rect 11660 17980 11694 18014
rect 11760 17980 11794 18014
rect 11860 17980 11894 18014
rect 11960 17980 11994 18014
rect 12060 17980 12094 18014
rect 12160 17980 12194 18014
rect 11660 17886 11694 17914
rect 11660 17880 11666 17886
rect 11666 17880 11694 17886
rect 11760 17880 11794 17914
rect 11860 17880 11894 17914
rect 11960 17886 11994 17914
rect 12060 17886 12094 17914
rect 12160 17886 12194 17914
rect 11960 17880 11992 17886
rect 11992 17880 11994 17886
rect 12060 17880 12082 17886
rect 12082 17880 12094 17886
rect 12160 17880 12172 17886
rect 12172 17880 12194 17886
rect 13020 18392 13026 18414
rect 13026 18392 13054 18414
rect 13020 18380 13054 18392
rect 13120 18380 13154 18414
rect 13220 18380 13254 18414
rect 13320 18392 13352 18414
rect 13352 18392 13354 18414
rect 13420 18392 13442 18414
rect 13442 18392 13454 18414
rect 13520 18392 13532 18414
rect 13532 18392 13554 18414
rect 13320 18380 13354 18392
rect 13420 18380 13454 18392
rect 13520 18380 13554 18392
rect 13020 18302 13026 18314
rect 13026 18302 13054 18314
rect 13020 18280 13054 18302
rect 13120 18280 13154 18314
rect 13220 18280 13254 18314
rect 13320 18302 13352 18314
rect 13352 18302 13354 18314
rect 13420 18302 13442 18314
rect 13442 18302 13454 18314
rect 13520 18302 13532 18314
rect 13532 18302 13554 18314
rect 13320 18280 13354 18302
rect 13420 18280 13454 18302
rect 13520 18280 13554 18302
rect 13020 18212 13026 18214
rect 13026 18212 13054 18214
rect 13020 18180 13054 18212
rect 13120 18180 13154 18214
rect 13220 18180 13254 18214
rect 13320 18212 13352 18214
rect 13352 18212 13354 18214
rect 13420 18212 13442 18214
rect 13442 18212 13454 18214
rect 13520 18212 13532 18214
rect 13532 18212 13554 18214
rect 13320 18180 13354 18212
rect 13420 18180 13454 18212
rect 13520 18180 13554 18212
rect 13020 18080 13054 18114
rect 13120 18080 13154 18114
rect 13220 18080 13254 18114
rect 13320 18080 13354 18114
rect 13420 18080 13454 18114
rect 13520 18080 13554 18114
rect 13020 17980 13054 18014
rect 13120 17980 13154 18014
rect 13220 17980 13254 18014
rect 13320 17980 13354 18014
rect 13420 17980 13454 18014
rect 13520 17980 13554 18014
rect 13020 17886 13054 17914
rect 13020 17880 13026 17886
rect 13026 17880 13054 17886
rect 13120 17880 13154 17914
rect 13220 17880 13254 17914
rect 13320 17886 13354 17914
rect 13420 17886 13454 17914
rect 13520 17886 13554 17914
rect 13320 17880 13352 17886
rect 13352 17880 13354 17886
rect 13420 17880 13442 17886
rect 13442 17880 13454 17886
rect 13520 17880 13532 17886
rect 13532 17880 13554 17886
rect 14380 18392 14386 18414
rect 14386 18392 14414 18414
rect 14380 18380 14414 18392
rect 14480 18380 14514 18414
rect 14580 18380 14614 18414
rect 14680 18392 14712 18414
rect 14712 18392 14714 18414
rect 14780 18392 14802 18414
rect 14802 18392 14814 18414
rect 14880 18392 14892 18414
rect 14892 18392 14914 18414
rect 14680 18380 14714 18392
rect 14780 18380 14814 18392
rect 14880 18380 14914 18392
rect 14380 18302 14386 18314
rect 14386 18302 14414 18314
rect 14380 18280 14414 18302
rect 14480 18280 14514 18314
rect 14580 18280 14614 18314
rect 14680 18302 14712 18314
rect 14712 18302 14714 18314
rect 14780 18302 14802 18314
rect 14802 18302 14814 18314
rect 14880 18302 14892 18314
rect 14892 18302 14914 18314
rect 14680 18280 14714 18302
rect 14780 18280 14814 18302
rect 14880 18280 14914 18302
rect 14380 18212 14386 18214
rect 14386 18212 14414 18214
rect 14380 18180 14414 18212
rect 14480 18180 14514 18214
rect 14580 18180 14614 18214
rect 14680 18212 14712 18214
rect 14712 18212 14714 18214
rect 14780 18212 14802 18214
rect 14802 18212 14814 18214
rect 14880 18212 14892 18214
rect 14892 18212 14914 18214
rect 14680 18180 14714 18212
rect 14780 18180 14814 18212
rect 14880 18180 14914 18212
rect 14380 18080 14414 18114
rect 14480 18080 14514 18114
rect 14580 18080 14614 18114
rect 14680 18080 14714 18114
rect 14780 18080 14814 18114
rect 14880 18080 14914 18114
rect 14380 17980 14414 18014
rect 14480 17980 14514 18014
rect 14580 17980 14614 18014
rect 14680 17980 14714 18014
rect 14780 17980 14814 18014
rect 14880 17980 14914 18014
rect 14380 17886 14414 17914
rect 14380 17880 14386 17886
rect 14386 17880 14414 17886
rect 14480 17880 14514 17914
rect 14580 17880 14614 17914
rect 14680 17886 14714 17914
rect 14780 17886 14814 17914
rect 14880 17886 14914 17914
rect 14680 17880 14712 17886
rect 14712 17880 14714 17886
rect 14780 17880 14802 17886
rect 14802 17880 14814 17886
rect 14880 17880 14892 17886
rect 14892 17880 14914 17886
rect 15690 18597 15730 18610
rect 15690 18570 15730 18597
rect 16800 18594 16840 18610
rect 17590 18597 17630 18610
rect 11660 17032 11666 17054
rect 11666 17032 11694 17054
rect 11660 17020 11694 17032
rect 11760 17020 11794 17054
rect 11860 17020 11894 17054
rect 11960 17032 11992 17054
rect 11992 17032 11994 17054
rect 12060 17032 12082 17054
rect 12082 17032 12094 17054
rect 12160 17032 12172 17054
rect 12172 17032 12194 17054
rect 11960 17020 11994 17032
rect 12060 17020 12094 17032
rect 12160 17020 12194 17032
rect 11660 16942 11666 16954
rect 11666 16942 11694 16954
rect 11660 16920 11694 16942
rect 11760 16920 11794 16954
rect 11860 16920 11894 16954
rect 11960 16942 11992 16954
rect 11992 16942 11994 16954
rect 12060 16942 12082 16954
rect 12082 16942 12094 16954
rect 12160 16942 12172 16954
rect 12172 16942 12194 16954
rect 11960 16920 11994 16942
rect 12060 16920 12094 16942
rect 12160 16920 12194 16942
rect 11660 16852 11666 16854
rect 11666 16852 11694 16854
rect 11660 16820 11694 16852
rect 11760 16820 11794 16854
rect 11860 16820 11894 16854
rect 11960 16852 11992 16854
rect 11992 16852 11994 16854
rect 12060 16852 12082 16854
rect 12082 16852 12094 16854
rect 12160 16852 12172 16854
rect 12172 16852 12194 16854
rect 11960 16820 11994 16852
rect 12060 16820 12094 16852
rect 12160 16820 12194 16852
rect 11660 16720 11694 16754
rect 11760 16720 11794 16754
rect 11860 16720 11894 16754
rect 11960 16720 11994 16754
rect 12060 16720 12094 16754
rect 12160 16720 12194 16754
rect 11660 16620 11694 16654
rect 11760 16620 11794 16654
rect 11860 16620 11894 16654
rect 11960 16620 11994 16654
rect 12060 16620 12094 16654
rect 12160 16620 12194 16654
rect 11660 16526 11694 16554
rect 11660 16520 11666 16526
rect 11666 16520 11694 16526
rect 11760 16520 11794 16554
rect 11860 16520 11894 16554
rect 11960 16526 11994 16554
rect 12060 16526 12094 16554
rect 12160 16526 12194 16554
rect 11960 16520 11992 16526
rect 11992 16520 11994 16526
rect 12060 16520 12082 16526
rect 12082 16520 12094 16526
rect 12160 16520 12172 16526
rect 12172 16520 12194 16526
rect 13020 17032 13026 17054
rect 13026 17032 13054 17054
rect 13020 17020 13054 17032
rect 13120 17020 13154 17054
rect 13220 17020 13254 17054
rect 13320 17032 13352 17054
rect 13352 17032 13354 17054
rect 13420 17032 13442 17054
rect 13442 17032 13454 17054
rect 13520 17032 13532 17054
rect 13532 17032 13554 17054
rect 13320 17020 13354 17032
rect 13420 17020 13454 17032
rect 13520 17020 13554 17032
rect 13020 16942 13026 16954
rect 13026 16942 13054 16954
rect 13020 16920 13054 16942
rect 13120 16920 13154 16954
rect 13220 16920 13254 16954
rect 13320 16942 13352 16954
rect 13352 16942 13354 16954
rect 13420 16942 13442 16954
rect 13442 16942 13454 16954
rect 13520 16942 13532 16954
rect 13532 16942 13554 16954
rect 13320 16920 13354 16942
rect 13420 16920 13454 16942
rect 13520 16920 13554 16942
rect 13020 16852 13026 16854
rect 13026 16852 13054 16854
rect 13020 16820 13054 16852
rect 13120 16820 13154 16854
rect 13220 16820 13254 16854
rect 13320 16852 13352 16854
rect 13352 16852 13354 16854
rect 13420 16852 13442 16854
rect 13442 16852 13454 16854
rect 13520 16852 13532 16854
rect 13532 16852 13554 16854
rect 13320 16820 13354 16852
rect 13420 16820 13454 16852
rect 13520 16820 13554 16852
rect 13020 16720 13054 16754
rect 13120 16720 13154 16754
rect 13220 16720 13254 16754
rect 13320 16720 13354 16754
rect 13420 16720 13454 16754
rect 13520 16720 13554 16754
rect 13020 16620 13054 16654
rect 13120 16620 13154 16654
rect 13220 16620 13254 16654
rect 13320 16620 13354 16654
rect 13420 16620 13454 16654
rect 13520 16620 13554 16654
rect 13020 16526 13054 16554
rect 13020 16520 13026 16526
rect 13026 16520 13054 16526
rect 13120 16520 13154 16554
rect 13220 16520 13254 16554
rect 13320 16526 13354 16554
rect 13420 16526 13454 16554
rect 13520 16526 13554 16554
rect 13320 16520 13352 16526
rect 13352 16520 13354 16526
rect 13420 16520 13442 16526
rect 13442 16520 13454 16526
rect 13520 16520 13532 16526
rect 13532 16520 13554 16526
rect 14380 17032 14386 17054
rect 14386 17032 14414 17054
rect 14380 17020 14414 17032
rect 14480 17020 14514 17054
rect 14580 17020 14614 17054
rect 14680 17032 14712 17054
rect 14712 17032 14714 17054
rect 14780 17032 14802 17054
rect 14802 17032 14814 17054
rect 14880 17032 14892 17054
rect 14892 17032 14914 17054
rect 14680 17020 14714 17032
rect 14780 17020 14814 17032
rect 14880 17020 14914 17032
rect 14380 16942 14386 16954
rect 14386 16942 14414 16954
rect 14380 16920 14414 16942
rect 14480 16920 14514 16954
rect 14580 16920 14614 16954
rect 14680 16942 14712 16954
rect 14712 16942 14714 16954
rect 14780 16942 14802 16954
rect 14802 16942 14814 16954
rect 14880 16942 14892 16954
rect 14892 16942 14914 16954
rect 14680 16920 14714 16942
rect 14780 16920 14814 16942
rect 14880 16920 14914 16942
rect 14380 16852 14386 16854
rect 14386 16852 14414 16854
rect 14380 16820 14414 16852
rect 14480 16820 14514 16854
rect 14580 16820 14614 16854
rect 14680 16852 14712 16854
rect 14712 16852 14714 16854
rect 14780 16852 14802 16854
rect 14802 16852 14814 16854
rect 14880 16852 14892 16854
rect 14892 16852 14914 16854
rect 14680 16820 14714 16852
rect 14780 16820 14814 16852
rect 14880 16820 14914 16852
rect 14380 16720 14414 16754
rect 14480 16720 14514 16754
rect 14580 16720 14614 16754
rect 14680 16720 14714 16754
rect 14780 16720 14814 16754
rect 14880 16720 14914 16754
rect 14380 16620 14414 16654
rect 14480 16620 14514 16654
rect 14580 16620 14614 16654
rect 14680 16620 14714 16654
rect 14780 16620 14814 16654
rect 14880 16620 14914 16654
rect 14380 16526 14414 16554
rect 14380 16520 14386 16526
rect 14386 16520 14414 16526
rect 14480 16520 14514 16554
rect 14580 16520 14614 16554
rect 14680 16526 14714 16554
rect 14780 16526 14814 16554
rect 14880 16526 14914 16554
rect 14680 16520 14712 16526
rect 14712 16520 14714 16526
rect 14780 16520 14802 16526
rect 14802 16520 14814 16526
rect 14880 16520 14892 16526
rect 14892 16520 14914 16526
rect 15690 18050 15730 18440
rect 16020 16310 16060 16700
rect 16800 18570 16840 18594
rect 16803 18040 16841 18437
rect 16803 17441 16841 17838
rect 17590 18570 17630 18597
rect 17590 18043 17628 18440
rect 17590 17234 17628 17631
rect 11660 15672 11666 15694
rect 11666 15672 11694 15694
rect 11660 15660 11694 15672
rect 11760 15660 11794 15694
rect 11860 15660 11894 15694
rect 11960 15672 11992 15694
rect 11992 15672 11994 15694
rect 12060 15672 12082 15694
rect 12082 15672 12094 15694
rect 12160 15672 12172 15694
rect 12172 15672 12194 15694
rect 11960 15660 11994 15672
rect 12060 15660 12094 15672
rect 12160 15660 12194 15672
rect 11660 15582 11666 15594
rect 11666 15582 11694 15594
rect 11660 15560 11694 15582
rect 11760 15560 11794 15594
rect 11860 15560 11894 15594
rect 11960 15582 11992 15594
rect 11992 15582 11994 15594
rect 12060 15582 12082 15594
rect 12082 15582 12094 15594
rect 12160 15582 12172 15594
rect 12172 15582 12194 15594
rect 11960 15560 11994 15582
rect 12060 15560 12094 15582
rect 12160 15560 12194 15582
rect 11660 15492 11666 15494
rect 11666 15492 11694 15494
rect 11660 15460 11694 15492
rect 11760 15460 11794 15494
rect 11860 15460 11894 15494
rect 11960 15492 11992 15494
rect 11992 15492 11994 15494
rect 12060 15492 12082 15494
rect 12082 15492 12094 15494
rect 12160 15492 12172 15494
rect 12172 15492 12194 15494
rect 11960 15460 11994 15492
rect 12060 15460 12094 15492
rect 12160 15460 12194 15492
rect 11660 15360 11694 15394
rect 11760 15360 11794 15394
rect 11860 15360 11894 15394
rect 11960 15360 11994 15394
rect 12060 15360 12094 15394
rect 12160 15360 12194 15394
rect 11660 15260 11694 15294
rect 11760 15260 11794 15294
rect 11860 15260 11894 15294
rect 11960 15260 11994 15294
rect 12060 15260 12094 15294
rect 12160 15260 12194 15294
rect 11660 15166 11694 15194
rect 11660 15160 11666 15166
rect 11666 15160 11694 15166
rect 11760 15160 11794 15194
rect 11860 15160 11894 15194
rect 11960 15166 11994 15194
rect 12060 15166 12094 15194
rect 12160 15166 12194 15194
rect 11960 15160 11992 15166
rect 11992 15160 11994 15166
rect 12060 15160 12082 15166
rect 12082 15160 12094 15166
rect 12160 15160 12172 15166
rect 12172 15160 12194 15166
rect 13020 15672 13026 15694
rect 13026 15672 13054 15694
rect 13020 15660 13054 15672
rect 13120 15660 13154 15694
rect 13220 15660 13254 15694
rect 13320 15672 13352 15694
rect 13352 15672 13354 15694
rect 13420 15672 13442 15694
rect 13442 15672 13454 15694
rect 13520 15672 13532 15694
rect 13532 15672 13554 15694
rect 13320 15660 13354 15672
rect 13420 15660 13454 15672
rect 13520 15660 13554 15672
rect 13020 15582 13026 15594
rect 13026 15582 13054 15594
rect 13020 15560 13054 15582
rect 13120 15560 13154 15594
rect 13220 15560 13254 15594
rect 13320 15582 13352 15594
rect 13352 15582 13354 15594
rect 13420 15582 13442 15594
rect 13442 15582 13454 15594
rect 13520 15582 13532 15594
rect 13532 15582 13554 15594
rect 13320 15560 13354 15582
rect 13420 15560 13454 15582
rect 13520 15560 13554 15582
rect 13020 15492 13026 15494
rect 13026 15492 13054 15494
rect 13020 15460 13054 15492
rect 13120 15460 13154 15494
rect 13220 15460 13254 15494
rect 13320 15492 13352 15494
rect 13352 15492 13354 15494
rect 13420 15492 13442 15494
rect 13442 15492 13454 15494
rect 13520 15492 13532 15494
rect 13532 15492 13554 15494
rect 13320 15460 13354 15492
rect 13420 15460 13454 15492
rect 13520 15460 13554 15492
rect 13020 15360 13054 15394
rect 13120 15360 13154 15394
rect 13220 15360 13254 15394
rect 13320 15360 13354 15394
rect 13420 15360 13454 15394
rect 13520 15360 13554 15394
rect 13020 15260 13054 15294
rect 13120 15260 13154 15294
rect 13220 15260 13254 15294
rect 13320 15260 13354 15294
rect 13420 15260 13454 15294
rect 13520 15260 13554 15294
rect 13020 15166 13054 15194
rect 13020 15160 13026 15166
rect 13026 15160 13054 15166
rect 13120 15160 13154 15194
rect 13220 15160 13254 15194
rect 13320 15166 13354 15194
rect 13420 15166 13454 15194
rect 13520 15166 13554 15194
rect 13320 15160 13352 15166
rect 13352 15160 13354 15166
rect 13420 15160 13442 15166
rect 13442 15160 13454 15166
rect 13520 15160 13532 15166
rect 13532 15160 13554 15166
rect 14380 15672 14386 15694
rect 14386 15672 14414 15694
rect 14380 15660 14414 15672
rect 14480 15660 14514 15694
rect 14580 15660 14614 15694
rect 14680 15672 14712 15694
rect 14712 15672 14714 15694
rect 14780 15672 14802 15694
rect 14802 15672 14814 15694
rect 14880 15672 14892 15694
rect 14892 15672 14914 15694
rect 14680 15660 14714 15672
rect 14780 15660 14814 15672
rect 14880 15660 14914 15672
rect 14380 15582 14386 15594
rect 14386 15582 14414 15594
rect 14380 15560 14414 15582
rect 14480 15560 14514 15594
rect 14580 15560 14614 15594
rect 14680 15582 14712 15594
rect 14712 15582 14714 15594
rect 14780 15582 14802 15594
rect 14802 15582 14814 15594
rect 14880 15582 14892 15594
rect 14892 15582 14914 15594
rect 14680 15560 14714 15582
rect 14780 15560 14814 15582
rect 14880 15560 14914 15582
rect 14380 15492 14386 15494
rect 14386 15492 14414 15494
rect 14380 15460 14414 15492
rect 14480 15460 14514 15494
rect 14580 15460 14614 15494
rect 14680 15492 14712 15494
rect 14712 15492 14714 15494
rect 14780 15492 14802 15494
rect 14802 15492 14814 15494
rect 14880 15492 14892 15494
rect 14892 15492 14914 15494
rect 14680 15460 14714 15492
rect 14780 15460 14814 15492
rect 14880 15460 14914 15492
rect 14380 15360 14414 15394
rect 14480 15360 14514 15394
rect 14580 15360 14614 15394
rect 14680 15360 14714 15394
rect 14780 15360 14814 15394
rect 14880 15360 14914 15394
rect 14380 15260 14414 15294
rect 14480 15260 14514 15294
rect 14580 15260 14614 15294
rect 14680 15260 14714 15294
rect 14780 15260 14814 15294
rect 14880 15260 14914 15294
rect 14380 15166 14414 15194
rect 14380 15160 14386 15166
rect 14386 15160 14414 15166
rect 14480 15160 14514 15194
rect 14580 15160 14614 15194
rect 14680 15166 14714 15194
rect 14780 15166 14814 15194
rect 14880 15166 14914 15194
rect 14680 15160 14712 15166
rect 14712 15160 14714 15166
rect 14780 15160 14802 15166
rect 14802 15160 14814 15166
rect 14880 15160 14892 15166
rect 14892 15160 14914 15166
rect 12562 14550 12612 14600
rect 13960 14550 14010 14600
rect 11100 14160 11140 14200
rect 15490 14200 15530 14240
rect 15490 14120 15530 14160
rect 11180 13990 11220 14030
rect 11340 13990 11380 14030
rect 11500 13990 11540 14030
rect 11660 13990 11700 14030
rect 11820 13990 11860 14030
rect 11980 13990 12020 14030
rect 12140 13990 12180 14030
rect 12300 13990 12340 14030
rect 12460 13990 12500 14030
rect 12620 13990 12660 14030
rect 12780 13990 12820 14030
rect 12940 13990 12980 14030
rect 13100 13990 13140 14030
rect 13260 13990 13300 14030
rect 13420 13990 13460 14030
rect 13580 13990 13620 14030
rect 13740 13990 13780 14030
rect 13900 13990 13940 14030
rect 14060 13990 14100 14030
rect 14220 13990 14260 14030
rect 14380 13990 14420 14030
rect 14540 13990 14580 14030
rect 14700 13990 14740 14030
rect 14860 13990 14900 14030
rect 15020 13990 15060 14030
rect 15180 13990 15220 14030
rect 11920 13720 11960 13760
rect 14600 13720 14640 13760
rect 10760 13120 10800 13160
rect 10940 13080 10980 13120
rect 11180 13080 11220 13120
rect 11420 13080 11460 13120
rect 11660 13080 11700 13120
rect 12300 13080 12340 13120
rect 12540 13080 12580 13120
rect 12780 13080 12820 13120
rect 13080 13110 13120 13150
rect 15760 13600 15800 13640
rect 15760 13500 15800 13540
rect 15760 13400 15800 13440
rect 15760 13300 15800 13340
rect 15760 13200 15800 13240
rect 13440 13110 13480 13150
rect 13740 13080 13780 13120
rect 13980 13080 14020 13120
rect 14220 13080 14260 13120
rect 14860 13080 14900 13120
rect 15100 13080 15140 13120
rect 15340 13080 15380 13120
rect 15580 13080 15620 13120
rect 11443 12708 11477 12742
rect 11803 12708 11837 12742
rect 11923 12708 11957 12742
rect 12283 12708 12317 12742
rect 12403 12708 12437 12742
rect 12820 12680 12860 12720
rect 11380 12590 11420 12630
rect 11500 12590 11540 12630
rect 11620 12590 11660 12630
rect 11740 12590 11780 12630
rect 11860 12590 11900 12630
rect 11980 12590 12020 12630
rect 12100 12590 12140 12630
rect 12220 12590 12260 12630
rect 12340 12590 12380 12630
rect 12460 12590 12500 12630
rect 12580 12590 12620 12630
rect 12820 12600 12860 12640
rect 11544 12478 11578 12512
rect 11702 12478 11736 12512
rect 12026 12478 12060 12512
rect 12180 12478 12214 12512
rect 12504 12478 12538 12512
rect 12820 12520 12860 12560
rect 13700 12680 13740 12720
rect 14123 12708 14157 12742
rect 14243 12708 14277 12742
rect 14603 12708 14637 12742
rect 14723 12708 14757 12742
rect 15083 12708 15117 12742
rect 13700 12600 13740 12640
rect 13940 12590 13980 12630
rect 14060 12590 14100 12630
rect 14180 12590 14220 12630
rect 14300 12590 14340 12630
rect 14420 12590 14460 12630
rect 14540 12590 14580 12630
rect 14660 12590 14700 12630
rect 14780 12590 14820 12630
rect 14900 12590 14940 12630
rect 15020 12590 15060 12630
rect 15140 12590 15180 12630
rect 13700 12520 13740 12560
rect 14022 12478 14056 12512
rect 14346 12478 14380 12512
rect 14500 12478 14534 12512
rect 14824 12478 14858 12512
rect 14982 12478 15016 12512
rect 10720 11880 10760 11920
rect 10900 11870 10940 11910
rect 11380 11870 11420 11910
rect 11620 11870 11660 11910
rect 12100 11870 12140 11910
rect 12340 11870 12380 11910
rect 12760 11870 12800 11910
rect 13760 11870 13800 11910
rect 14180 11870 14220 11910
rect 14420 11870 14460 11910
rect 14900 11870 14940 11910
rect 15140 11870 15180 11910
rect 15620 11870 15660 11910
rect 15800 11880 15840 11920
rect 10540 11750 10580 11790
rect 10540 11650 10580 11690
rect 10660 11750 10700 11790
rect 10660 11650 10700 11690
rect 10780 11750 10820 11790
rect 10780 11650 10820 11690
rect 10900 11750 10940 11790
rect 10900 11650 10940 11690
rect 11020 11750 11060 11790
rect 11020 11650 11060 11690
rect 11140 11750 11180 11790
rect 11140 11650 11180 11690
rect 11260 11750 11300 11790
rect 11260 11650 11300 11690
rect 11380 11750 11420 11790
rect 11380 11650 11420 11690
rect 11500 11750 11540 11790
rect 11500 11650 11540 11690
rect 11620 11750 11660 11790
rect 11620 11650 11660 11690
rect 11740 11750 11780 11790
rect 11740 11650 11780 11690
rect 11860 11750 11900 11790
rect 11860 11650 11900 11690
rect 11980 11750 12020 11790
rect 11980 11650 12020 11690
rect 12100 11750 12140 11790
rect 12100 11650 12140 11690
rect 12220 11750 12260 11790
rect 12220 11650 12260 11690
rect 12340 11750 12380 11790
rect 12340 11650 12380 11690
rect 12460 11750 12500 11790
rect 12460 11650 12500 11690
rect 12580 11750 12620 11790
rect 12580 11650 12620 11690
rect 12700 11750 12740 11790
rect 12700 11650 12740 11690
rect 12820 11750 12860 11790
rect 12820 11650 12860 11690
rect 12940 11750 12980 11790
rect 12940 11650 12980 11690
rect 13580 11750 13620 11790
rect 13580 11650 13620 11690
rect 13700 11750 13740 11790
rect 13700 11650 13740 11690
rect 13820 11750 13860 11790
rect 13820 11650 13860 11690
rect 13940 11750 13980 11790
rect 13940 11650 13980 11690
rect 14060 11750 14100 11790
rect 14060 11650 14100 11690
rect 14180 11750 14220 11790
rect 14180 11650 14220 11690
rect 14300 11750 14340 11790
rect 14300 11650 14340 11690
rect 14420 11750 14460 11790
rect 14420 11650 14460 11690
rect 14540 11750 14580 11790
rect 14540 11650 14580 11690
rect 14660 11750 14700 11790
rect 14660 11650 14700 11690
rect 14780 11750 14820 11790
rect 14780 11650 14820 11690
rect 14900 11750 14940 11790
rect 14900 11650 14940 11690
rect 15020 11750 15060 11790
rect 15020 11650 15060 11690
rect 15140 11750 15180 11790
rect 15140 11650 15180 11690
rect 15260 11750 15300 11790
rect 15260 11650 15300 11690
rect 15380 11750 15420 11790
rect 15380 11650 15420 11690
rect 15500 11750 15540 11790
rect 15500 11650 15540 11690
rect 15620 11750 15660 11790
rect 15620 11650 15660 11690
rect 15740 11750 15780 11790
rect 15740 11650 15780 11690
rect 15860 11750 15900 11790
rect 15860 11650 15900 11690
rect 15980 11750 16020 11790
rect 15980 11650 16020 11690
rect 10540 11530 10580 11570
rect 12940 11530 12980 11570
rect 13580 11530 13620 11570
rect 15980 11530 16020 11570
rect 11910 10710 11950 10750
rect 12090 10710 12130 10750
rect 12270 10710 12310 10750
rect 12450 10710 12490 10750
rect 12630 10710 12670 10750
rect 12810 10710 12850 10750
rect 12990 10710 13030 10750
rect 13170 10710 13210 10750
rect 13350 10710 13390 10750
rect 13530 10710 13570 10750
rect 13710 10710 13750 10750
rect 13890 10710 13930 10750
rect 14070 10710 14110 10750
rect 14250 10710 14290 10750
rect 14430 10710 14470 10750
rect 14610 10710 14650 10750
rect 11640 10590 11680 10630
rect 11640 10490 11680 10530
rect 11640 10390 11680 10430
rect 11640 10290 11680 10330
rect 11640 10190 11680 10230
rect 11640 10090 11680 10130
rect 11820 10590 11860 10630
rect 11820 10490 11860 10530
rect 11820 10390 11860 10430
rect 11820 10290 11860 10330
rect 11820 10190 11860 10230
rect 11820 10090 11860 10130
rect 12000 10590 12040 10630
rect 12000 10490 12040 10530
rect 12000 10390 12040 10430
rect 12000 10290 12040 10330
rect 12000 10190 12040 10230
rect 12000 10090 12040 10130
rect 12180 10590 12220 10630
rect 12180 10490 12220 10530
rect 12180 10390 12220 10430
rect 12180 10290 12220 10330
rect 12180 10190 12220 10230
rect 12180 10090 12220 10130
rect 12360 10590 12400 10630
rect 12360 10490 12400 10530
rect 12360 10390 12400 10430
rect 12360 10290 12400 10330
rect 12360 10190 12400 10230
rect 12360 10090 12400 10130
rect 12540 10590 12580 10630
rect 12540 10490 12580 10530
rect 12540 10390 12580 10430
rect 12540 10290 12580 10330
rect 12540 10190 12580 10230
rect 12540 10090 12580 10130
rect 12720 10590 12760 10630
rect 12720 10490 12760 10530
rect 12720 10390 12760 10430
rect 12720 10290 12760 10330
rect 12720 10190 12760 10230
rect 12720 10090 12760 10130
rect 12900 10590 12940 10630
rect 12900 10490 12940 10530
rect 12900 10390 12940 10430
rect 12900 10290 12940 10330
rect 12900 10190 12940 10230
rect 12900 10090 12940 10130
rect 13080 10590 13120 10630
rect 13080 10490 13120 10530
rect 13080 10390 13120 10430
rect 13080 10290 13120 10330
rect 13080 10190 13120 10230
rect 13080 10090 13120 10130
rect 13260 10590 13300 10630
rect 13260 10490 13300 10530
rect 13260 10390 13300 10430
rect 13260 10290 13300 10330
rect 13260 10190 13300 10230
rect 13260 10090 13300 10130
rect 13440 10590 13480 10630
rect 13440 10490 13480 10530
rect 13440 10390 13480 10430
rect 13440 10290 13480 10330
rect 13440 10190 13480 10230
rect 13440 10090 13480 10130
rect 13620 10590 13660 10630
rect 13620 10490 13660 10530
rect 13620 10390 13660 10430
rect 13620 10290 13660 10330
rect 13620 10190 13660 10230
rect 13620 10090 13660 10130
rect 13800 10590 13840 10630
rect 13800 10490 13840 10530
rect 13800 10390 13840 10430
rect 13800 10290 13840 10330
rect 13800 10190 13840 10230
rect 13800 10090 13840 10130
rect 13980 10590 14020 10630
rect 13980 10490 14020 10530
rect 13980 10390 14020 10430
rect 13980 10290 14020 10330
rect 13980 10190 14020 10230
rect 13980 10090 14020 10130
rect 14160 10590 14200 10630
rect 14160 10490 14200 10530
rect 14160 10390 14200 10430
rect 14160 10290 14200 10330
rect 14160 10190 14200 10230
rect 14160 10090 14200 10130
rect 14340 10590 14380 10630
rect 14340 10490 14380 10530
rect 14340 10390 14380 10430
rect 14340 10290 14380 10330
rect 14340 10190 14380 10230
rect 14340 10090 14380 10130
rect 14520 10590 14560 10630
rect 14520 10490 14560 10530
rect 14520 10390 14560 10430
rect 14520 10290 14560 10330
rect 14520 10190 14560 10230
rect 14520 10090 14560 10130
rect 14700 10590 14740 10630
rect 14700 10490 14740 10530
rect 14700 10390 14740 10430
rect 14700 10290 14740 10330
rect 14700 10190 14740 10230
rect 14700 10090 14740 10130
rect 14880 10590 14920 10630
rect 14880 10490 14920 10530
rect 15610 10510 15650 10550
rect 15730 10510 15770 10550
rect 15850 10510 15890 10550
rect 14880 10390 14920 10430
rect 14880 10290 14920 10330
rect 15510 10390 15550 10430
rect 15510 10290 15550 10330
rect 15620 10390 15660 10430
rect 15620 10290 15660 10330
rect 15730 10390 15770 10430
rect 15730 10290 15770 10330
rect 15840 10390 15880 10430
rect 15840 10290 15880 10330
rect 15950 10390 15990 10430
rect 15950 10290 15990 10330
rect 14880 10190 14920 10230
rect 15510 10170 15550 10210
rect 15730 10170 15770 10210
rect 15950 10170 15990 10210
rect 14880 10090 14920 10130
rect 11640 9970 11680 10010
rect 12000 9970 12040 10010
rect 12360 9970 12400 10010
rect 12720 9970 12760 10010
rect 13080 9970 13120 10010
rect 13440 9970 13480 10010
rect 13800 9970 13840 10010
rect 14160 9970 14200 10010
rect 14520 9970 14560 10010
rect 14880 9970 14920 10010
rect 11818 9708 11852 9742
rect 11928 9708 11962 9742
rect 12038 9708 12072 9742
rect 12148 9708 12182 9742
rect 12258 9708 12292 9742
rect 12368 9708 12402 9742
rect 12478 9708 12512 9742
rect 12588 9708 12622 9742
rect 12698 9708 12732 9742
rect 12808 9708 12842 9742
rect 13718 9708 13752 9742
rect 13828 9708 13862 9742
rect 13938 9708 13972 9742
rect 14048 9708 14082 9742
rect 14158 9708 14192 9742
rect 14268 9708 14302 9742
rect 14378 9708 14412 9742
rect 14488 9708 14522 9742
rect 14598 9708 14632 9742
rect 14708 9708 14742 9742
rect 11570 9590 11610 9630
rect 11650 9590 11690 9630
rect 11570 9490 11610 9530
rect 11650 9490 11690 9530
rect 11760 9590 11800 9630
rect 11760 9490 11800 9530
rect 11870 9590 11910 9630
rect 11870 9490 11910 9530
rect 11980 9590 12020 9630
rect 11980 9490 12020 9530
rect 12090 9590 12130 9630
rect 12090 9490 12130 9530
rect 12200 9590 12240 9630
rect 12200 9490 12240 9530
rect 12310 9590 12350 9630
rect 12310 9490 12350 9530
rect 12420 9590 12460 9630
rect 12420 9490 12460 9530
rect 12530 9590 12570 9630
rect 12530 9490 12570 9530
rect 12640 9590 12680 9630
rect 12640 9490 12680 9530
rect 12750 9590 12790 9630
rect 12750 9490 12790 9530
rect 12860 9590 12900 9630
rect 12860 9490 12900 9530
rect 12970 9590 13010 9630
rect 13050 9590 13090 9630
rect 12970 9490 13010 9530
rect 13050 9490 13090 9530
rect 13470 9590 13510 9630
rect 13550 9590 13590 9630
rect 13470 9490 13510 9530
rect 13550 9490 13590 9530
rect 13660 9590 13700 9630
rect 13660 9490 13700 9530
rect 13770 9590 13810 9630
rect 13770 9490 13810 9530
rect 13880 9590 13920 9630
rect 13880 9490 13920 9530
rect 13990 9590 14030 9630
rect 13990 9490 14030 9530
rect 14100 9590 14140 9630
rect 14100 9490 14140 9530
rect 14210 9590 14250 9630
rect 14210 9490 14250 9530
rect 14320 9590 14360 9630
rect 14320 9490 14360 9530
rect 14430 9590 14470 9630
rect 14430 9490 14470 9530
rect 14540 9590 14580 9630
rect 14540 9490 14580 9530
rect 14650 9590 14690 9630
rect 14650 9490 14690 9530
rect 14760 9590 14800 9630
rect 14760 9490 14800 9530
rect 14870 9590 14910 9630
rect 14950 9590 14990 9630
rect 14870 9490 14910 9530
rect 14950 9490 14990 9530
rect 11650 9370 11690 9410
rect 12970 9370 13010 9410
rect 13550 9370 13590 9410
rect 14870 9370 14910 9410
<< metal1 >>
rect 8870 19190 8950 19200
rect 8870 19130 8880 19190
rect 8940 19130 8950 19190
rect 8450 19080 8530 19090
rect 8450 19020 8460 19080
rect 8520 19020 8530 19080
rect 8450 19000 8530 19020
rect 8450 18940 8460 19000
rect 8520 18940 8530 19000
rect 8450 18920 8530 18940
rect 8450 18860 8460 18920
rect 8520 18860 8530 18920
rect 8450 18610 8530 18860
rect 8450 18570 8470 18610
rect 8510 18570 8530 18610
rect 8450 18550 8530 18570
rect 8450 18440 8530 18460
rect 8450 18040 8460 18440
rect 8520 18040 8530 18440
rect 8450 18030 8530 18040
rect 8870 18450 8950 19130
rect 8870 18390 8880 18450
rect 8940 18390 8950 18450
rect 8870 18370 8950 18390
rect 8870 18310 8880 18370
rect 8940 18310 8950 18370
rect 8870 18280 8950 18310
rect 8870 18220 8880 18280
rect 8940 18220 8950 18280
rect 8870 18190 8950 18220
rect 8870 18130 8880 18190
rect 8940 18130 8950 18190
rect 8870 18110 8950 18130
rect 8870 18050 8880 18110
rect 8940 18050 8950 18110
rect 8870 18030 8950 18050
rect 9240 19080 9320 19090
rect 9240 19020 9250 19080
rect 9310 19020 9320 19080
rect 9240 19000 9320 19020
rect 9240 18940 9250 19000
rect 9310 18940 9320 19000
rect 9240 18920 9320 18940
rect 9240 18860 9250 18920
rect 9310 18860 9320 18920
rect 9240 18610 9320 18860
rect 9240 18570 9260 18610
rect 9300 18570 9320 18610
rect 9240 18450 9320 18570
rect 9240 18060 9250 18450
rect 9290 18060 9320 18450
rect 9240 18030 9320 18060
rect 10680 19080 10760 19090
rect 10680 19020 10690 19080
rect 10750 19020 10760 19080
rect 10680 19000 10760 19020
rect 10680 18940 10690 19000
rect 10750 18940 10760 19000
rect 10680 18920 10760 18940
rect 10680 18860 10690 18920
rect 10750 18860 10760 18920
rect 10680 18610 10760 18860
rect 10680 18570 10700 18610
rect 10740 18570 10760 18610
rect 10680 18440 10760 18570
rect 10680 18050 10700 18440
rect 10740 18050 10760 18440
rect 10680 18030 10760 18050
rect 8464 17631 8514 17643
rect 8464 17234 8470 17631
rect 8508 17234 8514 17631
rect 8464 17230 8514 17234
rect 8450 11580 8530 17230
rect 9570 17226 9650 17246
rect 9570 16836 9590 17226
rect 9630 16836 9650 17226
rect 8450 11520 8460 11580
rect 8520 11520 8530 11580
rect 8450 9760 8530 11520
rect 9460 14210 9540 14220
rect 9460 14150 9470 14210
rect 9530 14150 9540 14210
rect 9460 11090 9540 14150
rect 9570 12520 9650 16836
rect 10350 16700 10430 16720
rect 10350 16310 10370 16700
rect 10410 16310 10430 16700
rect 10350 14720 10430 16310
rect 10350 14660 10360 14720
rect 10420 14660 10430 14720
rect 10350 14650 10430 14660
rect 9570 12460 9580 12520
rect 9640 12460 9650 12520
rect 9570 11200 9650 12460
rect 9570 11140 9580 11200
rect 9640 11140 9650 11200
rect 9570 11130 9650 11140
rect 9680 14490 9760 14500
rect 9680 14430 9690 14490
rect 9750 14430 9760 14490
rect 9680 12750 9760 14430
rect 9680 12690 9690 12750
rect 9750 12690 9760 12750
rect 9460 11030 9470 11090
rect 9530 11030 9540 11090
rect 9460 11020 9540 11030
rect 8450 9700 8460 9760
rect 8520 9700 8530 9760
rect 8450 9690 8530 9700
rect 9680 9310 9760 12690
rect 10620 14380 10700 14390
rect 10620 14320 10630 14380
rect 10690 14320 10700 14380
rect 10620 12050 10700 14320
rect 11030 14380 11110 19200
rect 18190 19190 18270 19200
rect 18190 19130 18200 19190
rect 18260 19130 18270 19190
rect 13240 19080 13320 19090
rect 13240 19020 13250 19080
rect 13310 19020 13320 19080
rect 13240 19000 13320 19020
rect 13240 18940 13250 19000
rect 13310 18940 13320 19000
rect 13240 18920 13320 18940
rect 13240 18860 13250 18920
rect 13310 18860 13320 18920
rect 13240 18850 13320 18860
rect 15670 19080 15750 19090
rect 15670 19020 15680 19080
rect 15740 19020 15750 19080
rect 15670 19000 15750 19020
rect 15670 18940 15680 19000
rect 15740 18940 15750 19000
rect 15670 18920 15750 18940
rect 15670 18860 15680 18920
rect 15740 18860 15750 18920
rect 15670 18610 15750 18860
rect 15670 18570 15690 18610
rect 15730 18570 15750 18610
rect 11570 18414 14990 18490
rect 11570 18380 11660 18414
rect 11694 18380 11760 18414
rect 11794 18380 11860 18414
rect 11894 18380 11960 18414
rect 11994 18380 12060 18414
rect 12094 18380 12160 18414
rect 12194 18380 13020 18414
rect 13054 18380 13120 18414
rect 13154 18380 13220 18414
rect 13254 18380 13320 18414
rect 13354 18380 13420 18414
rect 13454 18380 13520 18414
rect 13554 18380 14380 18414
rect 14414 18380 14480 18414
rect 14514 18380 14580 18414
rect 14614 18380 14680 18414
rect 14714 18380 14780 18414
rect 14814 18380 14880 18414
rect 14914 18380 14990 18414
rect 11570 18314 14990 18380
rect 11570 18280 11660 18314
rect 11694 18280 11760 18314
rect 11794 18280 11860 18314
rect 11894 18280 11960 18314
rect 11994 18280 12060 18314
rect 12094 18280 12160 18314
rect 12194 18280 13020 18314
rect 13054 18280 13120 18314
rect 13154 18280 13220 18314
rect 13254 18280 13320 18314
rect 13354 18280 13420 18314
rect 13454 18280 13520 18314
rect 13554 18280 14380 18314
rect 14414 18280 14480 18314
rect 14514 18280 14580 18314
rect 14614 18280 14680 18314
rect 14714 18280 14780 18314
rect 14814 18280 14880 18314
rect 14914 18280 14990 18314
rect 11570 18214 14990 18280
rect 11570 18180 11660 18214
rect 11694 18180 11760 18214
rect 11794 18180 11860 18214
rect 11894 18180 11960 18214
rect 11994 18180 12060 18214
rect 12094 18180 12160 18214
rect 12194 18180 13020 18214
rect 13054 18180 13120 18214
rect 13154 18180 13220 18214
rect 13254 18180 13320 18214
rect 13354 18180 13420 18214
rect 13454 18180 13520 18214
rect 13554 18180 14380 18214
rect 14414 18180 14480 18214
rect 14514 18180 14580 18214
rect 14614 18180 14680 18214
rect 14714 18180 14780 18214
rect 14814 18180 14880 18214
rect 14914 18180 14990 18214
rect 11570 18114 14990 18180
rect 11570 18080 11660 18114
rect 11694 18080 11760 18114
rect 11794 18080 11860 18114
rect 11894 18080 11960 18114
rect 11994 18080 12060 18114
rect 12094 18080 12160 18114
rect 12194 18080 13020 18114
rect 13054 18080 13120 18114
rect 13154 18080 13220 18114
rect 13254 18080 13320 18114
rect 13354 18080 13420 18114
rect 13454 18080 13520 18114
rect 13554 18080 14380 18114
rect 14414 18080 14480 18114
rect 14514 18080 14580 18114
rect 14614 18080 14680 18114
rect 14714 18080 14780 18114
rect 14814 18080 14880 18114
rect 14914 18080 14990 18114
rect 11570 18014 14990 18080
rect 15670 18440 15750 18570
rect 15670 18050 15690 18440
rect 15730 18050 15750 18440
rect 15670 18030 15750 18050
rect 16780 19080 16860 19090
rect 16780 19020 16790 19080
rect 16850 19020 16860 19080
rect 16780 19000 16860 19020
rect 16780 18940 16790 19000
rect 16850 18940 16860 19000
rect 16780 18920 16860 18940
rect 16780 18860 16790 18920
rect 16850 18860 16860 18920
rect 16780 18610 16860 18860
rect 16780 18570 16800 18610
rect 16840 18570 16860 18610
rect 16780 18437 16860 18570
rect 17570 19080 17650 19090
rect 17570 19020 17580 19080
rect 17640 19020 17650 19080
rect 17570 19000 17650 19020
rect 17570 18940 17580 19000
rect 17640 18940 17650 19000
rect 17570 18920 17650 18940
rect 17570 18860 17580 18920
rect 17640 18860 17650 18920
rect 17570 18610 17650 18860
rect 18190 18850 18270 19130
rect 18190 18790 18200 18850
rect 18260 18790 18270 18850
rect 18190 18780 18270 18790
rect 17570 18570 17590 18610
rect 17630 18570 17650 18610
rect 17570 18550 17650 18570
rect 16780 18040 16803 18437
rect 16841 18040 16860 18437
rect 16780 18030 16860 18040
rect 17570 18440 17650 18460
rect 17570 18040 17580 18440
rect 17640 18040 17650 18440
rect 17570 18030 17650 18040
rect 17950 18450 18030 18460
rect 17950 18390 17960 18450
rect 18020 18390 18030 18450
rect 17950 18370 18030 18390
rect 17950 18310 17960 18370
rect 18020 18310 18030 18370
rect 17950 18280 18030 18310
rect 17950 18220 17960 18280
rect 18020 18220 18030 18280
rect 17950 18190 18030 18220
rect 17950 18130 17960 18190
rect 18020 18130 18030 18190
rect 17950 18110 18030 18130
rect 17950 18050 17960 18110
rect 18020 18050 18030 18110
rect 18640 18150 18740 18170
rect 18640 18090 18660 18150
rect 18720 18090 18740 18150
rect 18640 18070 18740 18090
rect 16797 18028 16847 18030
rect 11570 17980 11660 18014
rect 11694 17980 11760 18014
rect 11794 17980 11860 18014
rect 11894 17980 11960 18014
rect 11994 17980 12060 18014
rect 12094 17980 12160 18014
rect 12194 17980 13020 18014
rect 13054 17980 13120 18014
rect 13154 17980 13220 18014
rect 13254 17980 13320 18014
rect 13354 17980 13420 18014
rect 13454 17980 13520 18014
rect 13554 17980 14380 18014
rect 14414 17980 14480 18014
rect 14514 17980 14580 18014
rect 14614 17980 14680 18014
rect 14714 17980 14780 18014
rect 14814 17980 14880 18014
rect 14914 17980 14990 18014
rect 11570 17914 14990 17980
rect 11570 17880 11660 17914
rect 11694 17880 11760 17914
rect 11794 17880 11860 17914
rect 11894 17880 11960 17914
rect 11994 17880 12060 17914
rect 12094 17880 12160 17914
rect 12194 17880 13020 17914
rect 13054 17880 13120 17914
rect 13154 17880 13220 17914
rect 13254 17880 13320 17914
rect 13354 17880 13420 17914
rect 13454 17880 13520 17914
rect 13554 17880 14380 17914
rect 14414 17880 14480 17914
rect 14514 17880 14580 17914
rect 14614 17880 14680 17914
rect 14714 17880 14780 17914
rect 14814 17880 14880 17914
rect 14914 17880 14990 17914
rect 11570 17790 14990 17880
rect 11570 17054 12270 17790
rect 11570 17020 11660 17054
rect 11694 17020 11760 17054
rect 11794 17020 11860 17054
rect 11894 17020 11960 17054
rect 11994 17020 12060 17054
rect 12094 17020 12160 17054
rect 12194 17020 12270 17054
rect 11570 16954 12270 17020
rect 11570 16920 11660 16954
rect 11694 16920 11760 16954
rect 11794 16920 11860 16954
rect 11894 16920 11960 16954
rect 11994 16920 12060 16954
rect 12094 16920 12160 16954
rect 12194 16920 12270 16954
rect 11570 16854 12270 16920
rect 11570 16820 11660 16854
rect 11694 16820 11760 16854
rect 11794 16820 11860 16854
rect 11894 16820 11960 16854
rect 11994 16820 12060 16854
rect 12094 16820 12160 16854
rect 12194 16820 12270 16854
rect 11140 16810 11220 16820
rect 11140 16750 11150 16810
rect 11210 16750 11220 16810
rect 11140 14610 11220 16750
rect 11570 16810 12270 16820
rect 11570 16750 11580 16810
rect 11640 16754 12270 16810
rect 11640 16750 11660 16754
rect 11570 16720 11660 16750
rect 11694 16720 11760 16754
rect 11794 16720 11860 16754
rect 11894 16720 11960 16754
rect 11994 16720 12060 16754
rect 12094 16720 12160 16754
rect 12194 16720 12270 16754
rect 11570 16654 12270 16720
rect 11570 16620 11660 16654
rect 11694 16620 11760 16654
rect 11794 16620 11860 16654
rect 11894 16620 11960 16654
rect 11994 16620 12060 16654
rect 12094 16620 12160 16654
rect 12194 16620 12270 16654
rect 11570 16554 12270 16620
rect 11570 16520 11660 16554
rect 11694 16520 11760 16554
rect 11794 16520 11860 16554
rect 11894 16520 11960 16554
rect 11994 16520 12060 16554
rect 12094 16520 12160 16554
rect 12194 16520 12270 16554
rect 11570 15770 12270 16520
rect 12930 17054 13630 17130
rect 12930 17020 13020 17054
rect 13054 17020 13120 17054
rect 13154 17020 13220 17054
rect 13254 17020 13320 17054
rect 13354 17020 13420 17054
rect 13454 17020 13520 17054
rect 13554 17020 13630 17054
rect 12930 16954 13630 17020
rect 12930 16920 13020 16954
rect 13054 16920 13120 16954
rect 13154 16920 13220 16954
rect 13254 16920 13320 16954
rect 13354 16920 13420 16954
rect 13454 16920 13520 16954
rect 13554 16920 13630 16954
rect 12930 16854 13630 16920
rect 12930 16820 13020 16854
rect 13054 16820 13120 16854
rect 13154 16820 13220 16854
rect 13254 16820 13320 16854
rect 13354 16820 13420 16854
rect 13454 16820 13520 16854
rect 13554 16820 13630 16854
rect 12930 16810 13630 16820
rect 12930 16754 13250 16810
rect 13310 16754 13630 16810
rect 12930 16720 13020 16754
rect 13054 16720 13120 16754
rect 13154 16720 13220 16754
rect 13310 16750 13320 16754
rect 13254 16720 13320 16750
rect 13354 16720 13420 16754
rect 13454 16720 13520 16754
rect 13554 16720 13630 16754
rect 12930 16654 13630 16720
rect 12930 16620 13020 16654
rect 13054 16620 13120 16654
rect 13154 16620 13220 16654
rect 13254 16620 13320 16654
rect 13354 16620 13420 16654
rect 13454 16620 13520 16654
rect 13554 16620 13630 16654
rect 12930 16554 13630 16620
rect 12930 16520 13020 16554
rect 13054 16520 13120 16554
rect 13154 16520 13220 16554
rect 13254 16520 13320 16554
rect 13354 16520 13420 16554
rect 13454 16520 13520 16554
rect 13554 16520 13630 16554
rect 12930 16430 13630 16520
rect 14290 17054 14990 17790
rect 14290 17020 14380 17054
rect 14414 17020 14480 17054
rect 14514 17020 14580 17054
rect 14614 17020 14680 17054
rect 14714 17020 14780 17054
rect 14814 17020 14880 17054
rect 14914 17020 14990 17054
rect 14290 16954 14990 17020
rect 14290 16920 14380 16954
rect 14414 16920 14480 16954
rect 14514 16920 14580 16954
rect 14614 16920 14680 16954
rect 14714 16920 14780 16954
rect 14814 16920 14880 16954
rect 14914 16920 14990 16954
rect 14290 16854 14990 16920
rect 14290 16820 14380 16854
rect 14414 16820 14480 16854
rect 14514 16820 14580 16854
rect 14614 16820 14680 16854
rect 14714 16820 14780 16854
rect 14814 16820 14880 16854
rect 14914 16820 14990 16854
rect 16780 17838 16860 17850
rect 16780 17441 16803 17838
rect 16841 17441 16860 17838
rect 14290 16754 14990 16820
rect 14290 16720 14380 16754
rect 14414 16720 14480 16754
rect 14514 16720 14580 16754
rect 14614 16720 14680 16754
rect 14714 16720 14780 16754
rect 14814 16720 14880 16754
rect 14914 16720 14990 16754
rect 14290 16654 14990 16720
rect 14290 16620 14380 16654
rect 14414 16620 14480 16654
rect 14514 16620 14580 16654
rect 14614 16620 14680 16654
rect 14714 16620 14780 16654
rect 14814 16620 14880 16654
rect 14914 16620 14990 16654
rect 14290 16554 14990 16620
rect 14290 16520 14380 16554
rect 14414 16520 14480 16554
rect 14514 16520 14580 16554
rect 14614 16520 14680 16554
rect 14714 16520 14780 16554
rect 14814 16520 14880 16554
rect 14914 16520 14990 16554
rect 14290 15770 14990 16520
rect 11570 15694 14990 15770
rect 11570 15660 11660 15694
rect 11694 15660 11760 15694
rect 11794 15660 11860 15694
rect 11894 15660 11960 15694
rect 11994 15660 12060 15694
rect 12094 15660 12160 15694
rect 12194 15660 13020 15694
rect 13054 15660 13120 15694
rect 13154 15660 13220 15694
rect 13254 15660 13320 15694
rect 13354 15660 13420 15694
rect 13454 15660 13520 15694
rect 13554 15660 14380 15694
rect 14414 15660 14480 15694
rect 14514 15660 14580 15694
rect 14614 15660 14680 15694
rect 14714 15660 14780 15694
rect 14814 15660 14880 15694
rect 14914 15660 14990 15694
rect 11570 15594 14990 15660
rect 11570 15560 11660 15594
rect 11694 15560 11760 15594
rect 11794 15560 11860 15594
rect 11894 15560 11960 15594
rect 11994 15560 12060 15594
rect 12094 15560 12160 15594
rect 12194 15560 13020 15594
rect 13054 15560 13120 15594
rect 13154 15560 13220 15594
rect 13254 15560 13320 15594
rect 13354 15560 13420 15594
rect 13454 15560 13520 15594
rect 13554 15560 14380 15594
rect 14414 15560 14480 15594
rect 14514 15560 14580 15594
rect 14614 15560 14680 15594
rect 14714 15560 14780 15594
rect 14814 15560 14880 15594
rect 14914 15560 14990 15594
rect 11570 15494 14990 15560
rect 11570 15460 11660 15494
rect 11694 15460 11760 15494
rect 11794 15460 11860 15494
rect 11894 15460 11960 15494
rect 11994 15460 12060 15494
rect 12094 15460 12160 15494
rect 12194 15460 13020 15494
rect 13054 15460 13120 15494
rect 13154 15460 13220 15494
rect 13254 15460 13320 15494
rect 13354 15460 13420 15494
rect 13454 15460 13520 15494
rect 13554 15460 14380 15494
rect 14414 15460 14480 15494
rect 14514 15460 14580 15494
rect 14614 15460 14680 15494
rect 14714 15460 14780 15494
rect 14814 15460 14880 15494
rect 14914 15460 14990 15494
rect 11570 15394 14990 15460
rect 11570 15360 11660 15394
rect 11694 15360 11760 15394
rect 11794 15360 11860 15394
rect 11894 15360 11960 15394
rect 11994 15360 12060 15394
rect 12094 15360 12160 15394
rect 12194 15360 13020 15394
rect 13054 15360 13120 15394
rect 13154 15360 13220 15394
rect 13254 15360 13320 15394
rect 13354 15360 13420 15394
rect 13454 15360 13520 15394
rect 13554 15360 14380 15394
rect 14414 15360 14480 15394
rect 14514 15360 14580 15394
rect 14614 15360 14680 15394
rect 14714 15360 14780 15394
rect 14814 15360 14880 15394
rect 14914 15360 14990 15394
rect 11570 15294 14990 15360
rect 11570 15260 11660 15294
rect 11694 15260 11760 15294
rect 11794 15260 11860 15294
rect 11894 15260 11960 15294
rect 11994 15260 12060 15294
rect 12094 15260 12160 15294
rect 12194 15260 13020 15294
rect 13054 15260 13120 15294
rect 13154 15260 13220 15294
rect 13254 15260 13320 15294
rect 13354 15260 13420 15294
rect 13454 15260 13520 15294
rect 13554 15260 14380 15294
rect 14414 15260 14480 15294
rect 14514 15260 14580 15294
rect 14614 15260 14680 15294
rect 14714 15260 14780 15294
rect 14814 15260 14880 15294
rect 14914 15260 14990 15294
rect 11570 15194 14990 15260
rect 11570 15160 11660 15194
rect 11694 15160 11760 15194
rect 11794 15160 11860 15194
rect 11894 15160 11960 15194
rect 11994 15160 12060 15194
rect 12094 15160 12160 15194
rect 12194 15160 13020 15194
rect 13054 15160 13120 15194
rect 13154 15160 13220 15194
rect 13254 15160 13320 15194
rect 13354 15160 13420 15194
rect 13454 15160 13520 15194
rect 13554 15160 14380 15194
rect 14414 15160 14480 15194
rect 14514 15160 14580 15194
rect 14614 15160 14680 15194
rect 14714 15160 14780 15194
rect 14814 15160 14880 15194
rect 14914 15160 14990 15194
rect 11570 15070 14990 15160
rect 15340 16810 15420 16820
rect 15340 16750 15350 16810
rect 15410 16750 15420 16810
rect 15340 14800 15420 16750
rect 15340 14740 15350 14800
rect 15410 14740 15420 14800
rect 15340 14730 15420 14740
rect 16000 16700 16080 16720
rect 16000 16310 16020 16700
rect 16060 16310 16080 16700
rect 16000 14800 16080 16310
rect 16350 15350 16590 15370
rect 16350 15290 16360 15350
rect 16420 15290 16440 15350
rect 16500 15290 16520 15350
rect 16580 15290 16590 15350
rect 16000 14740 16010 14800
rect 16070 14740 16080 14800
rect 16000 14730 16080 14740
rect 16240 14800 16320 14810
rect 16240 14740 16250 14800
rect 16310 14740 16320 14800
rect 16240 14730 16320 14740
rect 13950 14720 14030 14730
rect 13950 14660 13960 14720
rect 14020 14660 14030 14720
rect 13950 14610 14030 14660
rect 11140 14550 11150 14610
rect 11210 14550 11220 14610
rect 11140 14540 11220 14550
rect 12542 14540 12552 14610
rect 12622 14540 12632 14610
rect 13940 14540 13950 14610
rect 14020 14540 14030 14610
rect 16150 14600 16230 14610
rect 16150 14540 16160 14600
rect 16220 14540 16230 14600
rect 16150 14530 16230 14540
rect 11030 14320 11040 14380
rect 11100 14320 11110 14380
rect 11030 14310 11110 14320
rect 15470 14250 15550 14260
rect 11080 14210 11160 14220
rect 11080 14150 11090 14210
rect 11150 14150 11160 14210
rect 11080 14140 11160 14150
rect 15470 14190 15480 14250
rect 15540 14190 15550 14250
rect 15470 14170 15550 14190
rect 15470 14110 15480 14170
rect 15540 14110 15550 14170
rect 15470 14100 15550 14110
rect 11160 14040 11240 14050
rect 11160 13980 11170 14040
rect 11230 13980 11240 14040
rect 11160 13970 11240 13980
rect 11320 14040 11400 14050
rect 11320 13980 11330 14040
rect 11390 13980 11400 14040
rect 11320 13970 11400 13980
rect 11480 14040 11560 14050
rect 11480 13980 11490 14040
rect 11550 13980 11560 14040
rect 11480 13970 11560 13980
rect 11640 14040 11720 14050
rect 11640 13980 11650 14040
rect 11710 13980 11720 14040
rect 11640 13970 11720 13980
rect 11800 14040 11880 14050
rect 11800 13980 11810 14040
rect 11870 13980 11880 14040
rect 11800 13970 11880 13980
rect 11960 14040 12040 14050
rect 11960 13980 11970 14040
rect 12030 13980 12040 14040
rect 11960 13970 12040 13980
rect 12120 14040 12200 14050
rect 12120 13980 12130 14040
rect 12190 13980 12200 14040
rect 12120 13970 12200 13980
rect 12280 14040 12360 14050
rect 12280 13980 12290 14040
rect 12350 13980 12360 14040
rect 12280 13970 12360 13980
rect 12440 14040 12520 14050
rect 12440 13980 12450 14040
rect 12510 13980 12520 14040
rect 12440 13970 12520 13980
rect 12600 14040 12680 14050
rect 12600 13980 12610 14040
rect 12670 13980 12680 14040
rect 12600 13970 12680 13980
rect 12760 14040 12840 14050
rect 12760 13980 12770 14040
rect 12830 13980 12840 14040
rect 12760 13970 12840 13980
rect 12920 14040 13000 14050
rect 12920 13980 12930 14040
rect 12990 13980 13000 14040
rect 12920 13970 13000 13980
rect 13080 14040 13160 14050
rect 13080 13980 13090 14040
rect 13150 13980 13160 14040
rect 13080 13970 13160 13980
rect 13240 14040 13320 14050
rect 13240 13980 13250 14040
rect 13310 13980 13320 14040
rect 13240 13970 13320 13980
rect 13400 14040 13480 14050
rect 13400 13980 13410 14040
rect 13470 13980 13480 14040
rect 13400 13970 13480 13980
rect 13560 14040 13640 14050
rect 13560 13980 13570 14040
rect 13630 13980 13640 14040
rect 13560 13970 13640 13980
rect 13720 14040 13800 14050
rect 13720 13980 13730 14040
rect 13790 13980 13800 14040
rect 13720 13970 13800 13980
rect 13880 14040 13960 14050
rect 13880 13980 13890 14040
rect 13950 13980 13960 14040
rect 13880 13970 13960 13980
rect 14040 14040 14120 14050
rect 14040 13980 14050 14040
rect 14110 13980 14120 14040
rect 14040 13970 14120 13980
rect 14200 14040 14280 14050
rect 14200 13980 14210 14040
rect 14270 13980 14280 14040
rect 14200 13970 14280 13980
rect 14360 14040 14440 14050
rect 14360 13980 14370 14040
rect 14430 13980 14440 14040
rect 14360 13970 14440 13980
rect 14520 14040 14600 14050
rect 14520 13980 14530 14040
rect 14590 13980 14600 14040
rect 14520 13970 14600 13980
rect 14680 14040 14760 14050
rect 14680 13980 14690 14040
rect 14750 13980 14760 14040
rect 14680 13970 14760 13980
rect 14840 14040 14920 14050
rect 14840 13980 14850 14040
rect 14910 13980 14920 14040
rect 14840 13970 14920 13980
rect 15000 14040 15080 14050
rect 15000 13980 15010 14040
rect 15070 13980 15080 14040
rect 15000 13970 15080 13980
rect 15160 14040 15240 14050
rect 15160 13980 15170 14040
rect 15230 13980 15240 14040
rect 15160 13970 15240 13980
rect 11900 13930 11980 13940
rect 11900 13870 11910 13930
rect 11970 13870 11980 13930
rect 11900 13850 11980 13870
rect 11900 13790 11910 13850
rect 11970 13790 11980 13850
rect 11900 13770 11980 13790
rect 11900 13710 11910 13770
rect 11970 13710 11980 13770
rect 11900 13700 11980 13710
rect 13160 13930 13400 13940
rect 13160 13870 13170 13930
rect 13230 13870 13250 13930
rect 13310 13870 13330 13930
rect 13390 13870 13400 13930
rect 13160 13850 13400 13870
rect 13160 13790 13170 13850
rect 13230 13790 13250 13850
rect 13310 13790 13330 13850
rect 13390 13790 13400 13850
rect 13160 13770 13400 13790
rect 13160 13710 13170 13770
rect 13230 13710 13250 13770
rect 13310 13710 13330 13770
rect 13390 13710 13400 13770
rect 10740 13160 10820 13180
rect 10740 13120 10760 13160
rect 10800 13120 10820 13160
rect 13070 13150 13130 13170
rect 10740 12860 10820 13120
rect 10920 13130 11000 13140
rect 10920 13070 10930 13130
rect 10990 13070 11000 13130
rect 10920 13050 11000 13070
rect 10920 12990 10930 13050
rect 10990 12990 11000 13050
rect 10920 12970 11000 12990
rect 10920 12910 10930 12970
rect 10990 12910 11000 12970
rect 10920 12900 11000 12910
rect 11160 13130 11240 13140
rect 11160 13070 11170 13130
rect 11230 13070 11240 13130
rect 11160 13050 11240 13070
rect 11160 12990 11170 13050
rect 11230 12990 11240 13050
rect 11160 12970 11240 12990
rect 11160 12910 11170 12970
rect 11230 12910 11240 12970
rect 11160 12900 11240 12910
rect 11400 13130 11480 13140
rect 11400 13070 11410 13130
rect 11470 13070 11480 13130
rect 11400 13050 11480 13070
rect 11400 12990 11410 13050
rect 11470 12990 11480 13050
rect 11400 12970 11480 12990
rect 11400 12910 11410 12970
rect 11470 12910 11480 12970
rect 11400 12900 11480 12910
rect 11640 13130 11720 13140
rect 11640 13070 11650 13130
rect 11710 13070 11720 13130
rect 11640 13050 11720 13070
rect 11640 12990 11650 13050
rect 11710 12990 11720 13050
rect 11640 12970 11720 12990
rect 11640 12910 11650 12970
rect 11710 12910 11720 12970
rect 11640 12900 11720 12910
rect 12280 13130 12360 13140
rect 12280 13070 12290 13130
rect 12350 13070 12360 13130
rect 12280 13050 12360 13070
rect 12280 12990 12290 13050
rect 12350 12990 12360 13050
rect 12280 12970 12360 12990
rect 12280 12910 12290 12970
rect 12350 12910 12360 12970
rect 12280 12900 12360 12910
rect 12520 13130 12600 13140
rect 12520 13070 12530 13130
rect 12590 13070 12600 13130
rect 12520 13050 12600 13070
rect 12520 12990 12530 13050
rect 12590 12990 12600 13050
rect 12520 12970 12600 12990
rect 12520 12910 12530 12970
rect 12590 12910 12600 12970
rect 12520 12900 12600 12910
rect 12760 13130 12840 13140
rect 12760 13070 12770 13130
rect 12830 13070 12840 13130
rect 12760 13050 12840 13070
rect 12760 12990 12770 13050
rect 12830 12990 12840 13050
rect 12760 12970 12840 12990
rect 12760 12910 12770 12970
rect 12830 12910 12840 12970
rect 12760 12900 12840 12910
rect 13070 13110 13080 13150
rect 13120 13110 13130 13150
rect 10740 12800 10750 12860
rect 10810 12800 10820 12860
rect 10740 12790 10820 12800
rect 11490 12860 11570 12870
rect 11490 12800 11500 12860
rect 11560 12800 11570 12860
rect 11490 12790 11570 12800
rect 11710 12860 11790 12870
rect 11710 12800 11720 12860
rect 11780 12800 11790 12860
rect 11710 12790 11790 12800
rect 11970 12860 12050 12870
rect 11970 12800 11980 12860
rect 12040 12800 12050 12860
rect 11970 12790 12050 12800
rect 12190 12860 12270 12870
rect 12190 12800 12200 12860
rect 12260 12800 12270 12860
rect 12190 12790 12270 12800
rect 12450 12860 12530 12870
rect 12450 12800 12460 12860
rect 12520 12800 12530 12860
rect 12450 12790 12530 12800
rect 11431 12750 11489 12760
rect 11431 12698 11433 12750
rect 11485 12698 11489 12750
rect 11431 12690 11489 12698
rect 11520 12650 11550 12790
rect 11730 12650 11760 12790
rect 11791 12750 11849 12760
rect 11791 12698 11793 12750
rect 11845 12698 11849 12750
rect 11791 12690 11849 12698
rect 11911 12750 11969 12760
rect 11911 12698 11913 12750
rect 11965 12698 11969 12750
rect 11911 12690 11969 12698
rect 12000 12650 12030 12790
rect 12210 12650 12240 12790
rect 12271 12750 12329 12760
rect 12271 12698 12273 12750
rect 12325 12698 12329 12750
rect 12271 12690 12329 12698
rect 12391 12750 12449 12760
rect 12391 12698 12393 12750
rect 12445 12698 12449 12750
rect 12391 12690 12449 12698
rect 12480 12650 12510 12790
rect 12800 12730 12880 12740
rect 12800 12670 12810 12730
rect 12870 12670 12880 12730
rect 12800 12650 12880 12670
rect 11370 12630 11430 12650
rect 11370 12590 11380 12630
rect 11420 12590 11430 12630
rect 11370 12320 11430 12590
rect 11490 12630 11550 12650
rect 11490 12590 11500 12630
rect 11540 12590 11550 12630
rect 11490 12570 11550 12590
rect 11610 12630 11670 12650
rect 11610 12590 11620 12630
rect 11660 12590 11670 12630
rect 11610 12570 11670 12590
rect 11730 12630 11790 12650
rect 11730 12590 11740 12630
rect 11780 12590 11790 12630
rect 11730 12570 11790 12590
rect 11850 12630 11910 12650
rect 11850 12590 11860 12630
rect 11900 12590 11910 12630
rect 11850 12570 11910 12590
rect 11970 12630 12030 12650
rect 11970 12590 11980 12630
rect 12020 12590 12030 12630
rect 11970 12570 12030 12590
rect 12090 12630 12150 12650
rect 12090 12590 12100 12630
rect 12140 12590 12150 12630
rect 12090 12570 12150 12590
rect 12210 12630 12270 12650
rect 12210 12590 12220 12630
rect 12260 12590 12270 12630
rect 12210 12570 12270 12590
rect 12330 12630 12390 12650
rect 12330 12590 12340 12630
rect 12380 12590 12390 12630
rect 12330 12570 12390 12590
rect 12450 12630 12510 12650
rect 12450 12590 12460 12630
rect 12500 12590 12510 12630
rect 12450 12570 12510 12590
rect 12570 12630 12630 12650
rect 12570 12590 12580 12630
rect 12620 12590 12630 12630
rect 12570 12570 12630 12590
rect 12800 12590 12810 12650
rect 12870 12590 12880 12650
rect 12800 12570 12880 12590
rect 11532 12522 11590 12530
rect 11532 12470 11536 12522
rect 11588 12470 11590 12522
rect 11532 12460 11590 12470
rect 11620 12430 11660 12570
rect 11690 12522 11748 12530
rect 11690 12470 11694 12522
rect 11746 12470 11748 12522
rect 11690 12460 11748 12470
rect 11600 12420 11680 12430
rect 11600 12360 11610 12420
rect 11670 12360 11680 12420
rect 11360 12310 11440 12320
rect 11360 12250 11370 12310
rect 11430 12250 11440 12310
rect 10620 12040 10780 12050
rect 10620 11980 10630 12040
rect 10690 11980 10710 12040
rect 10770 11980 10780 12040
rect 10620 11970 10780 11980
rect 11120 12040 11200 12050
rect 11120 11980 11130 12040
rect 11190 11980 11200 12040
rect 11120 11970 11200 11980
rect 11360 12040 11440 12250
rect 11360 11980 11370 12040
rect 11430 11980 11440 12040
rect 11360 11970 11440 11980
rect 10710 11920 10770 11970
rect 10710 11880 10720 11920
rect 10760 11880 10770 11920
rect 10710 11860 10770 11880
rect 10880 11920 10960 11930
rect 10880 11860 10890 11920
rect 10950 11860 10960 11920
rect 10880 11850 10960 11860
rect 10530 11790 10590 11810
rect 10530 11750 10540 11790
rect 10580 11750 10590 11790
rect 10530 11690 10590 11750
rect 10530 11650 10540 11690
rect 10580 11650 10590 11690
rect 10530 11570 10590 11650
rect 10650 11790 10710 11810
rect 10650 11750 10660 11790
rect 10700 11750 10710 11790
rect 10650 11690 10710 11750
rect 10650 11650 10660 11690
rect 10700 11650 10710 11690
rect 10650 11590 10710 11650
rect 10770 11790 10830 11810
rect 10770 11750 10780 11790
rect 10820 11750 10830 11790
rect 10770 11690 10830 11750
rect 10770 11650 10780 11690
rect 10820 11650 10830 11690
rect 10530 11530 10540 11570
rect 10580 11530 10590 11570
rect 10530 11480 10590 11530
rect 10640 11580 10720 11590
rect 10640 11520 10650 11580
rect 10710 11520 10720 11580
rect 10640 11510 10720 11520
rect 10770 11480 10830 11650
rect 10890 11790 10950 11850
rect 10890 11750 10900 11790
rect 10940 11750 10950 11790
rect 10890 11690 10950 11750
rect 10890 11650 10900 11690
rect 10940 11650 10950 11690
rect 10890 11630 10950 11650
rect 11010 11790 11070 11810
rect 11010 11750 11020 11790
rect 11060 11750 11070 11790
rect 11010 11690 11070 11750
rect 11010 11650 11020 11690
rect 11060 11650 11070 11690
rect 11010 11480 11070 11650
rect 11130 11790 11190 11970
rect 11370 11910 11430 11970
rect 11370 11870 11380 11910
rect 11420 11870 11430 11910
rect 11370 11850 11430 11870
rect 11600 11920 11680 12360
rect 11860 12320 11900 12570
rect 12014 12522 12072 12530
rect 12014 12470 12018 12522
rect 12070 12470 12072 12522
rect 12014 12460 12072 12470
rect 12100 12430 12140 12570
rect 12168 12522 12226 12530
rect 12168 12470 12172 12522
rect 12224 12470 12226 12522
rect 12168 12460 12226 12470
rect 12080 12420 12160 12430
rect 12080 12360 12090 12420
rect 12150 12360 12160 12420
rect 12080 12350 12160 12360
rect 12340 12320 12380 12570
rect 12492 12522 12550 12530
rect 12492 12470 12496 12522
rect 12548 12470 12550 12522
rect 12492 12460 12550 12470
rect 12580 12430 12620 12570
rect 12800 12510 12810 12570
rect 12870 12510 12880 12570
rect 12800 12500 12880 12510
rect 12560 12420 12640 12430
rect 12560 12360 12570 12420
rect 12630 12360 12640 12420
rect 12560 12350 12640 12360
rect 11840 12310 11920 12320
rect 11840 12250 11850 12310
rect 11910 12250 11920 12310
rect 11840 12240 11920 12250
rect 12320 12310 12400 12320
rect 12320 12250 12330 12310
rect 12390 12250 12400 12310
rect 12320 12240 12400 12250
rect 11840 12040 11920 12050
rect 11840 11980 11850 12040
rect 11910 11980 11920 12040
rect 11840 11970 11920 11980
rect 12080 12040 12160 12050
rect 12080 11980 12090 12040
rect 12150 11980 12160 12040
rect 12080 11970 12160 11980
rect 12560 12040 12640 12050
rect 12560 11980 12570 12040
rect 12630 11980 12640 12040
rect 12560 11970 12640 11980
rect 12740 12040 12820 12050
rect 12740 11980 12750 12040
rect 12810 11980 12820 12040
rect 12740 11970 12820 11980
rect 11600 11860 11610 11920
rect 11670 11860 11680 11920
rect 11600 11850 11680 11860
rect 11130 11750 11140 11790
rect 11180 11750 11190 11790
rect 11130 11690 11190 11750
rect 11130 11650 11140 11690
rect 11180 11650 11190 11690
rect 11130 11630 11190 11650
rect 11250 11790 11310 11810
rect 11250 11750 11260 11790
rect 11300 11750 11310 11790
rect 11250 11690 11310 11750
rect 11250 11650 11260 11690
rect 11300 11650 11310 11690
rect 11250 11480 11310 11650
rect 11370 11790 11430 11810
rect 11370 11750 11380 11790
rect 11420 11750 11430 11790
rect 11370 11690 11430 11750
rect 11370 11650 11380 11690
rect 11420 11650 11430 11690
rect 11370 11590 11430 11650
rect 11490 11790 11550 11810
rect 11490 11750 11500 11790
rect 11540 11750 11550 11790
rect 11490 11690 11550 11750
rect 11490 11650 11500 11690
rect 11540 11650 11550 11690
rect 11360 11580 11440 11590
rect 11360 11520 11370 11580
rect 11430 11520 11440 11580
rect 11360 11510 11440 11520
rect 11490 11480 11550 11650
rect 11610 11790 11670 11850
rect 11610 11750 11620 11790
rect 11660 11750 11670 11790
rect 11610 11690 11670 11750
rect 11610 11650 11620 11690
rect 11660 11650 11670 11690
rect 11610 11630 11670 11650
rect 11730 11790 11790 11810
rect 11730 11750 11740 11790
rect 11780 11750 11790 11790
rect 11730 11690 11790 11750
rect 11730 11650 11740 11690
rect 11780 11650 11790 11690
rect 11730 11480 11790 11650
rect 11850 11790 11910 11970
rect 12090 11910 12150 11970
rect 12090 11870 12100 11910
rect 12140 11870 12150 11910
rect 12090 11850 12150 11870
rect 12320 11920 12400 11930
rect 12320 11860 12330 11920
rect 12390 11860 12400 11920
rect 12320 11850 12400 11860
rect 11850 11750 11860 11790
rect 11900 11750 11910 11790
rect 11850 11690 11910 11750
rect 11850 11650 11860 11690
rect 11900 11650 11910 11690
rect 11850 11630 11910 11650
rect 11970 11790 12030 11810
rect 11970 11750 11980 11790
rect 12020 11750 12030 11790
rect 11970 11690 12030 11750
rect 11970 11650 11980 11690
rect 12020 11650 12030 11690
rect 11970 11480 12030 11650
rect 12090 11790 12150 11810
rect 12090 11750 12100 11790
rect 12140 11750 12150 11790
rect 12090 11690 12150 11750
rect 12090 11650 12100 11690
rect 12140 11650 12150 11690
rect 12090 11590 12150 11650
rect 12210 11790 12270 11810
rect 12210 11750 12220 11790
rect 12260 11750 12270 11790
rect 12210 11690 12270 11750
rect 12210 11650 12220 11690
rect 12260 11650 12270 11690
rect 12080 11580 12160 11590
rect 12080 11520 12090 11580
rect 12150 11520 12160 11580
rect 12080 11510 12160 11520
rect 12210 11480 12270 11650
rect 12330 11790 12390 11850
rect 12330 11750 12340 11790
rect 12380 11750 12390 11790
rect 12330 11690 12390 11750
rect 12330 11650 12340 11690
rect 12380 11650 12390 11690
rect 12330 11630 12390 11650
rect 12450 11790 12510 11810
rect 12450 11750 12460 11790
rect 12500 11750 12510 11790
rect 12450 11690 12510 11750
rect 12450 11650 12460 11690
rect 12500 11650 12510 11690
rect 12450 11480 12510 11650
rect 12570 11790 12630 11970
rect 12750 11910 12810 11970
rect 12750 11870 12760 11910
rect 12800 11870 12810 11910
rect 12750 11850 12810 11870
rect 12570 11750 12580 11790
rect 12620 11750 12630 11790
rect 12570 11690 12630 11750
rect 12570 11650 12580 11690
rect 12620 11650 12630 11690
rect 12570 11630 12630 11650
rect 12690 11790 12750 11810
rect 12690 11750 12700 11790
rect 12740 11750 12750 11790
rect 12690 11690 12750 11750
rect 12690 11650 12700 11690
rect 12740 11650 12750 11690
rect 12690 11480 12750 11650
rect 12810 11790 12870 11810
rect 12810 11750 12820 11790
rect 12860 11750 12870 11790
rect 12810 11690 12870 11750
rect 12810 11650 12820 11690
rect 12860 11650 12870 11690
rect 12810 11590 12870 11650
rect 12930 11790 12990 11810
rect 12930 11750 12940 11790
rect 12980 11750 12990 11790
rect 12930 11690 12990 11750
rect 12930 11650 12940 11690
rect 12980 11650 12990 11690
rect 12800 11580 12880 11590
rect 12800 11520 12810 11580
rect 12870 11520 12880 11580
rect 12800 11510 12880 11520
rect 12930 11570 12990 11650
rect 13070 11590 13130 13110
rect 13160 12730 13400 13710
rect 14580 13930 14660 13940
rect 14580 13870 14590 13930
rect 14650 13870 14660 13930
rect 14580 13850 14660 13870
rect 14580 13790 14590 13850
rect 14650 13790 14660 13850
rect 14580 13770 14660 13790
rect 14580 13710 14590 13770
rect 14650 13710 14660 13770
rect 14580 13700 14660 13710
rect 15750 13640 15810 13660
rect 15750 13600 15760 13640
rect 15800 13600 15810 13640
rect 15750 13540 15810 13600
rect 15750 13500 15760 13540
rect 15800 13500 15810 13540
rect 15750 13440 15810 13500
rect 15750 13400 15760 13440
rect 15800 13400 15810 13440
rect 15750 13340 15810 13400
rect 15750 13300 15760 13340
rect 15800 13300 15810 13340
rect 15750 13240 15810 13300
rect 15750 13200 15760 13240
rect 15800 13200 15810 13240
rect 13160 12670 13170 12730
rect 13230 12670 13250 12730
rect 13310 12670 13330 12730
rect 13390 12670 13400 12730
rect 13160 12650 13400 12670
rect 13160 12590 13170 12650
rect 13230 12590 13250 12650
rect 13310 12590 13330 12650
rect 13390 12590 13400 12650
rect 13160 12570 13400 12590
rect 13160 12510 13170 12570
rect 13230 12510 13250 12570
rect 13310 12510 13330 12570
rect 13390 12510 13400 12570
rect 13160 12500 13400 12510
rect 13430 13150 13490 13170
rect 13430 13110 13440 13150
rect 13480 13110 13490 13150
rect 13430 11590 13490 13110
rect 13720 13130 13800 13140
rect 13720 13070 13730 13130
rect 13790 13070 13800 13130
rect 13720 13050 13800 13070
rect 13720 12990 13730 13050
rect 13790 12990 13800 13050
rect 13720 12970 13800 12990
rect 13720 12910 13730 12970
rect 13790 12910 13800 12970
rect 13720 12900 13800 12910
rect 13960 13130 14040 13140
rect 13960 13070 13970 13130
rect 14030 13070 14040 13130
rect 13960 13050 14040 13070
rect 13960 12990 13970 13050
rect 14030 12990 14040 13050
rect 13960 12970 14040 12990
rect 13960 12910 13970 12970
rect 14030 12910 14040 12970
rect 13960 12900 14040 12910
rect 14200 13130 14280 13140
rect 14200 13070 14210 13130
rect 14270 13070 14280 13130
rect 14200 13050 14280 13070
rect 14200 12990 14210 13050
rect 14270 12990 14280 13050
rect 14200 12970 14280 12990
rect 14200 12910 14210 12970
rect 14270 12910 14280 12970
rect 14200 12900 14280 12910
rect 14840 13130 14920 13140
rect 14840 13070 14850 13130
rect 14910 13070 14920 13130
rect 14840 13050 14920 13070
rect 14840 12990 14850 13050
rect 14910 12990 14920 13050
rect 14840 12970 14920 12990
rect 14840 12910 14850 12970
rect 14910 12910 14920 12970
rect 14840 12900 14920 12910
rect 15080 13130 15160 13140
rect 15080 13070 15090 13130
rect 15150 13070 15160 13130
rect 15080 13050 15160 13070
rect 15080 12990 15090 13050
rect 15150 12990 15160 13050
rect 15080 12970 15160 12990
rect 15080 12910 15090 12970
rect 15150 12910 15160 12970
rect 15080 12900 15160 12910
rect 15320 13130 15400 13140
rect 15320 13070 15330 13130
rect 15390 13070 15400 13130
rect 15320 13050 15400 13070
rect 15320 12990 15330 13050
rect 15390 12990 15400 13050
rect 15320 12970 15400 12990
rect 15320 12910 15330 12970
rect 15390 12910 15400 12970
rect 15320 12900 15400 12910
rect 15560 13130 15640 13140
rect 15560 13070 15570 13130
rect 15630 13070 15640 13130
rect 15560 13050 15640 13070
rect 15560 12990 15570 13050
rect 15630 12990 15640 13050
rect 15560 12970 15640 12990
rect 15560 12910 15570 12970
rect 15630 12910 15640 12970
rect 15560 12900 15640 12910
rect 15750 12870 15810 13200
rect 14030 12860 14110 12870
rect 14030 12800 14040 12860
rect 14100 12800 14110 12860
rect 14030 12790 14110 12800
rect 14290 12860 14370 12870
rect 14290 12800 14300 12860
rect 14360 12800 14370 12860
rect 14290 12790 14370 12800
rect 14510 12860 14590 12870
rect 14510 12800 14520 12860
rect 14580 12800 14590 12860
rect 14510 12790 14590 12800
rect 14770 12860 14850 12870
rect 14770 12800 14780 12860
rect 14840 12800 14850 12860
rect 14770 12790 14850 12800
rect 14990 12860 15070 12870
rect 14990 12800 15000 12860
rect 15060 12800 15070 12860
rect 14990 12790 15070 12800
rect 15740 12860 15820 12870
rect 15740 12800 15750 12860
rect 15810 12800 15820 12860
rect 15740 12790 15820 12800
rect 13680 12730 13760 12740
rect 13680 12670 13690 12730
rect 13750 12670 13760 12730
rect 13680 12650 13760 12670
rect 14050 12650 14080 12790
rect 14111 12750 14169 12760
rect 14111 12698 14115 12750
rect 14167 12698 14169 12750
rect 14111 12690 14169 12698
rect 14231 12750 14289 12760
rect 14231 12698 14235 12750
rect 14287 12698 14289 12750
rect 14231 12690 14289 12698
rect 14320 12650 14350 12790
rect 14530 12650 14560 12790
rect 14591 12750 14649 12760
rect 14591 12698 14595 12750
rect 14647 12698 14649 12750
rect 14591 12690 14649 12698
rect 14711 12750 14769 12760
rect 14711 12698 14715 12750
rect 14767 12698 14769 12750
rect 14711 12690 14769 12698
rect 14800 12650 14830 12790
rect 15010 12650 15040 12790
rect 16170 12760 16210 14530
rect 15071 12750 15129 12760
rect 15071 12698 15075 12750
rect 15127 12698 15129 12750
rect 15071 12690 15129 12698
rect 16150 12750 16230 12760
rect 16150 12690 16160 12750
rect 16220 12690 16230 12750
rect 16150 12680 16230 12690
rect 13680 12590 13690 12650
rect 13750 12590 13760 12650
rect 13680 12570 13760 12590
rect 13930 12630 13990 12650
rect 13930 12590 13940 12630
rect 13980 12590 13990 12630
rect 13930 12570 13990 12590
rect 14050 12630 14110 12650
rect 14050 12590 14060 12630
rect 14100 12590 14110 12630
rect 14050 12570 14110 12590
rect 14170 12630 14230 12650
rect 14170 12590 14180 12630
rect 14220 12590 14230 12630
rect 14170 12570 14230 12590
rect 14290 12630 14350 12650
rect 14290 12590 14300 12630
rect 14340 12590 14350 12630
rect 14290 12570 14350 12590
rect 14410 12630 14470 12650
rect 14410 12590 14420 12630
rect 14460 12590 14470 12630
rect 14410 12570 14470 12590
rect 14530 12630 14590 12650
rect 14530 12590 14540 12630
rect 14580 12590 14590 12630
rect 14530 12570 14590 12590
rect 14650 12630 14710 12650
rect 14650 12590 14660 12630
rect 14700 12590 14710 12630
rect 14650 12570 14710 12590
rect 14770 12630 14830 12650
rect 14770 12590 14780 12630
rect 14820 12590 14830 12630
rect 14770 12570 14830 12590
rect 14890 12630 14950 12650
rect 14890 12590 14900 12630
rect 14940 12590 14950 12630
rect 14890 12570 14950 12590
rect 15010 12630 15070 12650
rect 15010 12590 15020 12630
rect 15060 12590 15070 12630
rect 15010 12570 15070 12590
rect 15130 12630 15190 12650
rect 15130 12590 15140 12630
rect 15180 12590 15190 12630
rect 13680 12510 13690 12570
rect 13750 12510 13760 12570
rect 13680 12500 13760 12510
rect 13940 12430 13980 12570
rect 14010 12522 14068 12530
rect 14010 12470 14012 12522
rect 14064 12470 14068 12522
rect 14010 12460 14068 12470
rect 13920 12420 14000 12430
rect 13920 12360 13930 12420
rect 13990 12360 14000 12420
rect 13920 12350 14000 12360
rect 14180 12320 14220 12570
rect 14334 12522 14392 12530
rect 14334 12470 14336 12522
rect 14388 12470 14392 12522
rect 14334 12460 14392 12470
rect 14420 12430 14460 12570
rect 14488 12522 14546 12530
rect 14488 12470 14490 12522
rect 14542 12470 14546 12522
rect 14488 12460 14546 12470
rect 14400 12420 14480 12430
rect 14400 12360 14410 12420
rect 14470 12360 14480 12420
rect 14400 12350 14480 12360
rect 14660 12320 14700 12570
rect 14812 12522 14870 12530
rect 14812 12470 14814 12522
rect 14866 12470 14870 12522
rect 14812 12460 14870 12470
rect 14900 12430 14940 12570
rect 14970 12522 15028 12530
rect 14970 12470 14972 12522
rect 15024 12470 15028 12522
rect 14970 12460 15028 12470
rect 14880 12420 14960 12430
rect 14880 12360 14890 12420
rect 14950 12360 14960 12420
rect 14160 12310 14240 12320
rect 14160 12250 14170 12310
rect 14230 12250 14240 12310
rect 14160 12240 14240 12250
rect 14640 12310 14720 12320
rect 14640 12250 14650 12310
rect 14710 12250 14720 12310
rect 14640 12240 14720 12250
rect 13740 12200 13820 12210
rect 13740 12140 13750 12200
rect 13810 12140 13820 12200
rect 13740 12120 13820 12140
rect 13740 12060 13750 12120
rect 13810 12060 13820 12120
rect 13740 12040 13820 12060
rect 13740 11980 13750 12040
rect 13810 11980 13820 12040
rect 13740 11970 13820 11980
rect 13920 12200 14000 12210
rect 13920 12140 13930 12200
rect 13990 12140 14000 12200
rect 13920 12120 14000 12140
rect 13920 12060 13930 12120
rect 13990 12060 14000 12120
rect 13920 12040 14000 12060
rect 13920 11980 13930 12040
rect 13990 11980 14000 12040
rect 13920 11970 14000 11980
rect 14160 12200 14240 12210
rect 14160 12140 14170 12200
rect 14230 12140 14240 12200
rect 14160 12120 14240 12140
rect 14160 12060 14170 12120
rect 14230 12060 14240 12120
rect 14160 12040 14240 12060
rect 14160 11980 14170 12040
rect 14230 11980 14240 12040
rect 14160 11970 14240 11980
rect 14400 12200 14480 12210
rect 14400 12140 14410 12200
rect 14470 12140 14480 12200
rect 14400 12120 14480 12140
rect 14400 12060 14410 12120
rect 14470 12060 14480 12120
rect 14400 12040 14480 12060
rect 14400 11980 14410 12040
rect 14470 11980 14480 12040
rect 14400 11970 14480 11980
rect 14640 12200 14720 12210
rect 14640 12140 14650 12200
rect 14710 12140 14720 12200
rect 14640 12120 14720 12140
rect 14640 12060 14650 12120
rect 14710 12060 14720 12120
rect 14640 12040 14720 12060
rect 14640 11980 14650 12040
rect 14710 11980 14720 12040
rect 14640 11970 14720 11980
rect 13750 11910 13810 11970
rect 13750 11870 13760 11910
rect 13800 11870 13810 11910
rect 13750 11850 13810 11870
rect 13570 11790 13630 11810
rect 13570 11750 13580 11790
rect 13620 11750 13630 11790
rect 13570 11690 13630 11750
rect 13570 11650 13580 11690
rect 13620 11650 13630 11690
rect 12930 11530 12940 11570
rect 12980 11530 12990 11570
rect 12930 11480 12990 11530
rect 13060 11580 13140 11590
rect 13060 11520 13070 11580
rect 13130 11520 13140 11580
rect 13060 11510 13140 11520
rect 13420 11580 13500 11590
rect 13420 11520 13430 11580
rect 13490 11520 13500 11580
rect 10520 11470 10600 11480
rect 10520 11410 10530 11470
rect 10590 11410 10600 11470
rect 10520 11390 10600 11410
rect 10520 11330 10530 11390
rect 10590 11330 10600 11390
rect 10520 11310 10600 11330
rect 10520 11250 10530 11310
rect 10590 11250 10600 11310
rect 10520 11240 10600 11250
rect 10760 11470 10840 11480
rect 10760 11410 10770 11470
rect 10830 11410 10840 11470
rect 10760 11390 10840 11410
rect 10760 11330 10770 11390
rect 10830 11330 10840 11390
rect 10760 11310 10840 11330
rect 10760 11250 10770 11310
rect 10830 11250 10840 11310
rect 10760 11240 10840 11250
rect 11000 11470 11080 11480
rect 11000 11410 11010 11470
rect 11070 11410 11080 11470
rect 11000 11390 11080 11410
rect 11000 11330 11010 11390
rect 11070 11330 11080 11390
rect 11000 11310 11080 11330
rect 11000 11250 11010 11310
rect 11070 11250 11080 11310
rect 11000 11240 11080 11250
rect 11240 11470 11320 11480
rect 11240 11410 11250 11470
rect 11310 11410 11320 11470
rect 11240 11390 11320 11410
rect 11240 11330 11250 11390
rect 11310 11330 11320 11390
rect 11240 11310 11320 11330
rect 11240 11250 11250 11310
rect 11310 11250 11320 11310
rect 11240 11240 11320 11250
rect 11480 11470 11560 11480
rect 11480 11410 11490 11470
rect 11550 11410 11560 11470
rect 11480 11390 11560 11410
rect 11480 11330 11490 11390
rect 11550 11330 11560 11390
rect 11480 11310 11560 11330
rect 11480 11250 11490 11310
rect 11550 11250 11560 11310
rect 11480 11240 11560 11250
rect 11720 11470 11800 11480
rect 11720 11410 11730 11470
rect 11790 11410 11800 11470
rect 11720 11390 11800 11410
rect 11720 11330 11730 11390
rect 11790 11330 11800 11390
rect 11720 11310 11800 11330
rect 11720 11250 11730 11310
rect 11790 11250 11800 11310
rect 11720 11240 11800 11250
rect 11960 11470 12040 11480
rect 11960 11410 11970 11470
rect 12030 11410 12040 11470
rect 11960 11390 12040 11410
rect 11960 11330 11970 11390
rect 12030 11330 12040 11390
rect 11960 11310 12040 11330
rect 11960 11250 11970 11310
rect 12030 11250 12040 11310
rect 11960 11240 12040 11250
rect 12200 11470 12280 11480
rect 12200 11410 12210 11470
rect 12270 11410 12280 11470
rect 12200 11390 12280 11410
rect 12200 11330 12210 11390
rect 12270 11330 12280 11390
rect 12200 11310 12280 11330
rect 12200 11250 12210 11310
rect 12270 11250 12280 11310
rect 12200 11240 12280 11250
rect 12440 11470 12520 11480
rect 12440 11410 12450 11470
rect 12510 11410 12520 11470
rect 12440 11390 12520 11410
rect 12440 11330 12450 11390
rect 12510 11330 12520 11390
rect 12440 11310 12520 11330
rect 12440 11250 12450 11310
rect 12510 11250 12520 11310
rect 12440 11240 12520 11250
rect 12680 11470 12760 11480
rect 12680 11410 12690 11470
rect 12750 11410 12760 11470
rect 12680 11390 12760 11410
rect 12680 11330 12690 11390
rect 12750 11330 12760 11390
rect 12680 11310 12760 11330
rect 12680 11250 12690 11310
rect 12750 11250 12760 11310
rect 12680 11240 12760 11250
rect 12920 11470 13000 11480
rect 12920 11410 12930 11470
rect 12990 11410 13000 11470
rect 12920 11390 13000 11410
rect 12920 11330 12930 11390
rect 12990 11330 13000 11390
rect 12920 11310 13000 11330
rect 12920 11250 12930 11310
rect 12990 11250 13000 11310
rect 12920 11240 13000 11250
rect 11800 11200 11880 11210
rect 11800 11140 11810 11200
rect 11870 11140 11880 11200
rect 11800 11130 11880 11140
rect 13240 11200 13320 11210
rect 13240 11140 13250 11200
rect 13310 11140 13320 11200
rect 13240 11130 13320 11140
rect 11630 10630 11690 10650
rect 11630 10590 11640 10630
rect 11680 10590 11690 10630
rect 11630 10530 11690 10590
rect 11630 10490 11640 10530
rect 11680 10490 11690 10530
rect 11630 10430 11690 10490
rect 11630 10390 11640 10430
rect 11680 10390 11690 10430
rect 11630 10330 11690 10390
rect 11630 10290 11640 10330
rect 11680 10290 11690 10330
rect 11630 10230 11690 10290
rect 11630 10190 11640 10230
rect 11680 10190 11690 10230
rect 11630 10130 11690 10190
rect 11630 10090 11640 10130
rect 11680 10090 11690 10130
rect 11630 10070 11690 10090
rect 11810 10630 11870 11130
rect 12160 11090 12240 11100
rect 12160 11030 12170 11090
rect 12230 11030 12240 11090
rect 12160 11020 12240 11030
rect 11900 10760 11970 10770
rect 11960 10700 11970 10760
rect 11900 10690 11970 10700
rect 12070 10760 12150 10770
rect 12070 10700 12080 10760
rect 12140 10700 12150 10760
rect 12070 10690 12150 10700
rect 12180 10650 12220 11020
rect 12520 10980 12600 10990
rect 12520 10920 12530 10980
rect 12590 10920 12600 10980
rect 12520 10910 12600 10920
rect 12250 10760 12330 10770
rect 12250 10700 12260 10760
rect 12320 10700 12330 10760
rect 12250 10690 12330 10700
rect 12430 10760 12510 10770
rect 12430 10700 12440 10760
rect 12500 10700 12510 10760
rect 12430 10690 12510 10700
rect 12540 10650 12580 10910
rect 12880 10870 12960 10880
rect 12880 10810 12890 10870
rect 12950 10810 12960 10870
rect 12880 10800 12960 10810
rect 12610 10760 12690 10770
rect 12610 10700 12620 10760
rect 12680 10700 12690 10760
rect 12610 10690 12690 10700
rect 12790 10760 12870 10770
rect 12790 10700 12800 10760
rect 12860 10700 12870 10760
rect 12790 10690 12870 10700
rect 12900 10650 12940 10800
rect 12970 10760 13050 10770
rect 12970 10700 12980 10760
rect 13040 10700 13050 10760
rect 12970 10690 13050 10700
rect 13150 10760 13220 10770
rect 13150 10700 13160 10760
rect 13150 10690 13220 10700
rect 11810 10590 11820 10630
rect 11860 10590 11870 10630
rect 11810 10530 11870 10590
rect 11810 10490 11820 10530
rect 11860 10490 11870 10530
rect 11810 10430 11870 10490
rect 11810 10390 11820 10430
rect 11860 10390 11870 10430
rect 11810 10330 11870 10390
rect 11810 10290 11820 10330
rect 11860 10290 11870 10330
rect 11810 10230 11870 10290
rect 11810 10190 11820 10230
rect 11860 10190 11870 10230
rect 11810 10130 11870 10190
rect 11810 10090 11820 10130
rect 11860 10090 11870 10130
rect 11810 10070 11870 10090
rect 11990 10630 12050 10650
rect 11990 10590 12000 10630
rect 12040 10590 12050 10630
rect 11990 10530 12050 10590
rect 11990 10490 12000 10530
rect 12040 10490 12050 10530
rect 11990 10430 12050 10490
rect 11990 10390 12000 10430
rect 12040 10390 12050 10430
rect 11990 10330 12050 10390
rect 11990 10290 12000 10330
rect 12040 10290 12050 10330
rect 11990 10230 12050 10290
rect 11990 10190 12000 10230
rect 12040 10190 12050 10230
rect 11990 10130 12050 10190
rect 11990 10090 12000 10130
rect 12040 10090 12050 10130
rect 11990 10070 12050 10090
rect 12170 10630 12230 10650
rect 12170 10590 12180 10630
rect 12220 10590 12230 10630
rect 12170 10530 12230 10590
rect 12170 10490 12180 10530
rect 12220 10490 12230 10530
rect 12170 10430 12230 10490
rect 12170 10390 12180 10430
rect 12220 10390 12230 10430
rect 12170 10330 12230 10390
rect 12170 10290 12180 10330
rect 12220 10290 12230 10330
rect 12170 10230 12230 10290
rect 12170 10190 12180 10230
rect 12220 10190 12230 10230
rect 12170 10130 12230 10190
rect 12170 10090 12180 10130
rect 12220 10090 12230 10130
rect 12170 10070 12230 10090
rect 12350 10630 12410 10650
rect 12350 10590 12360 10630
rect 12400 10590 12410 10630
rect 12350 10530 12410 10590
rect 12350 10490 12360 10530
rect 12400 10490 12410 10530
rect 12350 10430 12410 10490
rect 12350 10390 12360 10430
rect 12400 10390 12410 10430
rect 12350 10330 12410 10390
rect 12350 10290 12360 10330
rect 12400 10290 12410 10330
rect 12350 10230 12410 10290
rect 12350 10190 12360 10230
rect 12400 10190 12410 10230
rect 12350 10130 12410 10190
rect 12350 10090 12360 10130
rect 12400 10090 12410 10130
rect 12350 10070 12410 10090
rect 12530 10630 12590 10650
rect 12530 10590 12540 10630
rect 12580 10590 12590 10630
rect 12530 10530 12590 10590
rect 12530 10490 12540 10530
rect 12580 10490 12590 10530
rect 12530 10430 12590 10490
rect 12530 10390 12540 10430
rect 12580 10390 12590 10430
rect 12530 10330 12590 10390
rect 12530 10290 12540 10330
rect 12580 10290 12590 10330
rect 12530 10230 12590 10290
rect 12530 10190 12540 10230
rect 12580 10190 12590 10230
rect 12530 10130 12590 10190
rect 12530 10090 12540 10130
rect 12580 10090 12590 10130
rect 12530 10070 12590 10090
rect 12710 10630 12770 10650
rect 12710 10590 12720 10630
rect 12760 10590 12770 10630
rect 12710 10530 12770 10590
rect 12710 10490 12720 10530
rect 12760 10490 12770 10530
rect 12710 10430 12770 10490
rect 12710 10390 12720 10430
rect 12760 10390 12770 10430
rect 12710 10330 12770 10390
rect 12710 10290 12720 10330
rect 12760 10290 12770 10330
rect 12710 10230 12770 10290
rect 12710 10190 12720 10230
rect 12760 10190 12770 10230
rect 12710 10130 12770 10190
rect 12710 10090 12720 10130
rect 12760 10090 12770 10130
rect 12710 10070 12770 10090
rect 12890 10630 12950 10650
rect 12890 10590 12900 10630
rect 12940 10590 12950 10630
rect 12890 10530 12950 10590
rect 12890 10490 12900 10530
rect 12940 10490 12950 10530
rect 12890 10430 12950 10490
rect 12890 10390 12900 10430
rect 12940 10390 12950 10430
rect 12890 10330 12950 10390
rect 12890 10290 12900 10330
rect 12940 10290 12950 10330
rect 12890 10230 12950 10290
rect 12890 10190 12900 10230
rect 12940 10190 12950 10230
rect 12890 10130 12950 10190
rect 12890 10090 12900 10130
rect 12940 10090 12950 10130
rect 12890 10070 12950 10090
rect 13070 10630 13130 10650
rect 13070 10590 13080 10630
rect 13120 10590 13130 10630
rect 13070 10530 13130 10590
rect 13070 10490 13080 10530
rect 13120 10490 13130 10530
rect 13070 10430 13130 10490
rect 13070 10390 13080 10430
rect 13120 10390 13130 10430
rect 13070 10330 13130 10390
rect 13070 10290 13080 10330
rect 13120 10290 13130 10330
rect 13070 10230 13130 10290
rect 13070 10190 13080 10230
rect 13120 10190 13130 10230
rect 13070 10130 13130 10190
rect 13070 10090 13080 10130
rect 13120 10090 13130 10130
rect 13070 10070 13130 10090
rect 13250 10630 13310 11130
rect 13420 10770 13500 11520
rect 13570 11570 13630 11650
rect 13690 11790 13750 11810
rect 13690 11750 13700 11790
rect 13740 11750 13750 11790
rect 13690 11690 13750 11750
rect 13690 11650 13700 11690
rect 13740 11650 13750 11690
rect 13690 11590 13750 11650
rect 13810 11790 13870 11810
rect 13810 11750 13820 11790
rect 13860 11750 13870 11790
rect 13810 11690 13870 11750
rect 13810 11650 13820 11690
rect 13860 11650 13870 11690
rect 13570 11530 13580 11570
rect 13620 11530 13630 11570
rect 13570 11480 13630 11530
rect 13680 11580 13760 11590
rect 13680 11520 13690 11580
rect 13750 11520 13760 11580
rect 13680 11510 13760 11520
rect 13810 11480 13870 11650
rect 13930 11790 13990 11970
rect 14160 11920 14240 11930
rect 14160 11860 14170 11920
rect 14230 11860 14240 11920
rect 14160 11850 14240 11860
rect 14410 11910 14470 11970
rect 14410 11870 14420 11910
rect 14460 11870 14470 11910
rect 14410 11850 14470 11870
rect 13930 11750 13940 11790
rect 13980 11750 13990 11790
rect 13930 11690 13990 11750
rect 13930 11650 13940 11690
rect 13980 11650 13990 11690
rect 13930 11630 13990 11650
rect 14050 11790 14110 11810
rect 14050 11750 14060 11790
rect 14100 11750 14110 11790
rect 14050 11690 14110 11750
rect 14050 11650 14060 11690
rect 14100 11650 14110 11690
rect 14050 11480 14110 11650
rect 14170 11790 14230 11850
rect 14170 11750 14180 11790
rect 14220 11750 14230 11790
rect 14170 11690 14230 11750
rect 14170 11650 14180 11690
rect 14220 11650 14230 11690
rect 14170 11630 14230 11650
rect 14290 11790 14350 11810
rect 14290 11750 14300 11790
rect 14340 11750 14350 11790
rect 14290 11690 14350 11750
rect 14290 11650 14300 11690
rect 14340 11650 14350 11690
rect 14290 11480 14350 11650
rect 14410 11790 14470 11810
rect 14410 11750 14420 11790
rect 14460 11750 14470 11790
rect 14410 11690 14470 11750
rect 14410 11650 14420 11690
rect 14460 11650 14470 11690
rect 14410 11590 14470 11650
rect 14530 11790 14590 11810
rect 14530 11750 14540 11790
rect 14580 11750 14590 11790
rect 14530 11690 14590 11750
rect 14530 11650 14540 11690
rect 14580 11650 14590 11690
rect 14400 11580 14480 11590
rect 14400 11520 14410 11580
rect 14470 11520 14480 11580
rect 14400 11510 14480 11520
rect 14530 11480 14590 11650
rect 14650 11790 14710 11970
rect 14880 11920 14960 12360
rect 15130 12320 15190 12590
rect 15120 12310 15200 12320
rect 15120 12250 15130 12310
rect 15190 12250 15200 12310
rect 15120 12200 15200 12250
rect 15120 12140 15130 12200
rect 15190 12140 15200 12200
rect 15120 12120 15200 12140
rect 15120 12060 15130 12120
rect 15190 12060 15200 12120
rect 15120 12040 15200 12060
rect 15120 11980 15130 12040
rect 15190 11980 15200 12040
rect 15120 11970 15200 11980
rect 15360 12200 15440 12210
rect 15360 12140 15370 12200
rect 15430 12140 15440 12200
rect 15360 12120 15440 12140
rect 15360 12060 15370 12120
rect 15430 12060 15440 12120
rect 15360 12040 15440 12060
rect 15360 11980 15370 12040
rect 15430 11980 15440 12040
rect 15360 11970 15440 11980
rect 15780 12200 15860 12210
rect 15780 12140 15790 12200
rect 15850 12140 15860 12200
rect 15780 12120 15860 12140
rect 15780 12060 15790 12120
rect 15850 12060 15860 12120
rect 15780 12040 15860 12060
rect 15780 11980 15790 12040
rect 15850 11980 15860 12040
rect 15780 11970 15860 11980
rect 14880 11860 14890 11920
rect 14950 11860 14960 11920
rect 14880 11850 14960 11860
rect 15130 11910 15190 11970
rect 15130 11870 15140 11910
rect 15180 11870 15190 11910
rect 15130 11850 15190 11870
rect 14650 11750 14660 11790
rect 14700 11750 14710 11790
rect 14650 11690 14710 11750
rect 14650 11650 14660 11690
rect 14700 11650 14710 11690
rect 14650 11630 14710 11650
rect 14770 11790 14830 11810
rect 14770 11750 14780 11790
rect 14820 11750 14830 11790
rect 14770 11690 14830 11750
rect 14770 11650 14780 11690
rect 14820 11650 14830 11690
rect 14770 11480 14830 11650
rect 14890 11790 14950 11850
rect 14890 11750 14900 11790
rect 14940 11750 14950 11790
rect 14890 11690 14950 11750
rect 14890 11650 14900 11690
rect 14940 11650 14950 11690
rect 14890 11630 14950 11650
rect 15010 11790 15070 11810
rect 15010 11750 15020 11790
rect 15060 11750 15070 11790
rect 15010 11690 15070 11750
rect 15010 11650 15020 11690
rect 15060 11650 15070 11690
rect 15010 11480 15070 11650
rect 15130 11790 15190 11810
rect 15130 11750 15140 11790
rect 15180 11750 15190 11790
rect 15130 11690 15190 11750
rect 15130 11650 15140 11690
rect 15180 11650 15190 11690
rect 15130 11590 15190 11650
rect 15250 11790 15310 11810
rect 15250 11750 15260 11790
rect 15300 11750 15310 11790
rect 15250 11690 15310 11750
rect 15250 11650 15260 11690
rect 15300 11650 15310 11690
rect 15120 11580 15200 11590
rect 15120 11520 15130 11580
rect 15190 11520 15200 11580
rect 15120 11510 15200 11520
rect 15250 11480 15310 11650
rect 15370 11790 15430 11970
rect 15600 11920 15680 11930
rect 15600 11860 15610 11920
rect 15670 11860 15680 11920
rect 15790 11920 15850 11970
rect 15790 11880 15800 11920
rect 15840 11880 15850 11920
rect 15790 11860 15850 11880
rect 15600 11850 15680 11860
rect 15370 11750 15380 11790
rect 15420 11750 15430 11790
rect 15370 11690 15430 11750
rect 15370 11650 15380 11690
rect 15420 11650 15430 11690
rect 15370 11630 15430 11650
rect 15490 11790 15550 11810
rect 15490 11750 15500 11790
rect 15540 11750 15550 11790
rect 15490 11690 15550 11750
rect 15490 11650 15500 11690
rect 15540 11650 15550 11690
rect 15490 11480 15550 11650
rect 15610 11790 15670 11850
rect 15610 11750 15620 11790
rect 15660 11750 15670 11790
rect 15610 11690 15670 11750
rect 15610 11650 15620 11690
rect 15660 11650 15670 11690
rect 15610 11630 15670 11650
rect 15730 11790 15790 11810
rect 15730 11750 15740 11790
rect 15780 11750 15790 11790
rect 15730 11690 15790 11750
rect 15730 11650 15740 11690
rect 15780 11650 15790 11690
rect 15730 11480 15790 11650
rect 15850 11790 15910 11810
rect 15850 11750 15860 11790
rect 15900 11750 15910 11790
rect 15850 11690 15910 11750
rect 15850 11650 15860 11690
rect 15900 11650 15910 11690
rect 15850 11590 15910 11650
rect 15970 11790 16030 11810
rect 15970 11750 15980 11790
rect 16020 11750 16030 11790
rect 15970 11690 16030 11750
rect 15970 11650 15980 11690
rect 16020 11650 16030 11690
rect 15840 11580 15920 11590
rect 15840 11520 15850 11580
rect 15910 11520 15920 11580
rect 13560 11470 13640 11480
rect 13560 11410 13570 11470
rect 13630 11410 13640 11470
rect 13560 11390 13640 11410
rect 13560 11330 13570 11390
rect 13630 11330 13640 11390
rect 13560 11310 13640 11330
rect 13560 11250 13570 11310
rect 13630 11250 13640 11310
rect 13560 11240 13640 11250
rect 13800 11470 13880 11480
rect 13800 11410 13810 11470
rect 13870 11410 13880 11470
rect 13800 11390 13880 11410
rect 13800 11330 13810 11390
rect 13870 11330 13880 11390
rect 13800 11310 13880 11330
rect 13800 11250 13810 11310
rect 13870 11250 13880 11310
rect 13800 11240 13880 11250
rect 14040 11470 14120 11480
rect 14040 11410 14050 11470
rect 14110 11410 14120 11470
rect 14040 11390 14120 11410
rect 14040 11330 14050 11390
rect 14110 11330 14120 11390
rect 14040 11310 14120 11330
rect 14040 11250 14050 11310
rect 14110 11250 14120 11310
rect 14040 11240 14120 11250
rect 14280 11470 14360 11480
rect 14280 11410 14290 11470
rect 14350 11410 14360 11470
rect 14280 11390 14360 11410
rect 14280 11330 14290 11390
rect 14350 11330 14360 11390
rect 14280 11310 14360 11330
rect 14280 11250 14290 11310
rect 14350 11250 14360 11310
rect 14280 11240 14360 11250
rect 14520 11470 14600 11480
rect 14520 11410 14530 11470
rect 14590 11410 14600 11470
rect 14520 11390 14600 11410
rect 14520 11330 14530 11390
rect 14590 11330 14600 11390
rect 14520 11310 14600 11330
rect 14520 11250 14530 11310
rect 14590 11250 14600 11310
rect 14520 11240 14600 11250
rect 14760 11470 14840 11480
rect 14760 11410 14770 11470
rect 14830 11410 14840 11470
rect 14760 11390 14840 11410
rect 14760 11330 14770 11390
rect 14830 11330 14840 11390
rect 14760 11310 14840 11330
rect 14760 11250 14770 11310
rect 14830 11250 14840 11310
rect 14760 11240 14840 11250
rect 15000 11470 15080 11480
rect 15000 11410 15010 11470
rect 15070 11410 15080 11470
rect 15000 11390 15080 11410
rect 15000 11330 15010 11390
rect 15070 11330 15080 11390
rect 15000 11310 15080 11330
rect 15000 11250 15010 11310
rect 15070 11250 15080 11310
rect 15000 11240 15080 11250
rect 15240 11470 15320 11480
rect 15240 11410 15250 11470
rect 15310 11410 15320 11470
rect 15240 11390 15320 11410
rect 15240 11330 15250 11390
rect 15310 11330 15320 11390
rect 15240 11310 15320 11330
rect 15240 11250 15250 11310
rect 15310 11250 15320 11310
rect 15240 11240 15320 11250
rect 15480 11470 15560 11480
rect 15480 11410 15490 11470
rect 15550 11410 15560 11470
rect 15480 11390 15560 11410
rect 15480 11330 15490 11390
rect 15550 11330 15560 11390
rect 15480 11310 15560 11330
rect 15480 11250 15490 11310
rect 15550 11250 15560 11310
rect 15480 11240 15560 11250
rect 15720 11470 15800 11480
rect 15720 11410 15730 11470
rect 15790 11410 15800 11470
rect 15720 11390 15800 11410
rect 15720 11330 15730 11390
rect 15790 11330 15800 11390
rect 15720 11310 15800 11330
rect 15720 11250 15730 11310
rect 15790 11250 15800 11310
rect 15720 11240 15800 11250
rect 14680 11200 14760 11210
rect 14680 11140 14690 11200
rect 14750 11140 14760 11200
rect 14680 11130 14760 11140
rect 14320 11090 14400 11100
rect 14320 11030 14330 11090
rect 14390 11030 14400 11090
rect 14320 11020 14400 11030
rect 13960 10980 14040 10990
rect 13960 10920 13970 10980
rect 14030 10920 14040 10980
rect 13960 10910 14040 10920
rect 13600 10870 13680 10880
rect 13600 10810 13610 10870
rect 13670 10810 13680 10870
rect 13600 10800 13680 10810
rect 13340 10760 13590 10770
rect 13400 10700 13430 10760
rect 13490 10700 13520 10760
rect 13580 10700 13590 10760
rect 13340 10690 13590 10700
rect 13620 10650 13660 10800
rect 13690 10760 13770 10770
rect 13690 10700 13700 10760
rect 13760 10700 13770 10760
rect 13690 10690 13770 10700
rect 13870 10760 13950 10770
rect 13870 10700 13880 10760
rect 13940 10700 13950 10760
rect 13870 10690 13950 10700
rect 13980 10650 14020 10910
rect 14050 10760 14130 10770
rect 14050 10700 14060 10760
rect 14120 10700 14130 10760
rect 14050 10690 14130 10700
rect 14230 10760 14310 10770
rect 14230 10700 14240 10760
rect 14300 10700 14310 10760
rect 14230 10690 14310 10700
rect 14340 10650 14380 11020
rect 14410 10760 14490 10770
rect 14410 10700 14420 10760
rect 14480 10700 14490 10760
rect 14410 10690 14490 10700
rect 14590 10760 14660 10770
rect 14590 10700 14600 10760
rect 14590 10690 14660 10700
rect 13250 10590 13260 10630
rect 13300 10590 13310 10630
rect 13250 10530 13310 10590
rect 13250 10490 13260 10530
rect 13300 10490 13310 10530
rect 13250 10430 13310 10490
rect 13250 10390 13260 10430
rect 13300 10390 13310 10430
rect 13250 10330 13310 10390
rect 13250 10290 13260 10330
rect 13300 10290 13310 10330
rect 13250 10230 13310 10290
rect 13250 10190 13260 10230
rect 13300 10190 13310 10230
rect 13250 10130 13310 10190
rect 13250 10090 13260 10130
rect 13300 10090 13310 10130
rect 13250 10070 13310 10090
rect 13430 10630 13490 10650
rect 13430 10590 13440 10630
rect 13480 10590 13490 10630
rect 13430 10530 13490 10590
rect 13430 10490 13440 10530
rect 13480 10490 13490 10530
rect 13430 10430 13490 10490
rect 13430 10390 13440 10430
rect 13480 10390 13490 10430
rect 13430 10330 13490 10390
rect 13430 10290 13440 10330
rect 13480 10290 13490 10330
rect 13430 10230 13490 10290
rect 13430 10190 13440 10230
rect 13480 10190 13490 10230
rect 13430 10130 13490 10190
rect 13430 10090 13440 10130
rect 13480 10090 13490 10130
rect 13430 10070 13490 10090
rect 13610 10630 13670 10650
rect 13610 10590 13620 10630
rect 13660 10590 13670 10630
rect 13610 10530 13670 10590
rect 13610 10490 13620 10530
rect 13660 10490 13670 10530
rect 13610 10430 13670 10490
rect 13610 10390 13620 10430
rect 13660 10390 13670 10430
rect 13610 10330 13670 10390
rect 13610 10290 13620 10330
rect 13660 10290 13670 10330
rect 13610 10230 13670 10290
rect 13610 10190 13620 10230
rect 13660 10190 13670 10230
rect 13610 10130 13670 10190
rect 13610 10090 13620 10130
rect 13660 10090 13670 10130
rect 13610 10070 13670 10090
rect 13790 10630 13850 10650
rect 13790 10590 13800 10630
rect 13840 10590 13850 10630
rect 13790 10530 13850 10590
rect 13790 10490 13800 10530
rect 13840 10490 13850 10530
rect 13790 10430 13850 10490
rect 13790 10390 13800 10430
rect 13840 10390 13850 10430
rect 13790 10330 13850 10390
rect 13790 10290 13800 10330
rect 13840 10290 13850 10330
rect 13790 10230 13850 10290
rect 13790 10190 13800 10230
rect 13840 10190 13850 10230
rect 13790 10130 13850 10190
rect 13790 10090 13800 10130
rect 13840 10090 13850 10130
rect 13790 10070 13850 10090
rect 13970 10630 14030 10650
rect 13970 10590 13980 10630
rect 14020 10590 14030 10630
rect 13970 10530 14030 10590
rect 13970 10490 13980 10530
rect 14020 10490 14030 10530
rect 13970 10430 14030 10490
rect 13970 10390 13980 10430
rect 14020 10390 14030 10430
rect 13970 10330 14030 10390
rect 13970 10290 13980 10330
rect 14020 10290 14030 10330
rect 13970 10230 14030 10290
rect 13970 10190 13980 10230
rect 14020 10190 14030 10230
rect 13970 10130 14030 10190
rect 13970 10090 13980 10130
rect 14020 10090 14030 10130
rect 13970 10070 14030 10090
rect 14150 10630 14210 10650
rect 14150 10590 14160 10630
rect 14200 10590 14210 10630
rect 14150 10530 14210 10590
rect 14150 10490 14160 10530
rect 14200 10490 14210 10530
rect 14150 10430 14210 10490
rect 14150 10390 14160 10430
rect 14200 10390 14210 10430
rect 14150 10330 14210 10390
rect 14150 10290 14160 10330
rect 14200 10290 14210 10330
rect 14150 10230 14210 10290
rect 14150 10190 14160 10230
rect 14200 10190 14210 10230
rect 14150 10130 14210 10190
rect 14150 10090 14160 10130
rect 14200 10090 14210 10130
rect 14150 10070 14210 10090
rect 14330 10630 14390 10650
rect 14330 10590 14340 10630
rect 14380 10590 14390 10630
rect 14330 10530 14390 10590
rect 14330 10490 14340 10530
rect 14380 10490 14390 10530
rect 14330 10430 14390 10490
rect 14330 10390 14340 10430
rect 14380 10390 14390 10430
rect 14330 10330 14390 10390
rect 14330 10290 14340 10330
rect 14380 10290 14390 10330
rect 14330 10230 14390 10290
rect 14330 10190 14340 10230
rect 14380 10190 14390 10230
rect 14330 10130 14390 10190
rect 14330 10090 14340 10130
rect 14380 10090 14390 10130
rect 14330 10070 14390 10090
rect 14510 10630 14570 10650
rect 14510 10590 14520 10630
rect 14560 10590 14570 10630
rect 14510 10530 14570 10590
rect 14510 10490 14520 10530
rect 14560 10490 14570 10530
rect 14510 10430 14570 10490
rect 14510 10390 14520 10430
rect 14560 10390 14570 10430
rect 14510 10330 14570 10390
rect 14510 10290 14520 10330
rect 14560 10290 14570 10330
rect 14510 10230 14570 10290
rect 14510 10190 14520 10230
rect 14560 10190 14570 10230
rect 14510 10130 14570 10190
rect 14510 10090 14520 10130
rect 14560 10090 14570 10130
rect 14510 10070 14570 10090
rect 14690 10630 14750 11130
rect 15710 11090 15790 11100
rect 15710 11030 15720 11090
rect 15780 11030 15790 11090
rect 15240 10980 15320 10990
rect 15240 10920 15250 10980
rect 15310 10920 15320 10980
rect 15240 10910 15320 10920
rect 14690 10590 14700 10630
rect 14740 10590 14750 10630
rect 14690 10530 14750 10590
rect 14690 10490 14700 10530
rect 14740 10490 14750 10530
rect 14690 10430 14750 10490
rect 14690 10390 14700 10430
rect 14740 10390 14750 10430
rect 14690 10330 14750 10390
rect 14690 10290 14700 10330
rect 14740 10290 14750 10330
rect 14690 10230 14750 10290
rect 14690 10190 14700 10230
rect 14740 10190 14750 10230
rect 14690 10130 14750 10190
rect 14690 10090 14700 10130
rect 14740 10090 14750 10130
rect 14690 10070 14750 10090
rect 14870 10630 14930 10650
rect 14870 10590 14880 10630
rect 14920 10590 14930 10630
rect 14870 10530 14930 10590
rect 14870 10490 14880 10530
rect 14920 10490 14930 10530
rect 14870 10430 14930 10490
rect 14870 10390 14880 10430
rect 14920 10390 14930 10430
rect 14870 10330 14930 10390
rect 14870 10290 14880 10330
rect 14920 10290 14930 10330
rect 14870 10230 14930 10290
rect 15260 10230 15300 10910
rect 15590 10560 15670 10570
rect 15590 10500 15600 10560
rect 15660 10500 15670 10560
rect 15590 10490 15670 10500
rect 15710 10550 15790 11030
rect 15840 10570 15920 11520
rect 15970 11570 16030 11650
rect 15970 11530 15980 11570
rect 16020 11530 16030 11570
rect 15970 11480 16030 11530
rect 15960 11470 16040 11480
rect 15960 11410 15970 11470
rect 16030 11410 16040 11470
rect 15960 11390 16040 11410
rect 15960 11330 15970 11390
rect 16030 11330 16040 11390
rect 15960 11310 16040 11330
rect 15960 11250 15970 11310
rect 16030 11250 16040 11310
rect 15960 11240 16040 11250
rect 16170 10880 16210 12680
rect 16260 12530 16300 14730
rect 16240 12520 16320 12530
rect 16240 12460 16250 12520
rect 16310 12460 16320 12520
rect 16240 12450 16320 12460
rect 16260 10990 16300 12450
rect 16350 12200 16590 15290
rect 16780 14490 16860 17441
rect 16780 14430 16790 14490
rect 16850 14430 16860 14490
rect 16780 14420 16860 14430
rect 17570 17631 17650 17650
rect 17570 17234 17590 17631
rect 17628 17234 17650 17631
rect 17570 16750 17650 17234
rect 17570 16690 17580 16750
rect 17640 16690 17650 16750
rect 16350 12140 16360 12200
rect 16420 12140 16440 12200
rect 16500 12140 16520 12200
rect 16580 12140 16590 12200
rect 16350 12120 16590 12140
rect 16350 12060 16360 12120
rect 16420 12060 16440 12120
rect 16500 12060 16520 12120
rect 16580 12060 16590 12120
rect 16350 12040 16590 12060
rect 16350 11980 16360 12040
rect 16420 11980 16440 12040
rect 16500 11980 16520 12040
rect 16580 11980 16590 12040
rect 16350 11970 16590 11980
rect 17570 11580 17650 16690
rect 17950 16050 18030 18050
rect 17950 15990 17960 16050
rect 18020 15990 18030 16050
rect 17950 15980 18030 15990
rect 18120 17450 18200 17460
rect 18120 17390 18130 17450
rect 18190 17390 18200 17450
rect 18120 13440 18200 17390
rect 18650 14380 18730 18070
rect 18780 16750 18880 16770
rect 18780 16690 18800 16750
rect 18860 16690 18880 16750
rect 18780 16670 18880 16690
rect 18780 15350 18880 15370
rect 18780 15290 18800 15350
rect 18860 15290 18880 15350
rect 18780 15270 18880 15290
rect 18650 14320 18660 14380
rect 18720 14320 18730 14380
rect 18650 14310 18730 14320
rect 17570 11520 17580 11580
rect 17640 11520 17650 11580
rect 17570 11510 17650 11520
rect 16240 10980 16320 10990
rect 16240 10920 16250 10980
rect 16310 10920 16320 10980
rect 16240 10910 16320 10920
rect 16150 10870 16230 10880
rect 16150 10810 16160 10870
rect 16220 10810 16230 10870
rect 16150 10800 16230 10810
rect 15710 10510 15730 10550
rect 15770 10510 15790 10550
rect 15710 10490 15790 10510
rect 15830 10560 15910 10570
rect 15830 10500 15840 10560
rect 15900 10500 15910 10560
rect 15830 10490 15910 10500
rect 15500 10430 15560 10450
rect 15500 10390 15510 10430
rect 15550 10390 15560 10430
rect 15500 10330 15560 10390
rect 15500 10290 15510 10330
rect 15550 10290 15560 10330
rect 15500 10230 15560 10290
rect 15610 10430 15670 10490
rect 15610 10390 15620 10430
rect 15660 10390 15670 10430
rect 15610 10330 15670 10390
rect 15610 10290 15620 10330
rect 15660 10290 15670 10330
rect 15610 10270 15670 10290
rect 15720 10430 15780 10450
rect 15720 10390 15730 10430
rect 15770 10390 15780 10430
rect 15720 10330 15780 10390
rect 15720 10290 15730 10330
rect 15770 10290 15780 10330
rect 15720 10230 15780 10290
rect 15830 10430 15890 10490
rect 15830 10390 15840 10430
rect 15880 10390 15890 10430
rect 15830 10330 15890 10390
rect 15830 10290 15840 10330
rect 15880 10290 15890 10330
rect 15830 10270 15890 10290
rect 15940 10430 16000 10450
rect 15940 10390 15950 10430
rect 15990 10390 16000 10430
rect 15940 10330 16000 10390
rect 15940 10290 15950 10330
rect 15990 10290 16000 10330
rect 15940 10230 16000 10290
rect 14870 10190 14880 10230
rect 14920 10190 14930 10230
rect 14870 10130 14930 10190
rect 15240 10220 15320 10230
rect 15240 10160 15250 10220
rect 15310 10160 15320 10220
rect 15240 10150 15320 10160
rect 15490 10210 15570 10230
rect 15490 10170 15510 10210
rect 15550 10170 15570 10210
rect 15490 10150 15570 10170
rect 15710 10220 15790 10230
rect 15710 10160 15720 10220
rect 15780 10160 15790 10220
rect 15710 10150 15790 10160
rect 15930 10210 16010 10230
rect 15930 10170 15950 10210
rect 15990 10170 16010 10210
rect 15930 10150 16010 10170
rect 14870 10090 14880 10130
rect 14920 10090 14930 10130
rect 14870 10070 14930 10090
rect 15500 10030 15560 10150
rect 15940 10030 16000 10150
rect 11620 10020 11700 10030
rect 11620 9960 11630 10020
rect 11690 9960 11700 10020
rect 11620 9940 11700 9960
rect 11620 9880 11630 9940
rect 11690 9880 11700 9940
rect 11620 9860 11700 9880
rect 11620 9800 11630 9860
rect 11690 9800 11700 9860
rect 11620 9790 11700 9800
rect 11980 10020 12060 10030
rect 11980 9960 11990 10020
rect 12050 9960 12060 10020
rect 11980 9940 12060 9960
rect 11980 9880 11990 9940
rect 12050 9880 12060 9940
rect 11980 9860 12060 9880
rect 11980 9800 11990 9860
rect 12050 9800 12060 9860
rect 11980 9790 12060 9800
rect 12340 10020 12420 10030
rect 12340 9960 12350 10020
rect 12410 9960 12420 10020
rect 12340 9940 12420 9960
rect 12340 9880 12350 9940
rect 12410 9880 12420 9940
rect 12340 9860 12420 9880
rect 12340 9800 12350 9860
rect 12410 9800 12420 9860
rect 12340 9790 12420 9800
rect 12700 10020 12780 10030
rect 12700 9960 12710 10020
rect 12770 9960 12780 10020
rect 12700 9940 12780 9960
rect 12700 9880 12710 9940
rect 12770 9880 12780 9940
rect 12700 9860 12780 9880
rect 12700 9800 12710 9860
rect 12770 9800 12780 9860
rect 12700 9790 12780 9800
rect 13060 10020 13140 10030
rect 13060 9960 13070 10020
rect 13130 9960 13140 10020
rect 13060 9940 13140 9960
rect 13060 9880 13070 9940
rect 13130 9880 13140 9940
rect 13060 9860 13140 9880
rect 13060 9800 13070 9860
rect 13130 9800 13140 9860
rect 13060 9790 13140 9800
rect 13420 10020 13500 10030
rect 13420 9960 13430 10020
rect 13490 9960 13500 10020
rect 13420 9940 13500 9960
rect 13420 9880 13430 9940
rect 13490 9880 13500 9940
rect 13420 9860 13500 9880
rect 13420 9800 13430 9860
rect 13490 9800 13500 9860
rect 13420 9790 13500 9800
rect 13780 10020 13860 10030
rect 13780 9960 13790 10020
rect 13850 9960 13860 10020
rect 13780 9940 13860 9960
rect 13780 9880 13790 9940
rect 13850 9880 13860 9940
rect 13780 9860 13860 9880
rect 13780 9800 13790 9860
rect 13850 9800 13860 9860
rect 13780 9790 13860 9800
rect 14140 10020 14220 10030
rect 14140 9960 14150 10020
rect 14210 9960 14220 10020
rect 14140 9940 14220 9960
rect 14140 9880 14150 9940
rect 14210 9880 14220 9940
rect 14140 9860 14220 9880
rect 14140 9800 14150 9860
rect 14210 9800 14220 9860
rect 14140 9790 14220 9800
rect 14500 10020 14580 10030
rect 14500 9960 14510 10020
rect 14570 9960 14580 10020
rect 14500 9940 14580 9960
rect 14500 9880 14510 9940
rect 14570 9880 14580 9940
rect 14500 9860 14580 9880
rect 14500 9800 14510 9860
rect 14570 9800 14580 9860
rect 14500 9790 14580 9800
rect 14860 10020 14940 10030
rect 14860 9960 14870 10020
rect 14930 9960 14940 10020
rect 14860 9940 14940 9960
rect 14860 9880 14870 9940
rect 14930 9880 14940 9940
rect 14860 9860 14940 9880
rect 14860 9800 14870 9860
rect 14930 9800 14940 9860
rect 14860 9790 14940 9800
rect 15490 10020 15570 10030
rect 15490 9960 15500 10020
rect 15560 9960 15570 10020
rect 15490 9940 15570 9960
rect 15490 9880 15500 9940
rect 15560 9880 15570 9940
rect 15490 9860 15570 9880
rect 15490 9800 15500 9860
rect 15560 9800 15570 9860
rect 15490 9790 15570 9800
rect 15930 10020 16010 10030
rect 15930 9960 15940 10020
rect 16000 9960 16010 10020
rect 15930 9940 16010 9960
rect 15930 9880 15940 9940
rect 16000 9880 16010 9940
rect 15930 9860 16010 9880
rect 15930 9800 15940 9860
rect 16000 9800 16010 9860
rect 15930 9790 16010 9800
rect 11806 9750 11864 9760
rect 11806 9698 11808 9750
rect 11860 9698 11864 9750
rect 11806 9690 11864 9698
rect 11916 9750 11974 9760
rect 11916 9698 11918 9750
rect 11970 9698 11974 9750
rect 11916 9690 11974 9698
rect 12026 9750 12084 9760
rect 12026 9698 12028 9750
rect 12080 9698 12084 9750
rect 12026 9690 12084 9698
rect 12136 9750 12194 9760
rect 12136 9698 12138 9750
rect 12190 9698 12194 9750
rect 12136 9690 12194 9698
rect 12246 9750 12304 9760
rect 12246 9698 12248 9750
rect 12300 9698 12304 9750
rect 12246 9690 12304 9698
rect 12356 9750 12414 9760
rect 12356 9698 12358 9750
rect 12410 9698 12414 9750
rect 12356 9690 12414 9698
rect 12466 9750 12524 9760
rect 12466 9698 12468 9750
rect 12520 9698 12524 9750
rect 12466 9690 12524 9698
rect 12576 9750 12634 9760
rect 12576 9698 12578 9750
rect 12630 9698 12634 9750
rect 12576 9690 12634 9698
rect 12686 9750 12744 9760
rect 12686 9698 12688 9750
rect 12740 9698 12744 9750
rect 12686 9690 12744 9698
rect 12796 9750 12854 9760
rect 12796 9698 12798 9750
rect 12850 9698 12854 9750
rect 12796 9690 12854 9698
rect 13706 9750 13764 9760
rect 13706 9698 13708 9750
rect 13760 9698 13764 9750
rect 13706 9690 13764 9698
rect 13816 9750 13874 9760
rect 13816 9698 13818 9750
rect 13870 9698 13874 9750
rect 13816 9690 13874 9698
rect 13926 9750 13984 9760
rect 13926 9698 13928 9750
rect 13980 9698 13984 9750
rect 13926 9690 13984 9698
rect 14036 9750 14094 9760
rect 14036 9698 14038 9750
rect 14090 9698 14094 9750
rect 14036 9690 14094 9698
rect 14146 9750 14204 9760
rect 14146 9698 14148 9750
rect 14200 9698 14204 9750
rect 14146 9690 14204 9698
rect 14256 9750 14314 9760
rect 14256 9698 14258 9750
rect 14310 9698 14314 9750
rect 14256 9690 14314 9698
rect 14366 9750 14424 9760
rect 14366 9698 14368 9750
rect 14420 9698 14424 9750
rect 14366 9690 14424 9698
rect 14476 9750 14534 9760
rect 14476 9698 14478 9750
rect 14530 9698 14534 9750
rect 14476 9690 14534 9698
rect 14586 9750 14644 9760
rect 14586 9698 14588 9750
rect 14640 9698 14644 9750
rect 14586 9690 14644 9698
rect 14696 9750 14754 9760
rect 14696 9698 14698 9750
rect 14750 9698 14754 9750
rect 14696 9690 14754 9698
rect 11560 9630 11700 9650
rect 11560 9590 11570 9630
rect 11610 9590 11650 9630
rect 11690 9590 11700 9630
rect 11560 9530 11700 9590
rect 11560 9490 11570 9530
rect 11610 9490 11650 9530
rect 11690 9490 11700 9530
rect 11560 9470 11700 9490
rect 11640 9430 11700 9470
rect 11750 9630 11810 9650
rect 11750 9590 11760 9630
rect 11800 9590 11810 9630
rect 11750 9530 11810 9590
rect 11750 9490 11760 9530
rect 11800 9490 11810 9530
rect 11630 9420 11710 9430
rect 11630 9360 11640 9420
rect 11700 9360 11710 9420
rect 11630 9350 11710 9360
rect 11750 9320 11810 9490
rect 11860 9630 11920 9650
rect 11860 9590 11870 9630
rect 11910 9590 11920 9630
rect 11860 9530 11920 9590
rect 11860 9490 11870 9530
rect 11910 9490 11920 9530
rect 11860 9430 11920 9490
rect 11970 9630 12030 9650
rect 11970 9590 11980 9630
rect 12020 9590 12030 9630
rect 11970 9530 12030 9590
rect 11970 9490 11980 9530
rect 12020 9490 12030 9530
rect 11850 9420 11930 9430
rect 11850 9360 11860 9420
rect 11920 9360 11930 9420
rect 11850 9350 11930 9360
rect 11970 9320 12030 9490
rect 12080 9630 12140 9650
rect 12080 9590 12090 9630
rect 12130 9590 12140 9630
rect 12080 9530 12140 9590
rect 12080 9490 12090 9530
rect 12130 9490 12140 9530
rect 12080 9430 12140 9490
rect 12190 9630 12250 9650
rect 12190 9590 12200 9630
rect 12240 9590 12250 9630
rect 12190 9530 12250 9590
rect 12190 9490 12200 9530
rect 12240 9490 12250 9530
rect 12070 9420 12150 9430
rect 12070 9360 12080 9420
rect 12140 9360 12150 9420
rect 12070 9350 12150 9360
rect 12190 9320 12250 9490
rect 12300 9630 12360 9650
rect 12300 9590 12310 9630
rect 12350 9590 12360 9630
rect 12300 9530 12360 9590
rect 12300 9490 12310 9530
rect 12350 9490 12360 9530
rect 12300 9430 12360 9490
rect 12410 9630 12470 9650
rect 12410 9590 12420 9630
rect 12460 9590 12470 9630
rect 12410 9530 12470 9590
rect 12410 9490 12420 9530
rect 12460 9490 12470 9530
rect 12290 9420 12370 9430
rect 12290 9360 12300 9420
rect 12360 9360 12370 9420
rect 12290 9350 12370 9360
rect 12410 9320 12470 9490
rect 12520 9630 12580 9650
rect 12520 9590 12530 9630
rect 12570 9590 12580 9630
rect 12520 9530 12580 9590
rect 12520 9490 12530 9530
rect 12570 9490 12580 9530
rect 12520 9430 12580 9490
rect 12630 9630 12690 9650
rect 12630 9590 12640 9630
rect 12680 9590 12690 9630
rect 12630 9530 12690 9590
rect 12630 9490 12640 9530
rect 12680 9490 12690 9530
rect 12510 9420 12590 9430
rect 12510 9360 12520 9420
rect 12580 9360 12590 9420
rect 12510 9350 12590 9360
rect 12630 9320 12690 9490
rect 12740 9630 12800 9650
rect 12740 9590 12750 9630
rect 12790 9590 12800 9630
rect 12740 9530 12800 9590
rect 12740 9490 12750 9530
rect 12790 9490 12800 9530
rect 12740 9430 12800 9490
rect 12850 9630 12910 9650
rect 12850 9590 12860 9630
rect 12900 9590 12910 9630
rect 12850 9530 12910 9590
rect 12850 9490 12860 9530
rect 12900 9490 12910 9530
rect 12730 9420 12810 9430
rect 12730 9360 12740 9420
rect 12800 9360 12810 9420
rect 12730 9350 12810 9360
rect 12850 9320 12910 9490
rect 12960 9630 13100 9650
rect 12960 9590 12970 9630
rect 13010 9590 13050 9630
rect 13090 9590 13100 9630
rect 12960 9530 13100 9590
rect 12960 9490 12970 9530
rect 13010 9490 13050 9530
rect 13090 9490 13100 9530
rect 12960 9470 13100 9490
rect 13460 9630 13600 9650
rect 13460 9590 13470 9630
rect 13510 9590 13550 9630
rect 13590 9590 13600 9630
rect 13460 9530 13600 9590
rect 13460 9490 13470 9530
rect 13510 9490 13550 9530
rect 13590 9490 13600 9530
rect 13460 9470 13600 9490
rect 12960 9430 13020 9470
rect 13540 9430 13600 9470
rect 13650 9630 13710 9650
rect 13650 9590 13660 9630
rect 13700 9590 13710 9630
rect 13650 9530 13710 9590
rect 13650 9490 13660 9530
rect 13700 9490 13710 9530
rect 12950 9420 13030 9430
rect 12950 9360 12960 9420
rect 13020 9360 13030 9420
rect 12950 9350 13030 9360
rect 13530 9420 13610 9430
rect 13530 9360 13540 9420
rect 13600 9360 13610 9420
rect 13530 9350 13610 9360
rect 9680 9250 9690 9310
rect 9750 9250 9760 9310
rect 9680 9240 9760 9250
rect 11740 9310 11820 9320
rect 11740 9250 11750 9310
rect 11810 9250 11820 9310
rect 11740 9240 11820 9250
rect 11960 9310 12040 9320
rect 11960 9250 11970 9310
rect 12030 9250 12040 9310
rect 11960 9240 12040 9250
rect 12180 9310 12260 9320
rect 12180 9250 12190 9310
rect 12250 9250 12260 9310
rect 12180 9240 12260 9250
rect 12400 9310 12480 9320
rect 12400 9250 12410 9310
rect 12470 9250 12480 9310
rect 12400 9240 12480 9250
rect 12620 9310 12700 9320
rect 12620 9250 12630 9310
rect 12690 9250 12700 9310
rect 12620 9240 12700 9250
rect 12840 9310 12920 9320
rect 13650 9310 13710 9490
rect 13760 9630 13820 9650
rect 13760 9590 13770 9630
rect 13810 9590 13820 9630
rect 13760 9530 13820 9590
rect 13760 9490 13770 9530
rect 13810 9490 13820 9530
rect 13760 9430 13820 9490
rect 13870 9630 13930 9650
rect 13870 9590 13880 9630
rect 13920 9590 13930 9630
rect 13870 9530 13930 9590
rect 13870 9490 13880 9530
rect 13920 9490 13930 9530
rect 13750 9420 13830 9430
rect 13750 9360 13760 9420
rect 13820 9360 13830 9420
rect 13750 9350 13830 9360
rect 13870 9310 13930 9490
rect 13980 9630 14040 9650
rect 13980 9590 13990 9630
rect 14030 9590 14040 9630
rect 13980 9530 14040 9590
rect 13980 9490 13990 9530
rect 14030 9490 14040 9530
rect 13980 9430 14040 9490
rect 14090 9630 14150 9650
rect 14090 9590 14100 9630
rect 14140 9590 14150 9630
rect 14090 9530 14150 9590
rect 14090 9490 14100 9530
rect 14140 9490 14150 9530
rect 13970 9420 14050 9430
rect 13970 9360 13980 9420
rect 14040 9360 14050 9420
rect 13970 9350 14050 9360
rect 14090 9310 14150 9490
rect 14200 9630 14260 9650
rect 14200 9590 14210 9630
rect 14250 9590 14260 9630
rect 14200 9530 14260 9590
rect 14200 9490 14210 9530
rect 14250 9490 14260 9530
rect 14200 9430 14260 9490
rect 14310 9630 14370 9650
rect 14310 9590 14320 9630
rect 14360 9590 14370 9630
rect 14310 9530 14370 9590
rect 14310 9490 14320 9530
rect 14360 9490 14370 9530
rect 14190 9420 14270 9430
rect 14190 9360 14200 9420
rect 14260 9360 14270 9420
rect 14190 9350 14270 9360
rect 14310 9310 14370 9490
rect 14420 9630 14480 9650
rect 14420 9590 14430 9630
rect 14470 9590 14480 9630
rect 14420 9530 14480 9590
rect 14420 9490 14430 9530
rect 14470 9490 14480 9530
rect 14420 9430 14480 9490
rect 14530 9630 14590 9650
rect 14530 9590 14540 9630
rect 14580 9590 14590 9630
rect 14530 9530 14590 9590
rect 14530 9490 14540 9530
rect 14580 9490 14590 9530
rect 14410 9420 14490 9430
rect 14410 9360 14420 9420
rect 14480 9360 14490 9420
rect 14410 9350 14490 9360
rect 14530 9310 14590 9490
rect 14640 9630 14700 9650
rect 14640 9590 14650 9630
rect 14690 9590 14700 9630
rect 14640 9530 14700 9590
rect 14640 9490 14650 9530
rect 14690 9490 14700 9530
rect 14640 9430 14700 9490
rect 14750 9630 14810 9650
rect 14750 9590 14760 9630
rect 14800 9590 14810 9630
rect 14750 9530 14810 9590
rect 14750 9490 14760 9530
rect 14800 9490 14810 9530
rect 14630 9420 14710 9430
rect 14630 9360 14640 9420
rect 14700 9360 14710 9420
rect 14630 9350 14710 9360
rect 14750 9310 14810 9490
rect 14860 9630 15000 9650
rect 14860 9590 14870 9630
rect 14910 9590 14950 9630
rect 14990 9590 15000 9630
rect 14860 9530 15000 9590
rect 14860 9490 14870 9530
rect 14910 9490 14950 9530
rect 14990 9490 15000 9530
rect 14860 9470 15000 9490
rect 14860 9430 14920 9470
rect 14850 9420 14930 9430
rect 14850 9360 14860 9420
rect 14920 9360 14930 9420
rect 14850 9350 14930 9360
rect 12840 9250 12850 9310
rect 12910 9250 12920 9310
rect 12840 9240 12920 9250
rect 13640 9300 13720 9310
rect 13640 9240 13650 9300
rect 13710 9240 13720 9300
rect 13640 9220 13720 9240
rect 13640 9160 13650 9220
rect 13710 9160 13720 9220
rect 13640 9140 13720 9160
rect 13640 9080 13650 9140
rect 13710 9080 13720 9140
rect 13640 9070 13720 9080
rect 13860 9300 13940 9310
rect 13860 9240 13870 9300
rect 13930 9240 13940 9300
rect 13860 9220 13940 9240
rect 13860 9160 13870 9220
rect 13930 9160 13940 9220
rect 13860 9140 13940 9160
rect 13860 9080 13870 9140
rect 13930 9080 13940 9140
rect 13860 9070 13940 9080
rect 14080 9300 14160 9310
rect 14080 9240 14090 9300
rect 14150 9240 14160 9300
rect 14080 9220 14160 9240
rect 14080 9160 14090 9220
rect 14150 9160 14160 9220
rect 14080 9140 14160 9160
rect 14080 9080 14090 9140
rect 14150 9080 14160 9140
rect 14080 9070 14160 9080
rect 14300 9300 14380 9310
rect 14300 9240 14310 9300
rect 14370 9240 14380 9300
rect 14300 9220 14380 9240
rect 14300 9160 14310 9220
rect 14370 9160 14380 9220
rect 14300 9140 14380 9160
rect 14300 9080 14310 9140
rect 14370 9080 14380 9140
rect 14300 9070 14380 9080
rect 14520 9300 14600 9310
rect 14520 9240 14530 9300
rect 14590 9240 14600 9300
rect 14520 9220 14600 9240
rect 14520 9160 14530 9220
rect 14590 9160 14600 9220
rect 14520 9140 14600 9160
rect 14520 9080 14530 9140
rect 14590 9080 14600 9140
rect 14520 9070 14600 9080
rect 14740 9300 14820 9310
rect 14740 9240 14750 9300
rect 14810 9240 14820 9300
rect 14740 9220 14820 9240
rect 14740 9160 14750 9220
rect 14810 9160 14820 9220
rect 14740 9140 14820 9160
rect 14740 9080 14750 9140
rect 14810 9080 14820 9140
rect 14740 9070 14820 9080
<< via1 >>
rect 8880 19130 8940 19190
rect 8460 19020 8520 19080
rect 8460 18940 8520 19000
rect 8460 18860 8520 18920
rect 8460 18043 8470 18440
rect 8470 18043 8508 18440
rect 8508 18043 8520 18440
rect 8460 18040 8520 18043
rect 8880 18390 8940 18450
rect 8880 18310 8940 18370
rect 8880 18220 8940 18280
rect 8880 18130 8940 18190
rect 8880 18050 8940 18110
rect 9250 19020 9310 19080
rect 9250 18940 9310 19000
rect 9250 18860 9310 18920
rect 10690 19020 10750 19080
rect 10690 18940 10750 19000
rect 10690 18860 10750 18920
rect 8460 11520 8520 11580
rect 9470 14150 9530 14210
rect 10360 14660 10420 14720
rect 9580 12460 9640 12520
rect 9580 11140 9640 11200
rect 9690 14430 9750 14490
rect 9690 12690 9750 12750
rect 9470 11030 9530 11090
rect 8460 9700 8520 9760
rect 10630 14320 10690 14380
rect 18200 19130 18260 19190
rect 13250 19070 13310 19080
rect 13250 19030 13260 19070
rect 13260 19030 13300 19070
rect 13300 19030 13310 19070
rect 13250 19020 13310 19030
rect 13250 18990 13310 19000
rect 13250 18950 13260 18990
rect 13260 18950 13300 18990
rect 13300 18950 13310 18990
rect 13250 18940 13310 18950
rect 13250 18910 13310 18920
rect 13250 18870 13260 18910
rect 13260 18870 13300 18910
rect 13300 18870 13310 18910
rect 13250 18860 13310 18870
rect 15680 19020 15740 19080
rect 15680 18940 15740 19000
rect 15680 18860 15740 18920
rect 16790 19020 16850 19080
rect 16790 18940 16850 19000
rect 16790 18860 16850 18920
rect 17580 19020 17640 19080
rect 17580 18940 17640 19000
rect 17580 18860 17640 18920
rect 18200 18790 18260 18850
rect 17580 18043 17590 18440
rect 17590 18043 17628 18440
rect 17628 18043 17640 18440
rect 17580 18040 17640 18043
rect 17960 18390 18020 18450
rect 17960 18310 18020 18370
rect 17960 18220 18020 18280
rect 17960 18130 18020 18190
rect 17960 18050 18020 18110
rect 18660 18090 18720 18150
rect 11150 16750 11210 16810
rect 11580 16750 11640 16810
rect 13250 16754 13310 16810
rect 13250 16750 13254 16754
rect 13254 16750 13310 16754
rect 15350 16750 15410 16810
rect 15350 14740 15410 14800
rect 16360 15290 16420 15350
rect 16440 15290 16500 15350
rect 16520 15290 16580 15350
rect 16010 14740 16070 14800
rect 16250 14740 16310 14800
rect 13960 14660 14020 14720
rect 11150 14550 11210 14610
rect 12552 14600 12622 14610
rect 12552 14550 12562 14600
rect 12562 14550 12612 14600
rect 12612 14550 12622 14600
rect 12552 14540 12622 14550
rect 13950 14600 14020 14610
rect 13950 14550 13960 14600
rect 13960 14550 14010 14600
rect 14010 14550 14020 14600
rect 13950 14540 14020 14550
rect 16160 14540 16220 14600
rect 11040 14320 11100 14380
rect 11090 14200 11150 14210
rect 11090 14160 11100 14200
rect 11100 14160 11140 14200
rect 11140 14160 11150 14200
rect 11090 14150 11150 14160
rect 15480 14240 15540 14250
rect 15480 14200 15490 14240
rect 15490 14200 15530 14240
rect 15530 14200 15540 14240
rect 15480 14190 15540 14200
rect 15480 14160 15540 14170
rect 15480 14120 15490 14160
rect 15490 14120 15530 14160
rect 15530 14120 15540 14160
rect 15480 14110 15540 14120
rect 11170 14030 11230 14040
rect 11170 13990 11180 14030
rect 11180 13990 11220 14030
rect 11220 13990 11230 14030
rect 11170 13980 11230 13990
rect 11330 14030 11390 14040
rect 11330 13990 11340 14030
rect 11340 13990 11380 14030
rect 11380 13990 11390 14030
rect 11330 13980 11390 13990
rect 11490 14030 11550 14040
rect 11490 13990 11500 14030
rect 11500 13990 11540 14030
rect 11540 13990 11550 14030
rect 11490 13980 11550 13990
rect 11650 14030 11710 14040
rect 11650 13990 11660 14030
rect 11660 13990 11700 14030
rect 11700 13990 11710 14030
rect 11650 13980 11710 13990
rect 11810 14030 11870 14040
rect 11810 13990 11820 14030
rect 11820 13990 11860 14030
rect 11860 13990 11870 14030
rect 11810 13980 11870 13990
rect 11970 14030 12030 14040
rect 11970 13990 11980 14030
rect 11980 13990 12020 14030
rect 12020 13990 12030 14030
rect 11970 13980 12030 13990
rect 12130 14030 12190 14040
rect 12130 13990 12140 14030
rect 12140 13990 12180 14030
rect 12180 13990 12190 14030
rect 12130 13980 12190 13990
rect 12290 14030 12350 14040
rect 12290 13990 12300 14030
rect 12300 13990 12340 14030
rect 12340 13990 12350 14030
rect 12290 13980 12350 13990
rect 12450 14030 12510 14040
rect 12450 13990 12460 14030
rect 12460 13990 12500 14030
rect 12500 13990 12510 14030
rect 12450 13980 12510 13990
rect 12610 14030 12670 14040
rect 12610 13990 12620 14030
rect 12620 13990 12660 14030
rect 12660 13990 12670 14030
rect 12610 13980 12670 13990
rect 12770 14030 12830 14040
rect 12770 13990 12780 14030
rect 12780 13990 12820 14030
rect 12820 13990 12830 14030
rect 12770 13980 12830 13990
rect 12930 14030 12990 14040
rect 12930 13990 12940 14030
rect 12940 13990 12980 14030
rect 12980 13990 12990 14030
rect 12930 13980 12990 13990
rect 13090 14030 13150 14040
rect 13090 13990 13100 14030
rect 13100 13990 13140 14030
rect 13140 13990 13150 14030
rect 13090 13980 13150 13990
rect 13250 14030 13310 14040
rect 13250 13990 13260 14030
rect 13260 13990 13300 14030
rect 13300 13990 13310 14030
rect 13250 13980 13310 13990
rect 13410 14030 13470 14040
rect 13410 13990 13420 14030
rect 13420 13990 13460 14030
rect 13460 13990 13470 14030
rect 13410 13980 13470 13990
rect 13570 14030 13630 14040
rect 13570 13990 13580 14030
rect 13580 13990 13620 14030
rect 13620 13990 13630 14030
rect 13570 13980 13630 13990
rect 13730 14030 13790 14040
rect 13730 13990 13740 14030
rect 13740 13990 13780 14030
rect 13780 13990 13790 14030
rect 13730 13980 13790 13990
rect 13890 14030 13950 14040
rect 13890 13990 13900 14030
rect 13900 13990 13940 14030
rect 13940 13990 13950 14030
rect 13890 13980 13950 13990
rect 14050 14030 14110 14040
rect 14050 13990 14060 14030
rect 14060 13990 14100 14030
rect 14100 13990 14110 14030
rect 14050 13980 14110 13990
rect 14210 14030 14270 14040
rect 14210 13990 14220 14030
rect 14220 13990 14260 14030
rect 14260 13990 14270 14030
rect 14210 13980 14270 13990
rect 14370 14030 14430 14040
rect 14370 13990 14380 14030
rect 14380 13990 14420 14030
rect 14420 13990 14430 14030
rect 14370 13980 14430 13990
rect 14530 14030 14590 14040
rect 14530 13990 14540 14030
rect 14540 13990 14580 14030
rect 14580 13990 14590 14030
rect 14530 13980 14590 13990
rect 14690 14030 14750 14040
rect 14690 13990 14700 14030
rect 14700 13990 14740 14030
rect 14740 13990 14750 14030
rect 14690 13980 14750 13990
rect 14850 14030 14910 14040
rect 14850 13990 14860 14030
rect 14860 13990 14900 14030
rect 14900 13990 14910 14030
rect 14850 13980 14910 13990
rect 15010 14030 15070 14040
rect 15010 13990 15020 14030
rect 15020 13990 15060 14030
rect 15060 13990 15070 14030
rect 15010 13980 15070 13990
rect 15170 14030 15230 14040
rect 15170 13990 15180 14030
rect 15180 13990 15220 14030
rect 15220 13990 15230 14030
rect 15170 13980 15230 13990
rect 11910 13870 11970 13930
rect 11910 13790 11970 13850
rect 11910 13760 11970 13770
rect 11910 13720 11920 13760
rect 11920 13720 11960 13760
rect 11960 13720 11970 13760
rect 11910 13710 11970 13720
rect 13170 13870 13230 13930
rect 13250 13870 13310 13930
rect 13330 13870 13390 13930
rect 13170 13790 13230 13850
rect 13250 13790 13310 13850
rect 13330 13790 13390 13850
rect 13170 13710 13230 13770
rect 13250 13710 13310 13770
rect 13330 13710 13390 13770
rect 10930 13120 10990 13130
rect 10930 13080 10940 13120
rect 10940 13080 10980 13120
rect 10980 13080 10990 13120
rect 10930 13070 10990 13080
rect 10930 12990 10990 13050
rect 10930 12910 10990 12970
rect 11170 13120 11230 13130
rect 11170 13080 11180 13120
rect 11180 13080 11220 13120
rect 11220 13080 11230 13120
rect 11170 13070 11230 13080
rect 11170 12990 11230 13050
rect 11170 12910 11230 12970
rect 11410 13120 11470 13130
rect 11410 13080 11420 13120
rect 11420 13080 11460 13120
rect 11460 13080 11470 13120
rect 11410 13070 11470 13080
rect 11410 12990 11470 13050
rect 11410 12910 11470 12970
rect 11650 13120 11710 13130
rect 11650 13080 11660 13120
rect 11660 13080 11700 13120
rect 11700 13080 11710 13120
rect 11650 13070 11710 13080
rect 11650 12990 11710 13050
rect 11650 12910 11710 12970
rect 12290 13120 12350 13130
rect 12290 13080 12300 13120
rect 12300 13080 12340 13120
rect 12340 13080 12350 13120
rect 12290 13070 12350 13080
rect 12290 12990 12350 13050
rect 12290 12910 12350 12970
rect 12530 13120 12590 13130
rect 12530 13080 12540 13120
rect 12540 13080 12580 13120
rect 12580 13080 12590 13120
rect 12530 13070 12590 13080
rect 12530 12990 12590 13050
rect 12530 12910 12590 12970
rect 12770 13120 12830 13130
rect 12770 13080 12780 13120
rect 12780 13080 12820 13120
rect 12820 13080 12830 13120
rect 12770 13070 12830 13080
rect 12770 12990 12830 13050
rect 12770 12910 12830 12970
rect 10750 12800 10810 12860
rect 11500 12800 11560 12860
rect 11720 12800 11780 12860
rect 11980 12800 12040 12860
rect 12200 12800 12260 12860
rect 12460 12800 12520 12860
rect 11433 12742 11485 12750
rect 11433 12708 11443 12742
rect 11443 12708 11477 12742
rect 11477 12708 11485 12742
rect 11433 12698 11485 12708
rect 11793 12742 11845 12750
rect 11793 12708 11803 12742
rect 11803 12708 11837 12742
rect 11837 12708 11845 12742
rect 11793 12698 11845 12708
rect 11913 12742 11965 12750
rect 11913 12708 11923 12742
rect 11923 12708 11957 12742
rect 11957 12708 11965 12742
rect 11913 12698 11965 12708
rect 12273 12742 12325 12750
rect 12273 12708 12283 12742
rect 12283 12708 12317 12742
rect 12317 12708 12325 12742
rect 12273 12698 12325 12708
rect 12393 12742 12445 12750
rect 12393 12708 12403 12742
rect 12403 12708 12437 12742
rect 12437 12708 12445 12742
rect 12393 12698 12445 12708
rect 12810 12720 12870 12730
rect 12810 12680 12820 12720
rect 12820 12680 12860 12720
rect 12860 12680 12870 12720
rect 12810 12670 12870 12680
rect 12810 12640 12870 12650
rect 12810 12600 12820 12640
rect 12820 12600 12860 12640
rect 12860 12600 12870 12640
rect 12810 12590 12870 12600
rect 11536 12512 11588 12522
rect 11536 12478 11544 12512
rect 11544 12478 11578 12512
rect 11578 12478 11588 12512
rect 11536 12470 11588 12478
rect 11694 12512 11746 12522
rect 11694 12478 11702 12512
rect 11702 12478 11736 12512
rect 11736 12478 11746 12512
rect 11694 12470 11746 12478
rect 11610 12360 11670 12420
rect 11370 12250 11430 12310
rect 10630 11980 10690 12040
rect 10710 11980 10770 12040
rect 11130 11980 11190 12040
rect 11370 11980 11430 12040
rect 10890 11910 10950 11920
rect 10890 11870 10900 11910
rect 10900 11870 10940 11910
rect 10940 11870 10950 11910
rect 10890 11860 10950 11870
rect 10650 11520 10710 11580
rect 12018 12512 12070 12522
rect 12018 12478 12026 12512
rect 12026 12478 12060 12512
rect 12060 12478 12070 12512
rect 12018 12470 12070 12478
rect 12172 12512 12224 12522
rect 12172 12478 12180 12512
rect 12180 12478 12214 12512
rect 12214 12478 12224 12512
rect 12172 12470 12224 12478
rect 12090 12360 12150 12420
rect 12496 12512 12548 12522
rect 12496 12478 12504 12512
rect 12504 12478 12538 12512
rect 12538 12478 12548 12512
rect 12496 12470 12548 12478
rect 12810 12560 12870 12570
rect 12810 12520 12820 12560
rect 12820 12520 12860 12560
rect 12860 12520 12870 12560
rect 12810 12510 12870 12520
rect 12570 12360 12630 12420
rect 11850 12250 11910 12310
rect 12330 12250 12390 12310
rect 11850 11980 11910 12040
rect 12090 11980 12150 12040
rect 12570 11980 12630 12040
rect 12750 11980 12810 12040
rect 11610 11910 11670 11920
rect 11610 11870 11620 11910
rect 11620 11870 11660 11910
rect 11660 11870 11670 11910
rect 11610 11860 11670 11870
rect 11370 11520 11430 11580
rect 12330 11910 12390 11920
rect 12330 11870 12340 11910
rect 12340 11870 12380 11910
rect 12380 11870 12390 11910
rect 12330 11860 12390 11870
rect 12090 11520 12150 11580
rect 12810 11520 12870 11580
rect 14590 13870 14650 13930
rect 14590 13790 14650 13850
rect 14590 13760 14650 13770
rect 14590 13720 14600 13760
rect 14600 13720 14640 13760
rect 14640 13720 14650 13760
rect 14590 13710 14650 13720
rect 13170 12670 13230 12730
rect 13250 12670 13310 12730
rect 13330 12670 13390 12730
rect 13170 12590 13230 12650
rect 13250 12590 13310 12650
rect 13330 12590 13390 12650
rect 13170 12510 13230 12570
rect 13250 12510 13310 12570
rect 13330 12510 13390 12570
rect 13730 13120 13790 13130
rect 13730 13080 13740 13120
rect 13740 13080 13780 13120
rect 13780 13080 13790 13120
rect 13730 13070 13790 13080
rect 13730 12990 13790 13050
rect 13730 12910 13790 12970
rect 13970 13120 14030 13130
rect 13970 13080 13980 13120
rect 13980 13080 14020 13120
rect 14020 13080 14030 13120
rect 13970 13070 14030 13080
rect 13970 12990 14030 13050
rect 13970 12910 14030 12970
rect 14210 13120 14270 13130
rect 14210 13080 14220 13120
rect 14220 13080 14260 13120
rect 14260 13080 14270 13120
rect 14210 13070 14270 13080
rect 14210 12990 14270 13050
rect 14210 12910 14270 12970
rect 14850 13120 14910 13130
rect 14850 13080 14860 13120
rect 14860 13080 14900 13120
rect 14900 13080 14910 13120
rect 14850 13070 14910 13080
rect 14850 12990 14910 13050
rect 14850 12910 14910 12970
rect 15090 13120 15150 13130
rect 15090 13080 15100 13120
rect 15100 13080 15140 13120
rect 15140 13080 15150 13120
rect 15090 13070 15150 13080
rect 15090 12990 15150 13050
rect 15090 12910 15150 12970
rect 15330 13120 15390 13130
rect 15330 13080 15340 13120
rect 15340 13080 15380 13120
rect 15380 13080 15390 13120
rect 15330 13070 15390 13080
rect 15330 12990 15390 13050
rect 15330 12910 15390 12970
rect 15570 13120 15630 13130
rect 15570 13080 15580 13120
rect 15580 13080 15620 13120
rect 15620 13080 15630 13120
rect 15570 13070 15630 13080
rect 15570 12990 15630 13050
rect 15570 12910 15630 12970
rect 14040 12800 14100 12860
rect 14300 12800 14360 12860
rect 14520 12800 14580 12860
rect 14780 12800 14840 12860
rect 15000 12800 15060 12860
rect 15750 12800 15810 12860
rect 13690 12720 13750 12730
rect 13690 12680 13700 12720
rect 13700 12680 13740 12720
rect 13740 12680 13750 12720
rect 13690 12670 13750 12680
rect 14115 12742 14167 12750
rect 14115 12708 14123 12742
rect 14123 12708 14157 12742
rect 14157 12708 14167 12742
rect 14115 12698 14167 12708
rect 14235 12742 14287 12750
rect 14235 12708 14243 12742
rect 14243 12708 14277 12742
rect 14277 12708 14287 12742
rect 14235 12698 14287 12708
rect 14595 12742 14647 12750
rect 14595 12708 14603 12742
rect 14603 12708 14637 12742
rect 14637 12708 14647 12742
rect 14595 12698 14647 12708
rect 14715 12742 14767 12750
rect 14715 12708 14723 12742
rect 14723 12708 14757 12742
rect 14757 12708 14767 12742
rect 14715 12698 14767 12708
rect 15075 12742 15127 12750
rect 15075 12708 15083 12742
rect 15083 12708 15117 12742
rect 15117 12708 15127 12742
rect 15075 12698 15127 12708
rect 16160 12690 16220 12750
rect 13690 12640 13750 12650
rect 13690 12600 13700 12640
rect 13700 12600 13740 12640
rect 13740 12600 13750 12640
rect 13690 12590 13750 12600
rect 13690 12560 13750 12570
rect 13690 12520 13700 12560
rect 13700 12520 13740 12560
rect 13740 12520 13750 12560
rect 13690 12510 13750 12520
rect 14012 12512 14064 12522
rect 14012 12478 14022 12512
rect 14022 12478 14056 12512
rect 14056 12478 14064 12512
rect 14012 12470 14064 12478
rect 13930 12360 13990 12420
rect 14336 12512 14388 12522
rect 14336 12478 14346 12512
rect 14346 12478 14380 12512
rect 14380 12478 14388 12512
rect 14336 12470 14388 12478
rect 14490 12512 14542 12522
rect 14490 12478 14500 12512
rect 14500 12478 14534 12512
rect 14534 12478 14542 12512
rect 14490 12470 14542 12478
rect 14410 12360 14470 12420
rect 14814 12512 14866 12522
rect 14814 12478 14824 12512
rect 14824 12478 14858 12512
rect 14858 12478 14866 12512
rect 14814 12470 14866 12478
rect 14972 12512 15024 12522
rect 14972 12478 14982 12512
rect 14982 12478 15016 12512
rect 15016 12478 15024 12512
rect 14972 12470 15024 12478
rect 14890 12360 14950 12420
rect 14170 12250 14230 12310
rect 14650 12250 14710 12310
rect 13750 12140 13810 12200
rect 13750 12060 13810 12120
rect 13750 11980 13810 12040
rect 13930 12140 13990 12200
rect 13930 12060 13990 12120
rect 13930 11980 13990 12040
rect 14170 12140 14230 12200
rect 14170 12060 14230 12120
rect 14170 11980 14230 12040
rect 14410 12140 14470 12200
rect 14410 12060 14470 12120
rect 14410 11980 14470 12040
rect 14650 12140 14710 12200
rect 14650 12060 14710 12120
rect 14650 11980 14710 12040
rect 13070 11520 13130 11580
rect 13430 11520 13490 11580
rect 10530 11410 10590 11470
rect 10530 11330 10590 11390
rect 10530 11250 10590 11310
rect 10770 11410 10830 11470
rect 10770 11330 10830 11390
rect 10770 11250 10830 11310
rect 11010 11410 11070 11470
rect 11010 11330 11070 11390
rect 11010 11250 11070 11310
rect 11250 11410 11310 11470
rect 11250 11330 11310 11390
rect 11250 11250 11310 11310
rect 11490 11410 11550 11470
rect 11490 11330 11550 11390
rect 11490 11250 11550 11310
rect 11730 11410 11790 11470
rect 11730 11330 11790 11390
rect 11730 11250 11790 11310
rect 11970 11410 12030 11470
rect 11970 11330 12030 11390
rect 11970 11250 12030 11310
rect 12210 11410 12270 11470
rect 12210 11330 12270 11390
rect 12210 11250 12270 11310
rect 12450 11410 12510 11470
rect 12450 11330 12510 11390
rect 12450 11250 12510 11310
rect 12690 11410 12750 11470
rect 12690 11330 12750 11390
rect 12690 11250 12750 11310
rect 12930 11410 12990 11470
rect 12930 11330 12990 11390
rect 12930 11250 12990 11310
rect 11810 11140 11870 11200
rect 13250 11140 13310 11200
rect 12170 11030 12230 11090
rect 11900 10750 11960 10760
rect 11900 10710 11910 10750
rect 11910 10710 11950 10750
rect 11950 10710 11960 10750
rect 11900 10700 11960 10710
rect 12080 10750 12140 10760
rect 12080 10710 12090 10750
rect 12090 10710 12130 10750
rect 12130 10710 12140 10750
rect 12080 10700 12140 10710
rect 12530 10920 12590 10980
rect 12260 10750 12320 10760
rect 12260 10710 12270 10750
rect 12270 10710 12310 10750
rect 12310 10710 12320 10750
rect 12260 10700 12320 10710
rect 12440 10750 12500 10760
rect 12440 10710 12450 10750
rect 12450 10710 12490 10750
rect 12490 10710 12500 10750
rect 12440 10700 12500 10710
rect 12890 10810 12950 10870
rect 12620 10750 12680 10760
rect 12620 10710 12630 10750
rect 12630 10710 12670 10750
rect 12670 10710 12680 10750
rect 12620 10700 12680 10710
rect 12800 10750 12860 10760
rect 12800 10710 12810 10750
rect 12810 10710 12850 10750
rect 12850 10710 12860 10750
rect 12800 10700 12860 10710
rect 12980 10750 13040 10760
rect 12980 10710 12990 10750
rect 12990 10710 13030 10750
rect 13030 10710 13040 10750
rect 12980 10700 13040 10710
rect 13160 10750 13220 10760
rect 13160 10710 13170 10750
rect 13170 10710 13210 10750
rect 13210 10710 13220 10750
rect 13160 10700 13220 10710
rect 13690 11520 13750 11580
rect 14170 11910 14230 11920
rect 14170 11870 14180 11910
rect 14180 11870 14220 11910
rect 14220 11870 14230 11910
rect 14170 11860 14230 11870
rect 14410 11520 14470 11580
rect 15130 12250 15190 12310
rect 15130 12140 15190 12200
rect 15130 12060 15190 12120
rect 15130 11980 15190 12040
rect 15370 12140 15430 12200
rect 15370 12060 15430 12120
rect 15370 11980 15430 12040
rect 15790 12140 15850 12200
rect 15790 12060 15850 12120
rect 15790 11980 15850 12040
rect 14890 11910 14950 11920
rect 14890 11870 14900 11910
rect 14900 11870 14940 11910
rect 14940 11870 14950 11910
rect 14890 11860 14950 11870
rect 15130 11520 15190 11580
rect 15610 11910 15670 11920
rect 15610 11870 15620 11910
rect 15620 11870 15660 11910
rect 15660 11870 15670 11910
rect 15610 11860 15670 11870
rect 15850 11520 15910 11580
rect 13570 11410 13630 11470
rect 13570 11330 13630 11390
rect 13570 11250 13630 11310
rect 13810 11410 13870 11470
rect 13810 11330 13870 11390
rect 13810 11250 13870 11310
rect 14050 11410 14110 11470
rect 14050 11330 14110 11390
rect 14050 11250 14110 11310
rect 14290 11410 14350 11470
rect 14290 11330 14350 11390
rect 14290 11250 14350 11310
rect 14530 11410 14590 11470
rect 14530 11330 14590 11390
rect 14530 11250 14590 11310
rect 14770 11410 14830 11470
rect 14770 11330 14830 11390
rect 14770 11250 14830 11310
rect 15010 11410 15070 11470
rect 15010 11330 15070 11390
rect 15010 11250 15070 11310
rect 15250 11410 15310 11470
rect 15250 11330 15310 11390
rect 15250 11250 15310 11310
rect 15490 11410 15550 11470
rect 15490 11330 15550 11390
rect 15490 11250 15550 11310
rect 15730 11410 15790 11470
rect 15730 11330 15790 11390
rect 15730 11250 15790 11310
rect 14690 11140 14750 11200
rect 14330 11030 14390 11090
rect 13970 10920 14030 10980
rect 13610 10810 13670 10870
rect 13340 10750 13400 10760
rect 13340 10710 13350 10750
rect 13350 10710 13390 10750
rect 13390 10710 13400 10750
rect 13340 10700 13400 10710
rect 13430 10700 13490 10760
rect 13520 10750 13580 10760
rect 13520 10710 13530 10750
rect 13530 10710 13570 10750
rect 13570 10710 13580 10750
rect 13520 10700 13580 10710
rect 13700 10750 13760 10760
rect 13700 10710 13710 10750
rect 13710 10710 13750 10750
rect 13750 10710 13760 10750
rect 13700 10700 13760 10710
rect 13880 10750 13940 10760
rect 13880 10710 13890 10750
rect 13890 10710 13930 10750
rect 13930 10710 13940 10750
rect 13880 10700 13940 10710
rect 14060 10750 14120 10760
rect 14060 10710 14070 10750
rect 14070 10710 14110 10750
rect 14110 10710 14120 10750
rect 14060 10700 14120 10710
rect 14240 10750 14300 10760
rect 14240 10710 14250 10750
rect 14250 10710 14290 10750
rect 14290 10710 14300 10750
rect 14240 10700 14300 10710
rect 14420 10750 14480 10760
rect 14420 10710 14430 10750
rect 14430 10710 14470 10750
rect 14470 10710 14480 10750
rect 14420 10700 14480 10710
rect 14600 10750 14660 10760
rect 14600 10710 14610 10750
rect 14610 10710 14650 10750
rect 14650 10710 14660 10750
rect 14600 10700 14660 10710
rect 15720 11030 15780 11090
rect 15250 10920 15310 10980
rect 15600 10550 15660 10560
rect 15600 10510 15610 10550
rect 15610 10510 15650 10550
rect 15650 10510 15660 10550
rect 15600 10500 15660 10510
rect 15970 11410 16030 11470
rect 15970 11330 16030 11390
rect 15970 11250 16030 11310
rect 16250 12460 16310 12520
rect 16790 14430 16850 14490
rect 17580 16690 17640 16750
rect 16360 12140 16420 12200
rect 16440 12140 16500 12200
rect 16520 12140 16580 12200
rect 16360 12060 16420 12120
rect 16440 12060 16500 12120
rect 16520 12060 16580 12120
rect 16360 11980 16420 12040
rect 16440 11980 16500 12040
rect 16520 11980 16580 12040
rect 17960 15990 18020 16050
rect 18130 17390 18190 17450
rect 18800 16690 18860 16750
rect 18800 15290 18860 15350
rect 18660 14320 18720 14380
rect 17580 11520 17640 11580
rect 16250 10920 16310 10980
rect 16160 10810 16220 10870
rect 15840 10550 15900 10560
rect 15840 10510 15850 10550
rect 15850 10510 15890 10550
rect 15890 10510 15900 10550
rect 15840 10500 15900 10510
rect 15250 10160 15310 10220
rect 15720 10210 15780 10220
rect 15720 10170 15730 10210
rect 15730 10170 15770 10210
rect 15770 10170 15780 10210
rect 15720 10160 15780 10170
rect 11630 10010 11690 10020
rect 11630 9970 11640 10010
rect 11640 9970 11680 10010
rect 11680 9970 11690 10010
rect 11630 9960 11690 9970
rect 11630 9880 11690 9940
rect 11630 9800 11690 9860
rect 11990 10010 12050 10020
rect 11990 9970 12000 10010
rect 12000 9970 12040 10010
rect 12040 9970 12050 10010
rect 11990 9960 12050 9970
rect 11990 9880 12050 9940
rect 11990 9800 12050 9860
rect 12350 10010 12410 10020
rect 12350 9970 12360 10010
rect 12360 9970 12400 10010
rect 12400 9970 12410 10010
rect 12350 9960 12410 9970
rect 12350 9880 12410 9940
rect 12350 9800 12410 9860
rect 12710 10010 12770 10020
rect 12710 9970 12720 10010
rect 12720 9970 12760 10010
rect 12760 9970 12770 10010
rect 12710 9960 12770 9970
rect 12710 9880 12770 9940
rect 12710 9800 12770 9860
rect 13070 10010 13130 10020
rect 13070 9970 13080 10010
rect 13080 9970 13120 10010
rect 13120 9970 13130 10010
rect 13070 9960 13130 9970
rect 13070 9880 13130 9940
rect 13070 9800 13130 9860
rect 13430 10010 13490 10020
rect 13430 9970 13440 10010
rect 13440 9970 13480 10010
rect 13480 9970 13490 10010
rect 13430 9960 13490 9970
rect 13430 9880 13490 9940
rect 13430 9800 13490 9860
rect 13790 10010 13850 10020
rect 13790 9970 13800 10010
rect 13800 9970 13840 10010
rect 13840 9970 13850 10010
rect 13790 9960 13850 9970
rect 13790 9880 13850 9940
rect 13790 9800 13850 9860
rect 14150 10010 14210 10020
rect 14150 9970 14160 10010
rect 14160 9970 14200 10010
rect 14200 9970 14210 10010
rect 14150 9960 14210 9970
rect 14150 9880 14210 9940
rect 14150 9800 14210 9860
rect 14510 10010 14570 10020
rect 14510 9970 14520 10010
rect 14520 9970 14560 10010
rect 14560 9970 14570 10010
rect 14510 9960 14570 9970
rect 14510 9880 14570 9940
rect 14510 9800 14570 9860
rect 14870 10010 14930 10020
rect 14870 9970 14880 10010
rect 14880 9970 14920 10010
rect 14920 9970 14930 10010
rect 14870 9960 14930 9970
rect 14870 9880 14930 9940
rect 14870 9800 14930 9860
rect 15500 9960 15560 10020
rect 15500 9880 15560 9940
rect 15500 9800 15560 9860
rect 15940 9960 16000 10020
rect 15940 9880 16000 9940
rect 15940 9800 16000 9860
rect 11808 9742 11860 9750
rect 11808 9708 11818 9742
rect 11818 9708 11852 9742
rect 11852 9708 11860 9742
rect 11808 9698 11860 9708
rect 11918 9742 11970 9750
rect 11918 9708 11928 9742
rect 11928 9708 11962 9742
rect 11962 9708 11970 9742
rect 11918 9698 11970 9708
rect 12028 9742 12080 9750
rect 12028 9708 12038 9742
rect 12038 9708 12072 9742
rect 12072 9708 12080 9742
rect 12028 9698 12080 9708
rect 12138 9742 12190 9750
rect 12138 9708 12148 9742
rect 12148 9708 12182 9742
rect 12182 9708 12190 9742
rect 12138 9698 12190 9708
rect 12248 9742 12300 9750
rect 12248 9708 12258 9742
rect 12258 9708 12292 9742
rect 12292 9708 12300 9742
rect 12248 9698 12300 9708
rect 12358 9742 12410 9750
rect 12358 9708 12368 9742
rect 12368 9708 12402 9742
rect 12402 9708 12410 9742
rect 12358 9698 12410 9708
rect 12468 9742 12520 9750
rect 12468 9708 12478 9742
rect 12478 9708 12512 9742
rect 12512 9708 12520 9742
rect 12468 9698 12520 9708
rect 12578 9742 12630 9750
rect 12578 9708 12588 9742
rect 12588 9708 12622 9742
rect 12622 9708 12630 9742
rect 12578 9698 12630 9708
rect 12688 9742 12740 9750
rect 12688 9708 12698 9742
rect 12698 9708 12732 9742
rect 12732 9708 12740 9742
rect 12688 9698 12740 9708
rect 12798 9742 12850 9750
rect 12798 9708 12808 9742
rect 12808 9708 12842 9742
rect 12842 9708 12850 9742
rect 12798 9698 12850 9708
rect 13708 9742 13760 9750
rect 13708 9708 13718 9742
rect 13718 9708 13752 9742
rect 13752 9708 13760 9742
rect 13708 9698 13760 9708
rect 13818 9742 13870 9750
rect 13818 9708 13828 9742
rect 13828 9708 13862 9742
rect 13862 9708 13870 9742
rect 13818 9698 13870 9708
rect 13928 9742 13980 9750
rect 13928 9708 13938 9742
rect 13938 9708 13972 9742
rect 13972 9708 13980 9742
rect 13928 9698 13980 9708
rect 14038 9742 14090 9750
rect 14038 9708 14048 9742
rect 14048 9708 14082 9742
rect 14082 9708 14090 9742
rect 14038 9698 14090 9708
rect 14148 9742 14200 9750
rect 14148 9708 14158 9742
rect 14158 9708 14192 9742
rect 14192 9708 14200 9742
rect 14148 9698 14200 9708
rect 14258 9742 14310 9750
rect 14258 9708 14268 9742
rect 14268 9708 14302 9742
rect 14302 9708 14310 9742
rect 14258 9698 14310 9708
rect 14368 9742 14420 9750
rect 14368 9708 14378 9742
rect 14378 9708 14412 9742
rect 14412 9708 14420 9742
rect 14368 9698 14420 9708
rect 14478 9742 14530 9750
rect 14478 9708 14488 9742
rect 14488 9708 14522 9742
rect 14522 9708 14530 9742
rect 14478 9698 14530 9708
rect 14588 9742 14640 9750
rect 14588 9708 14598 9742
rect 14598 9708 14632 9742
rect 14632 9708 14640 9742
rect 14588 9698 14640 9708
rect 14698 9742 14750 9750
rect 14698 9708 14708 9742
rect 14708 9708 14742 9742
rect 14742 9708 14750 9742
rect 14698 9698 14750 9708
rect 11640 9410 11700 9420
rect 11640 9370 11650 9410
rect 11650 9370 11690 9410
rect 11690 9370 11700 9410
rect 11640 9360 11700 9370
rect 11860 9360 11920 9420
rect 12080 9360 12140 9420
rect 12300 9360 12360 9420
rect 12520 9360 12580 9420
rect 12740 9360 12800 9420
rect 12960 9410 13020 9420
rect 12960 9370 12970 9410
rect 12970 9370 13010 9410
rect 13010 9370 13020 9410
rect 12960 9360 13020 9370
rect 13540 9410 13600 9420
rect 13540 9370 13550 9410
rect 13550 9370 13590 9410
rect 13590 9370 13600 9410
rect 13540 9360 13600 9370
rect 9690 9250 9750 9310
rect 11750 9250 11810 9310
rect 11970 9250 12030 9310
rect 12190 9250 12250 9310
rect 12410 9250 12470 9310
rect 12630 9250 12690 9310
rect 13760 9360 13820 9420
rect 13980 9360 14040 9420
rect 14200 9360 14260 9420
rect 14420 9360 14480 9420
rect 14640 9360 14700 9420
rect 14860 9410 14920 9420
rect 14860 9370 14870 9410
rect 14870 9370 14910 9410
rect 14910 9370 14920 9410
rect 14860 9360 14920 9370
rect 12850 9250 12910 9310
rect 13650 9240 13710 9300
rect 13650 9160 13710 9220
rect 13650 9080 13710 9140
rect 13870 9240 13930 9300
rect 13870 9160 13930 9220
rect 13870 9080 13930 9140
rect 14090 9240 14150 9300
rect 14090 9160 14150 9220
rect 14090 9080 14150 9140
rect 14310 9240 14370 9300
rect 14310 9160 14370 9220
rect 14310 9080 14370 9140
rect 14530 9240 14590 9300
rect 14530 9160 14590 9220
rect 14530 9080 14590 9140
rect 14750 9240 14810 9300
rect 14750 9160 14810 9220
rect 14750 9080 14810 9140
<< metal2 >>
rect 8870 19190 18270 19200
rect 8870 19130 8880 19190
rect 8940 19130 18200 19190
rect 18260 19130 18270 19190
rect 8870 19120 18270 19130
rect 8450 19080 17650 19090
rect 8450 19020 8460 19080
rect 8520 19020 9250 19080
rect 9310 19020 10690 19080
rect 10750 19020 13250 19080
rect 13310 19020 15680 19080
rect 15740 19020 16790 19080
rect 16850 19020 17580 19080
rect 17640 19020 17650 19080
rect 8450 19000 17650 19020
rect 8450 18940 8460 19000
rect 8520 18940 9250 19000
rect 9310 18940 10690 19000
rect 10750 18940 13250 19000
rect 13310 18940 15680 19000
rect 15740 18940 16790 19000
rect 16850 18940 17580 19000
rect 17640 18940 17650 19000
rect 8450 18920 17650 18940
rect 8450 18860 8460 18920
rect 8520 18860 9250 18920
rect 9310 18860 10690 18920
rect 10750 18860 13250 18920
rect 13310 18860 15680 18920
rect 15740 18860 16790 18920
rect 16850 18860 17580 18920
rect 17640 18860 17650 18920
rect 8450 18850 17650 18860
rect 18190 18850 18270 18860
rect 18190 18790 18200 18850
rect 18260 18790 18270 18850
rect 18190 18780 18270 18790
rect 8450 18450 8950 18460
rect 8450 18440 8880 18450
rect 8450 18040 8460 18440
rect 8520 18390 8880 18440
rect 8940 18390 8950 18450
rect 8520 18370 8950 18390
rect 8520 18310 8880 18370
rect 8940 18310 8950 18370
rect 8520 18280 8950 18310
rect 8520 18220 8880 18280
rect 8940 18220 8950 18280
rect 8520 18190 8950 18220
rect 8520 18130 8880 18190
rect 8940 18130 8950 18190
rect 8520 18110 8950 18130
rect 8520 18050 8880 18110
rect 8940 18050 8950 18110
rect 8520 18040 8950 18050
rect 8450 18030 8950 18040
rect 17570 18450 18030 18460
rect 17570 18440 17960 18450
rect 17570 18040 17580 18440
rect 17640 18390 17960 18440
rect 18020 18390 18030 18450
rect 17640 18370 18030 18390
rect 17640 18310 17960 18370
rect 18020 18310 18030 18370
rect 17640 18280 18030 18310
rect 17640 18220 17960 18280
rect 18020 18220 18030 18280
rect 17640 18190 18030 18220
rect 17640 18130 17960 18190
rect 18020 18130 18030 18190
rect 17640 18110 18030 18130
rect 17640 18050 17960 18110
rect 18020 18050 18030 18110
rect 18640 18150 18740 18170
rect 18640 18090 18660 18150
rect 18720 18090 18740 18150
rect 18640 18070 18740 18090
rect 17640 18040 18030 18050
rect 17570 18030 18030 18040
rect 18120 17450 18200 17460
rect 18120 17390 18130 17450
rect 18190 17390 18200 17450
rect 18120 17380 18200 17390
rect 11140 16810 11650 16820
rect 11140 16750 11150 16810
rect 11210 16750 11580 16810
rect 11640 16750 11650 16810
rect 11140 16740 11650 16750
rect 13240 16810 15420 16820
rect 13240 16750 13250 16810
rect 13310 16750 15350 16810
rect 15410 16750 15420 16810
rect 13240 16740 15420 16750
rect 17570 16750 18880 16770
rect 17570 16690 17580 16750
rect 17640 16690 18800 16750
rect 18860 16690 18880 16750
rect 17570 16670 18880 16690
rect 17950 16050 19070 16060
rect 17950 15990 17960 16050
rect 18020 15990 19000 16050
rect 19060 15990 19070 16050
rect 17950 15980 19070 15990
rect 16350 15350 18880 15370
rect 16350 15290 16360 15350
rect 16420 15290 16440 15350
rect 16500 15290 16520 15350
rect 16580 15290 18800 15350
rect 18860 15290 18880 15350
rect 16350 15270 18880 15290
rect 15340 14800 16320 14810
rect 15340 14740 15350 14800
rect 15410 14740 16010 14800
rect 16070 14740 16250 14800
rect 16310 14740 16320 14800
rect 15340 14730 16320 14740
rect 10350 14720 14030 14730
rect 10350 14660 10360 14720
rect 10420 14660 13960 14720
rect 14020 14660 14030 14720
rect 10350 14650 14030 14660
rect 11140 14610 12550 14620
rect 11140 14550 11150 14610
rect 11210 14550 12552 14610
rect 11140 14540 12552 14550
rect 12622 14540 12632 14610
rect 13940 14540 13950 14610
rect 14020 14590 14030 14610
rect 16150 14600 16230 14610
rect 16150 14590 16160 14600
rect 14020 14550 16160 14590
rect 14020 14540 14030 14550
rect 16150 14540 16160 14550
rect 16220 14540 16230 14600
rect 16150 14530 16230 14540
rect 9680 14490 16860 14500
rect 9680 14430 9690 14490
rect 9750 14430 16790 14490
rect 16850 14430 16860 14490
rect 9680 14420 16860 14430
rect 10620 14380 18730 14390
rect 10620 14320 10630 14380
rect 10690 14320 11040 14380
rect 11100 14320 18660 14380
rect 18720 14320 18730 14380
rect 10620 14310 18730 14320
rect 15470 14250 15550 14260
rect 9460 14210 11160 14220
rect 9460 14150 9470 14210
rect 9530 14150 11090 14210
rect 11150 14150 11160 14210
rect 9460 14140 11160 14150
rect 15470 14190 15480 14250
rect 15540 14190 15550 14250
rect 15470 14170 15550 14190
rect 15470 14110 15480 14170
rect 15540 14110 15550 14170
rect 15470 14100 15550 14110
rect 11160 14040 11240 14050
rect 11160 13980 11170 14040
rect 11230 14030 11240 14040
rect 11320 14040 11400 14050
rect 11320 14030 11330 14040
rect 11230 13990 11330 14030
rect 11230 13980 11240 13990
rect 11160 13970 11240 13980
rect 11320 13980 11330 13990
rect 11390 14030 11400 14040
rect 11480 14040 11560 14050
rect 11480 14030 11490 14040
rect 11390 13990 11490 14030
rect 11390 13980 11400 13990
rect 11320 13970 11400 13980
rect 11480 13980 11490 13990
rect 11550 14030 11560 14040
rect 11640 14040 11720 14050
rect 11640 14030 11650 14040
rect 11550 13990 11650 14030
rect 11550 13980 11560 13990
rect 11480 13970 11560 13980
rect 11640 13980 11650 13990
rect 11710 14030 11720 14040
rect 11800 14040 11880 14050
rect 11800 14030 11810 14040
rect 11710 13990 11810 14030
rect 11710 13980 11720 13990
rect 11640 13970 11720 13980
rect 11800 13980 11810 13990
rect 11870 14030 11880 14040
rect 11960 14040 12040 14050
rect 11960 14030 11970 14040
rect 11870 13990 11970 14030
rect 11870 13980 11880 13990
rect 11800 13970 11880 13980
rect 11960 13980 11970 13990
rect 12030 14030 12040 14040
rect 12120 14040 12200 14050
rect 12120 14030 12130 14040
rect 12030 13990 12130 14030
rect 12030 13980 12040 13990
rect 11960 13970 12040 13980
rect 12120 13980 12130 13990
rect 12190 14030 12200 14040
rect 12280 14040 12360 14050
rect 12280 14030 12290 14040
rect 12190 13990 12290 14030
rect 12190 13980 12200 13990
rect 12120 13970 12200 13980
rect 12280 13980 12290 13990
rect 12350 14030 12360 14040
rect 12440 14040 12520 14050
rect 12440 14030 12450 14040
rect 12350 13990 12450 14030
rect 12350 13980 12360 13990
rect 12280 13970 12360 13980
rect 12440 13980 12450 13990
rect 12510 14030 12520 14040
rect 12600 14040 12680 14050
rect 12600 14030 12610 14040
rect 12510 13990 12610 14030
rect 12510 13980 12520 13990
rect 12440 13970 12520 13980
rect 12600 13980 12610 13990
rect 12670 14030 12680 14040
rect 12760 14040 12840 14050
rect 12760 14030 12770 14040
rect 12670 13990 12770 14030
rect 12670 13980 12680 13990
rect 12600 13970 12680 13980
rect 12760 13980 12770 13990
rect 12830 14030 12840 14040
rect 12920 14040 13000 14050
rect 12920 14030 12930 14040
rect 12830 13990 12930 14030
rect 12830 13980 12840 13990
rect 12760 13970 12840 13980
rect 12920 13980 12930 13990
rect 12990 14030 13000 14040
rect 13080 14040 13160 14050
rect 13080 14030 13090 14040
rect 12990 13990 13090 14030
rect 12990 13980 13000 13990
rect 12920 13970 13000 13980
rect 13080 13980 13090 13990
rect 13150 13980 13160 14040
rect 13080 13970 13160 13980
rect 13240 14040 13320 14050
rect 13240 13980 13250 14040
rect 13310 14030 13320 14040
rect 13400 14040 13480 14050
rect 13400 14030 13410 14040
rect 13310 13990 13410 14030
rect 13310 13980 13320 13990
rect 13240 13970 13320 13980
rect 13400 13980 13410 13990
rect 13470 14030 13480 14040
rect 13560 14040 13640 14050
rect 13560 14030 13570 14040
rect 13470 13990 13570 14030
rect 13470 13980 13480 13990
rect 13400 13970 13480 13980
rect 13560 13980 13570 13990
rect 13630 14030 13640 14040
rect 13720 14040 13800 14050
rect 13720 14030 13730 14040
rect 13630 13990 13730 14030
rect 13630 13980 13640 13990
rect 13560 13970 13640 13980
rect 13720 13980 13730 13990
rect 13790 14030 13800 14040
rect 13880 14040 13960 14050
rect 13880 14030 13890 14040
rect 13790 13990 13890 14030
rect 13790 13980 13800 13990
rect 13720 13970 13800 13980
rect 13880 13980 13890 13990
rect 13950 14030 13960 14040
rect 14040 14040 14120 14050
rect 14040 14030 14050 14040
rect 13950 13990 14050 14030
rect 13950 13980 13960 13990
rect 13880 13970 13960 13980
rect 14040 13980 14050 13990
rect 14110 14030 14120 14040
rect 14200 14040 14280 14050
rect 14200 14030 14210 14040
rect 14110 13990 14210 14030
rect 14110 13980 14120 13990
rect 14040 13970 14120 13980
rect 14200 13980 14210 13990
rect 14270 14030 14280 14040
rect 14360 14040 14440 14050
rect 14360 14030 14370 14040
rect 14270 13990 14370 14030
rect 14270 13980 14280 13990
rect 14200 13970 14280 13980
rect 14360 13980 14370 13990
rect 14430 14030 14440 14040
rect 14520 14040 14600 14050
rect 14520 14030 14530 14040
rect 14430 13990 14530 14030
rect 14430 13980 14440 13990
rect 14360 13970 14440 13980
rect 14520 13980 14530 13990
rect 14590 14030 14600 14040
rect 14680 14040 14760 14050
rect 14680 14030 14690 14040
rect 14590 13990 14690 14030
rect 14590 13980 14600 13990
rect 14520 13970 14600 13980
rect 14680 13980 14690 13990
rect 14750 14030 14760 14040
rect 14840 14040 14920 14050
rect 14840 14030 14850 14040
rect 14750 13990 14850 14030
rect 14750 13980 14760 13990
rect 14680 13970 14760 13980
rect 14840 13980 14850 13990
rect 14910 14030 14920 14040
rect 15000 14040 15080 14050
rect 15000 14030 15010 14040
rect 14910 13990 15010 14030
rect 14910 13980 14920 13990
rect 14840 13970 14920 13980
rect 15000 13980 15010 13990
rect 15070 14030 15080 14040
rect 15160 14040 15240 14050
rect 15160 14030 15170 14040
rect 15070 13990 15170 14030
rect 15070 13980 15080 13990
rect 15000 13970 15080 13980
rect 15160 13980 15170 13990
rect 15230 13980 15240 14040
rect 15160 13970 15240 13980
rect 11900 13930 14660 13940
rect 11900 13870 11910 13930
rect 11970 13870 13170 13930
rect 13230 13870 13250 13930
rect 13310 13870 13330 13930
rect 13390 13870 14590 13930
rect 14650 13870 14660 13930
rect 11900 13850 14660 13870
rect 11900 13790 11910 13850
rect 11970 13790 13170 13850
rect 13230 13790 13250 13850
rect 13310 13790 13330 13850
rect 13390 13790 14590 13850
rect 14650 13790 14660 13850
rect 11900 13770 14660 13790
rect 11900 13710 11910 13770
rect 11970 13710 13170 13770
rect 13230 13710 13250 13770
rect 13310 13710 13330 13770
rect 13390 13710 14590 13770
rect 14650 13710 14660 13770
rect 11900 13700 14660 13710
rect 10920 13130 15640 13140
rect 10920 13070 10930 13130
rect 10990 13070 11170 13130
rect 11230 13070 11410 13130
rect 11470 13070 11650 13130
rect 11710 13070 12290 13130
rect 12350 13070 12530 13130
rect 12590 13070 12770 13130
rect 12830 13070 13730 13130
rect 13790 13070 13970 13130
rect 14030 13070 14210 13130
rect 14270 13070 14850 13130
rect 14910 13070 15090 13130
rect 15150 13070 15330 13130
rect 15390 13070 15570 13130
rect 15630 13070 15640 13130
rect 10920 13050 15640 13070
rect 10920 12990 10930 13050
rect 10990 12990 11170 13050
rect 11230 12990 11410 13050
rect 11470 12990 11650 13050
rect 11710 12990 12290 13050
rect 12350 12990 12530 13050
rect 12590 12990 12770 13050
rect 12830 12990 13730 13050
rect 13790 12990 13970 13050
rect 14030 12990 14210 13050
rect 14270 12990 14850 13050
rect 14910 12990 15090 13050
rect 15150 12990 15330 13050
rect 15390 12990 15570 13050
rect 15630 12990 15640 13050
rect 10920 12970 15640 12990
rect 10920 12910 10930 12970
rect 10990 12910 11170 12970
rect 11230 12910 11410 12970
rect 11470 12910 11650 12970
rect 11710 12910 12290 12970
rect 12350 12910 12530 12970
rect 12590 12910 12770 12970
rect 12830 12910 13730 12970
rect 13790 12910 13970 12970
rect 14030 12910 14210 12970
rect 14270 12910 14850 12970
rect 14910 12910 15090 12970
rect 15150 12910 15330 12970
rect 15390 12910 15570 12970
rect 15630 12910 15640 12970
rect 10920 12900 15640 12910
rect 10740 12860 12530 12870
rect 10740 12800 10750 12860
rect 10810 12800 11500 12860
rect 11560 12800 11720 12860
rect 11780 12800 11980 12860
rect 12040 12800 12200 12860
rect 12260 12800 12460 12860
rect 12520 12800 12530 12860
rect 10740 12790 12530 12800
rect 14030 12860 15820 12870
rect 14030 12800 14040 12860
rect 14100 12800 14300 12860
rect 14360 12800 14520 12860
rect 14580 12800 14780 12860
rect 14840 12800 15000 12860
rect 15060 12800 15750 12860
rect 15810 12800 15820 12860
rect 14030 12790 15820 12800
rect 9680 12750 12449 12760
rect 9680 12690 9690 12750
rect 9750 12698 11433 12750
rect 11485 12698 11793 12750
rect 11845 12698 11913 12750
rect 11965 12698 12273 12750
rect 12325 12698 12393 12750
rect 12445 12698 12449 12750
rect 14111 12750 16230 12760
rect 9750 12690 12449 12698
rect 12800 12730 13760 12740
rect 9680 12680 9760 12690
rect 12800 12670 12810 12730
rect 12870 12670 13170 12730
rect 13230 12670 13250 12730
rect 13310 12670 13330 12730
rect 13390 12670 13690 12730
rect 13750 12670 13760 12730
rect 14111 12698 14115 12750
rect 14167 12698 14235 12750
rect 14287 12698 14595 12750
rect 14647 12698 14715 12750
rect 14767 12698 15075 12750
rect 15127 12698 16160 12750
rect 14111 12690 16160 12698
rect 16220 12690 16230 12750
rect 16150 12680 16230 12690
rect 12800 12650 13760 12670
rect 12800 12590 12810 12650
rect 12870 12590 13170 12650
rect 13230 12590 13250 12650
rect 13310 12590 13330 12650
rect 13390 12590 13690 12650
rect 13750 12590 13760 12650
rect 12800 12570 13760 12590
rect 9570 12522 12550 12530
rect 9570 12520 11536 12522
rect 9570 12460 9580 12520
rect 9640 12470 11536 12520
rect 11588 12470 11694 12522
rect 11746 12470 12018 12522
rect 12070 12470 12172 12522
rect 12224 12470 12496 12522
rect 12548 12470 12550 12522
rect 12800 12510 12810 12570
rect 12870 12510 13170 12570
rect 13230 12510 13250 12570
rect 13310 12510 13330 12570
rect 13390 12510 13690 12570
rect 13750 12510 13760 12570
rect 12800 12500 13760 12510
rect 14010 12522 16320 12530
rect 9640 12460 12550 12470
rect 14010 12470 14012 12522
rect 14064 12470 14336 12522
rect 14388 12470 14490 12522
rect 14542 12470 14814 12522
rect 14866 12470 14972 12522
rect 15024 12520 16320 12522
rect 15024 12470 16250 12520
rect 14010 12460 16250 12470
rect 16310 12460 16320 12520
rect 9570 12450 9650 12460
rect 16240 12450 16320 12460
rect 11600 12420 12640 12430
rect 11600 12360 11610 12420
rect 11670 12360 12090 12420
rect 12150 12360 12570 12420
rect 12630 12360 12640 12420
rect 11600 12350 12640 12360
rect 13920 12420 14960 12430
rect 13920 12360 13930 12420
rect 13990 12360 14410 12420
rect 14470 12360 14890 12420
rect 14950 12360 14960 12420
rect 13920 12350 14960 12360
rect 11360 12310 12400 12320
rect 11360 12250 11370 12310
rect 11430 12250 11850 12310
rect 11910 12250 12330 12310
rect 12390 12250 12400 12310
rect 11360 12240 12400 12250
rect 14160 12310 15200 12320
rect 14160 12250 14170 12310
rect 14230 12250 14650 12310
rect 14710 12250 15130 12310
rect 15190 12250 15200 12310
rect 14160 12240 15200 12250
rect 13740 12200 16590 12210
rect 13740 12140 13750 12200
rect 13810 12140 13930 12200
rect 13990 12140 14170 12200
rect 14230 12140 14410 12200
rect 14470 12140 14650 12200
rect 14710 12140 15130 12200
rect 15190 12140 15370 12200
rect 15430 12140 15790 12200
rect 15850 12140 16360 12200
rect 16420 12140 16440 12200
rect 16500 12140 16520 12200
rect 16580 12140 16590 12200
rect 13740 12120 16590 12140
rect 13740 12060 13750 12120
rect 13810 12060 13930 12120
rect 13990 12060 14170 12120
rect 14230 12060 14410 12120
rect 14470 12060 14650 12120
rect 14710 12060 15130 12120
rect 15190 12060 15370 12120
rect 15430 12060 15790 12120
rect 15850 12060 16360 12120
rect 16420 12060 16440 12120
rect 16500 12060 16520 12120
rect 16580 12060 16590 12120
rect 10620 12040 12820 12050
rect 10620 11980 10630 12040
rect 10690 11980 10710 12040
rect 10770 11980 11130 12040
rect 11190 11980 11370 12040
rect 11430 11980 11850 12040
rect 11910 11980 12090 12040
rect 12150 11980 12570 12040
rect 12630 11980 12750 12040
rect 12810 11980 12820 12040
rect 10620 11970 12820 11980
rect 13740 12040 16590 12060
rect 13740 11980 13750 12040
rect 13810 11980 13930 12040
rect 13990 11980 14170 12040
rect 14230 11980 14410 12040
rect 14470 11980 14650 12040
rect 14710 11980 15130 12040
rect 15190 11980 15370 12040
rect 15430 11980 15790 12040
rect 15850 11980 16360 12040
rect 16420 11980 16440 12040
rect 16500 11980 16520 12040
rect 16580 11980 16590 12040
rect 13740 11970 16590 11980
rect 10880 11920 10960 11930
rect 10880 11860 10890 11920
rect 10950 11910 10960 11920
rect 11600 11920 11680 11930
rect 11600 11910 11610 11920
rect 10950 11870 11610 11910
rect 10950 11860 10960 11870
rect 10880 11850 10960 11860
rect 11600 11860 11610 11870
rect 11670 11910 11680 11920
rect 12320 11920 12400 11930
rect 12320 11910 12330 11920
rect 11670 11870 12330 11910
rect 11670 11860 11680 11870
rect 11600 11850 11680 11860
rect 12320 11860 12330 11870
rect 12390 11860 12400 11920
rect 12320 11850 12400 11860
rect 14160 11920 14240 11930
rect 14160 11860 14170 11920
rect 14230 11910 14240 11920
rect 14880 11920 14960 11930
rect 14880 11910 14890 11920
rect 14230 11870 14890 11910
rect 14230 11860 14240 11870
rect 14160 11850 14240 11860
rect 14880 11860 14890 11870
rect 14950 11910 14960 11920
rect 15600 11920 15680 11930
rect 15600 11910 15610 11920
rect 14950 11870 15610 11910
rect 14950 11860 14960 11870
rect 14880 11850 14960 11860
rect 15600 11860 15610 11870
rect 15670 11860 15680 11920
rect 15600 11850 15680 11860
rect 11370 11590 11430 11620
rect 15130 11590 15190 11630
rect 8450 11580 13140 11590
rect 8450 11520 8460 11580
rect 8520 11520 10650 11580
rect 10710 11520 11370 11580
rect 11430 11520 12090 11580
rect 12150 11520 12810 11580
rect 12870 11520 13070 11580
rect 13130 11520 13140 11580
rect 8450 11510 13140 11520
rect 13420 11580 17650 11590
rect 13420 11520 13430 11580
rect 13490 11520 13690 11580
rect 13750 11520 14410 11580
rect 14470 11520 15130 11580
rect 15190 11520 15850 11580
rect 15910 11520 17580 11580
rect 17640 11520 17650 11580
rect 13420 11510 17650 11520
rect 10520 11470 16040 11480
rect 10520 11410 10530 11470
rect 10590 11410 10770 11470
rect 10830 11410 11010 11470
rect 11070 11410 11250 11470
rect 11310 11410 11490 11470
rect 11550 11410 11730 11470
rect 11790 11410 11970 11470
rect 12030 11410 12210 11470
rect 12270 11410 12450 11470
rect 12510 11410 12690 11470
rect 12750 11410 12930 11470
rect 12990 11410 13570 11470
rect 13630 11410 13810 11470
rect 13870 11410 14050 11470
rect 14110 11410 14290 11470
rect 14350 11410 14530 11470
rect 14590 11410 14770 11470
rect 14830 11410 15010 11470
rect 15070 11410 15250 11470
rect 15310 11410 15490 11470
rect 15550 11410 15730 11470
rect 15790 11410 15970 11470
rect 16030 11410 16040 11470
rect 10520 11390 16040 11410
rect 10520 11330 10530 11390
rect 10590 11330 10770 11390
rect 10830 11330 11010 11390
rect 11070 11330 11250 11390
rect 11310 11330 11490 11390
rect 11550 11330 11730 11390
rect 11790 11330 11970 11390
rect 12030 11330 12210 11390
rect 12270 11330 12450 11390
rect 12510 11330 12690 11390
rect 12750 11330 12930 11390
rect 12990 11330 13570 11390
rect 13630 11330 13810 11390
rect 13870 11330 14050 11390
rect 14110 11330 14290 11390
rect 14350 11330 14530 11390
rect 14590 11330 14770 11390
rect 14830 11330 15010 11390
rect 15070 11330 15250 11390
rect 15310 11330 15490 11390
rect 15550 11330 15730 11390
rect 15790 11330 15970 11390
rect 16030 11330 16040 11390
rect 10520 11310 16040 11330
rect 10520 11250 10530 11310
rect 10590 11250 10770 11310
rect 10830 11250 11010 11310
rect 11070 11250 11250 11310
rect 11310 11250 11490 11310
rect 11550 11250 11730 11310
rect 11790 11250 11970 11310
rect 12030 11250 12210 11310
rect 12270 11250 12450 11310
rect 12510 11250 12690 11310
rect 12750 11250 12930 11310
rect 12990 11250 13570 11310
rect 13630 11250 13810 11310
rect 13870 11250 14050 11310
rect 14110 11250 14290 11310
rect 14350 11250 14530 11310
rect 14590 11250 14770 11310
rect 14830 11250 15010 11310
rect 15070 11250 15250 11310
rect 15310 11250 15490 11310
rect 15550 11250 15730 11310
rect 15790 11250 15970 11310
rect 16030 11250 16040 11310
rect 10520 11240 16040 11250
rect 9570 11200 14760 11210
rect 9570 11140 9580 11200
rect 9640 11140 11810 11200
rect 11870 11140 13250 11200
rect 13310 11140 14690 11200
rect 14750 11140 14760 11200
rect 9570 11130 14760 11140
rect 9460 11090 15790 11100
rect 9460 11030 9470 11090
rect 9530 11030 12170 11090
rect 12230 11030 14330 11090
rect 14390 11030 15720 11090
rect 15780 11030 15790 11090
rect 9460 11020 15790 11030
rect 12520 10980 16320 10990
rect 12520 10920 12530 10980
rect 12590 10920 13970 10980
rect 14030 10920 15250 10980
rect 15310 10920 16250 10980
rect 16310 10920 16320 10980
rect 12520 10910 16320 10920
rect 12880 10870 16230 10880
rect 12880 10810 12890 10870
rect 12950 10810 13610 10870
rect 13670 10810 16160 10870
rect 16220 10810 16230 10870
rect 12880 10800 16230 10810
rect 11900 10760 14660 10770
rect 11960 10700 12080 10760
rect 12140 10700 12260 10760
rect 12320 10700 12440 10760
rect 12500 10700 12620 10760
rect 12680 10700 12800 10760
rect 12860 10700 12980 10760
rect 13040 10700 13160 10760
rect 13220 10700 13340 10760
rect 13400 10700 13430 10760
rect 13490 10700 13520 10760
rect 13580 10700 13700 10760
rect 13760 10700 13880 10760
rect 13940 10700 14060 10760
rect 14120 10700 14240 10760
rect 14300 10700 14420 10760
rect 14480 10700 14600 10760
rect 11900 10690 14660 10700
rect 15590 10560 15910 10570
rect 15590 10500 15600 10560
rect 15660 10500 15840 10560
rect 15900 10500 15910 10560
rect 15590 10490 15910 10500
rect 15240 10220 15320 10230
rect 15240 10160 15250 10220
rect 15310 10210 15320 10220
rect 15710 10220 15790 10230
rect 15710 10210 15720 10220
rect 15310 10170 15720 10210
rect 15310 10160 15320 10170
rect 15240 10150 15320 10160
rect 15710 10160 15720 10170
rect 15780 10160 15790 10220
rect 15710 10150 15790 10160
rect 11620 10020 16010 10030
rect 11620 9960 11630 10020
rect 11690 9960 11990 10020
rect 12050 9960 12350 10020
rect 12410 9960 12710 10020
rect 12770 9960 13070 10020
rect 13130 9960 13430 10020
rect 13490 9960 13790 10020
rect 13850 9960 14150 10020
rect 14210 9960 14510 10020
rect 14570 9960 14870 10020
rect 14930 9960 15500 10020
rect 15560 9960 15940 10020
rect 16000 9960 16010 10020
rect 11620 9940 16010 9960
rect 11620 9880 11630 9940
rect 11690 9880 11990 9940
rect 12050 9880 12350 9940
rect 12410 9880 12710 9940
rect 12770 9880 13070 9940
rect 13130 9880 13430 9940
rect 13490 9880 13790 9940
rect 13850 9880 14150 9940
rect 14210 9880 14510 9940
rect 14570 9880 14870 9940
rect 14930 9880 15500 9940
rect 15560 9880 15940 9940
rect 16000 9880 16010 9940
rect 11620 9860 16010 9880
rect 11620 9800 11630 9860
rect 11690 9800 11990 9860
rect 12050 9800 12350 9860
rect 12410 9800 12710 9860
rect 12770 9800 13070 9860
rect 13130 9800 13430 9860
rect 13490 9800 13790 9860
rect 13850 9800 14150 9860
rect 14210 9800 14510 9860
rect 14570 9800 14870 9860
rect 14930 9800 15500 9860
rect 15560 9800 15940 9860
rect 16000 9800 16010 9860
rect 11620 9790 16010 9800
rect 8450 9700 8460 9760
rect 8520 9750 14754 9760
rect 8520 9700 11808 9750
rect 8450 9698 11808 9700
rect 11860 9698 11918 9750
rect 11970 9698 12028 9750
rect 12080 9698 12138 9750
rect 12190 9698 12248 9750
rect 12300 9698 12358 9750
rect 12410 9698 12468 9750
rect 12520 9698 12578 9750
rect 12630 9698 12688 9750
rect 12740 9698 12798 9750
rect 12850 9698 13708 9750
rect 13760 9698 13818 9750
rect 13870 9698 13928 9750
rect 13980 9698 14038 9750
rect 14090 9698 14148 9750
rect 14200 9698 14258 9750
rect 14310 9698 14368 9750
rect 14420 9698 14478 9750
rect 14530 9698 14588 9750
rect 14640 9698 14698 9750
rect 14750 9698 14754 9750
rect 8450 9690 14754 9698
rect 11630 9420 14930 9430
rect 11630 9360 11640 9420
rect 11700 9360 11860 9420
rect 11920 9360 12080 9420
rect 12140 9360 12300 9420
rect 12360 9360 12520 9420
rect 12580 9360 12740 9420
rect 12800 9360 12960 9420
rect 13020 9360 13540 9420
rect 13600 9360 13760 9420
rect 13820 9360 13980 9420
rect 14040 9360 14200 9420
rect 14260 9360 14420 9420
rect 14480 9360 14640 9420
rect 14700 9360 14860 9420
rect 14920 9360 14930 9420
rect 11630 9350 14930 9360
rect 9680 9310 12920 9320
rect 9680 9250 9690 9310
rect 9750 9250 11750 9310
rect 11810 9250 11970 9310
rect 12030 9250 12190 9310
rect 12250 9250 12410 9310
rect 12470 9250 12630 9310
rect 12690 9250 12850 9310
rect 12910 9250 12920 9310
rect 9680 9240 12920 9250
rect 13640 9300 14820 9310
rect 13640 9240 13650 9300
rect 13710 9240 13870 9300
rect 13930 9240 14090 9300
rect 14150 9240 14310 9300
rect 14370 9240 14530 9300
rect 14590 9240 14750 9300
rect 14810 9240 14820 9300
rect 13640 9220 14820 9240
rect 13640 9160 13650 9220
rect 13710 9160 13870 9220
rect 13930 9160 14090 9220
rect 14150 9160 14310 9220
rect 14370 9160 14530 9220
rect 14590 9160 14750 9220
rect 14810 9160 14820 9220
rect 13640 9140 14820 9160
rect 13640 9080 13650 9140
rect 13710 9080 13870 9140
rect 13930 9080 14090 9140
rect 14150 9080 14310 9140
rect 14370 9080 14530 9140
rect 14590 9080 14750 9140
rect 14810 9080 14820 9140
rect 13640 9070 14820 9080
<< via2 >>
rect 18200 18790 18260 18850
rect 18660 18090 18720 18150
rect 18130 17390 18190 17450
rect 18800 16690 18860 16750
rect 19000 15990 19060 16050
rect 18800 15290 18860 15350
<< metal3 >>
rect 19120 18870 19580 19040
rect 19820 18870 20280 19040
rect 20520 18870 20980 19040
rect 21220 18870 21680 19040
rect 21920 18870 22380 19040
rect 22620 18870 23080 19040
rect 23320 18870 23780 19040
rect 24020 18870 24480 19040
rect 24720 18870 25180 19040
rect 25420 18870 25880 19040
rect 19120 18860 25880 18870
rect 18190 18850 25880 18860
rect 18190 18790 18200 18850
rect 18260 18790 25880 18850
rect 18190 18780 25880 18790
rect 19120 18770 25880 18780
rect 19120 18580 19580 18770
rect 19820 18580 20280 18770
rect 20520 18580 20980 18770
rect 21220 18580 21680 18770
rect 21920 18580 22380 18770
rect 22620 18580 23080 18770
rect 23320 18580 23780 18770
rect 24020 18580 24480 18770
rect 24720 18580 25180 18770
rect 25420 18580 25880 18770
rect 25600 18340 25700 18580
rect 19120 18170 19580 18340
rect 19820 18170 20280 18340
rect 20520 18170 20980 18340
rect 21220 18170 21680 18340
rect 21920 18170 22380 18340
rect 22620 18170 23080 18340
rect 23320 18170 23780 18340
rect 24020 18170 24480 18340
rect 24720 18170 25180 18340
rect 25420 18170 25880 18340
rect 18640 18160 18740 18170
rect 18640 18080 18650 18160
rect 18730 18080 18740 18160
rect 18640 18070 18740 18080
rect 19120 18070 25880 18170
rect 19120 17880 19580 18070
rect 19820 17880 20280 18070
rect 20520 17880 20980 18070
rect 21220 17880 21680 18070
rect 21920 17880 22380 18070
rect 22620 17880 23080 18070
rect 23320 17880 23780 18070
rect 24020 17880 24480 18070
rect 24720 17880 25180 18070
rect 25420 17880 25880 18070
rect 19120 17470 19580 17640
rect 19820 17470 20280 17640
rect 20520 17470 20980 17640
rect 21220 17470 21680 17640
rect 21920 17470 22380 17640
rect 22620 17470 23080 17640
rect 23320 17470 23780 17640
rect 24020 17470 24480 17640
rect 24720 17470 25180 17640
rect 25420 17470 25880 17640
rect 19120 17460 25880 17470
rect 18120 17450 25880 17460
rect 18120 17390 18130 17450
rect 18190 17390 25880 17450
rect 18120 17380 25880 17390
rect 19120 17370 25880 17380
rect 19120 17180 19580 17370
rect 19820 17180 20280 17370
rect 20520 17180 20980 17370
rect 21220 17180 21680 17370
rect 21920 17180 22380 17370
rect 22620 17180 23080 17370
rect 23320 17180 23780 17370
rect 24020 17180 24480 17370
rect 24720 17180 25180 17370
rect 25420 17180 25880 17370
rect 25600 16940 25700 17180
rect 19120 16770 19580 16940
rect 19820 16770 20280 16940
rect 20520 16770 20980 16940
rect 21220 16770 21680 16940
rect 21920 16770 22380 16940
rect 22620 16770 23080 16940
rect 23320 16770 23780 16940
rect 24020 16770 24480 16940
rect 24720 16770 25180 16940
rect 25420 16770 25880 16940
rect 18780 16760 18880 16770
rect 18780 16680 18790 16760
rect 18870 16680 18880 16760
rect 18780 16670 18880 16680
rect 19120 16670 25880 16770
rect 19120 16480 19580 16670
rect 19820 16480 20280 16670
rect 20520 16480 20980 16670
rect 21220 16480 21680 16670
rect 21920 16480 22380 16670
rect 22620 16480 23080 16670
rect 23320 16480 23780 16670
rect 24020 16480 24480 16670
rect 24720 16480 25180 16670
rect 25420 16480 25880 16670
rect 19120 16070 19580 16240
rect 19820 16070 20280 16240
rect 20520 16070 20980 16240
rect 21220 16070 21680 16240
rect 21920 16070 22380 16240
rect 22620 16070 23080 16240
rect 23320 16070 23780 16240
rect 24020 16070 24480 16240
rect 24720 16070 25180 16240
rect 25420 16070 25880 16240
rect 19120 16060 25880 16070
rect 18990 16050 25880 16060
rect 18990 15990 19000 16050
rect 19060 15990 25880 16050
rect 18990 15980 25880 15990
rect 19120 15970 25880 15980
rect 19120 15780 19580 15970
rect 19820 15780 20280 15970
rect 20520 15780 20980 15970
rect 21220 15780 21680 15970
rect 21920 15780 22380 15970
rect 22620 15780 23080 15970
rect 23320 15780 23780 15970
rect 24020 15780 24480 15970
rect 24720 15780 25180 15970
rect 25420 15780 25880 15970
rect 25600 15540 25700 15780
rect 19120 15370 19580 15540
rect 19820 15370 20280 15540
rect 20520 15370 20980 15540
rect 21220 15370 21680 15540
rect 21920 15370 22380 15540
rect 22620 15370 23080 15540
rect 23320 15370 23780 15540
rect 24020 15370 24480 15540
rect 24720 15370 25180 15540
rect 25420 15370 25880 15540
rect 18780 15360 18880 15370
rect 18780 15280 18790 15360
rect 18870 15280 18880 15360
rect 18780 15270 18880 15280
rect 19120 15270 25880 15370
rect 19120 15080 19580 15270
rect 19820 15080 20280 15270
rect 20520 15080 20980 15270
rect 21220 15080 21680 15270
rect 21920 15080 22380 15270
rect 22620 15080 23080 15270
rect 23320 15080 23780 15270
rect 24020 15080 24480 15270
rect 24720 15080 25180 15270
rect 25420 15080 25880 15270
<< via3 >>
rect 18650 18150 18730 18160
rect 18650 18090 18660 18150
rect 18660 18090 18720 18150
rect 18720 18090 18730 18150
rect 18650 18080 18730 18090
rect 18790 16750 18870 16760
rect 18790 16690 18800 16750
rect 18800 16690 18860 16750
rect 18860 16690 18870 16750
rect 18790 16680 18870 16690
rect 18790 15350 18870 15360
rect 18790 15290 18800 15350
rect 18800 15290 18860 15350
rect 18860 15290 18870 15350
rect 18790 15280 18870 15290
<< mimcap >>
rect 19150 18860 19550 19010
rect 19150 18780 19320 18860
rect 19400 18780 19550 18860
rect 19150 18610 19550 18780
rect 19850 18860 20250 19010
rect 19850 18780 20010 18860
rect 20090 18780 20250 18860
rect 19850 18610 20250 18780
rect 20550 18860 20950 19010
rect 20550 18780 20710 18860
rect 20790 18780 20950 18860
rect 20550 18610 20950 18780
rect 21250 18860 21650 19010
rect 21250 18780 21410 18860
rect 21490 18780 21650 18860
rect 21250 18610 21650 18780
rect 21950 18860 22350 19010
rect 21950 18780 22110 18860
rect 22190 18780 22350 18860
rect 21950 18610 22350 18780
rect 22650 18860 23050 19010
rect 22650 18780 22810 18860
rect 22890 18780 23050 18860
rect 22650 18610 23050 18780
rect 23350 18860 23750 19010
rect 23350 18780 23510 18860
rect 23590 18780 23750 18860
rect 23350 18610 23750 18780
rect 24050 18860 24450 19010
rect 24050 18780 24210 18860
rect 24290 18780 24450 18860
rect 24050 18610 24450 18780
rect 24750 18860 25150 19010
rect 24750 18780 24910 18860
rect 24990 18780 25150 18860
rect 24750 18610 25150 18780
rect 25450 18860 25850 19010
rect 25450 18780 25610 18860
rect 25690 18780 25850 18860
rect 25450 18610 25850 18780
rect 19150 18160 19550 18310
rect 19150 18080 19320 18160
rect 19400 18080 19550 18160
rect 19150 17910 19550 18080
rect 19850 18160 20250 18310
rect 19850 18080 20010 18160
rect 20090 18080 20250 18160
rect 19850 17910 20250 18080
rect 20550 18160 20950 18310
rect 20550 18080 20710 18160
rect 20790 18080 20950 18160
rect 20550 17910 20950 18080
rect 21250 18160 21650 18310
rect 21250 18080 21410 18160
rect 21490 18080 21650 18160
rect 21250 17910 21650 18080
rect 21950 18160 22350 18310
rect 21950 18080 22110 18160
rect 22190 18080 22350 18160
rect 21950 17910 22350 18080
rect 22650 18160 23050 18310
rect 22650 18080 22810 18160
rect 22890 18080 23050 18160
rect 22650 17910 23050 18080
rect 23350 18160 23750 18310
rect 23350 18080 23510 18160
rect 23590 18080 23750 18160
rect 23350 17910 23750 18080
rect 24050 18160 24450 18310
rect 24050 18080 24210 18160
rect 24290 18080 24450 18160
rect 24050 17910 24450 18080
rect 24750 18160 25150 18310
rect 24750 18080 24910 18160
rect 24990 18080 25150 18160
rect 24750 17910 25150 18080
rect 25450 18160 25850 18310
rect 25450 18080 25610 18160
rect 25690 18080 25850 18160
rect 25450 17910 25850 18080
rect 19150 17460 19550 17610
rect 19150 17380 19320 17460
rect 19400 17380 19550 17460
rect 19150 17210 19550 17380
rect 19850 17460 20250 17610
rect 19850 17380 20010 17460
rect 20090 17380 20250 17460
rect 19850 17210 20250 17380
rect 20550 17460 20950 17610
rect 20550 17380 20710 17460
rect 20790 17380 20950 17460
rect 20550 17210 20950 17380
rect 21250 17460 21650 17610
rect 21250 17380 21410 17460
rect 21490 17380 21650 17460
rect 21250 17210 21650 17380
rect 21950 17460 22350 17610
rect 21950 17380 22110 17460
rect 22190 17380 22350 17460
rect 21950 17210 22350 17380
rect 22650 17460 23050 17610
rect 22650 17380 22810 17460
rect 22890 17380 23050 17460
rect 22650 17210 23050 17380
rect 23350 17460 23750 17610
rect 23350 17380 23510 17460
rect 23590 17380 23750 17460
rect 23350 17210 23750 17380
rect 24050 17460 24450 17610
rect 24050 17380 24210 17460
rect 24290 17380 24450 17460
rect 24050 17210 24450 17380
rect 24750 17460 25150 17610
rect 24750 17380 24910 17460
rect 24990 17380 25150 17460
rect 24750 17210 25150 17380
rect 25450 17460 25850 17610
rect 25450 17380 25610 17460
rect 25690 17380 25850 17460
rect 25450 17210 25850 17380
rect 19150 16760 19550 16910
rect 19150 16680 19320 16760
rect 19400 16680 19550 16760
rect 19150 16510 19550 16680
rect 19850 16760 20250 16910
rect 19850 16680 20010 16760
rect 20090 16680 20250 16760
rect 19850 16510 20250 16680
rect 20550 16760 20950 16910
rect 20550 16680 20710 16760
rect 20790 16680 20950 16760
rect 20550 16510 20950 16680
rect 21250 16760 21650 16910
rect 21250 16680 21410 16760
rect 21490 16680 21650 16760
rect 21250 16510 21650 16680
rect 21950 16760 22350 16910
rect 21950 16680 22110 16760
rect 22190 16680 22350 16760
rect 21950 16510 22350 16680
rect 22650 16760 23050 16910
rect 22650 16680 22810 16760
rect 22890 16680 23050 16760
rect 22650 16510 23050 16680
rect 23350 16760 23750 16910
rect 23350 16680 23510 16760
rect 23590 16680 23750 16760
rect 23350 16510 23750 16680
rect 24050 16760 24450 16910
rect 24050 16680 24210 16760
rect 24290 16680 24450 16760
rect 24050 16510 24450 16680
rect 24750 16760 25150 16910
rect 24750 16680 24910 16760
rect 24990 16680 25150 16760
rect 24750 16510 25150 16680
rect 25450 16760 25850 16910
rect 25450 16680 25610 16760
rect 25690 16680 25850 16760
rect 25450 16510 25850 16680
rect 19150 16060 19550 16210
rect 19150 15980 19320 16060
rect 19400 15980 19550 16060
rect 19150 15810 19550 15980
rect 19850 16060 20250 16210
rect 19850 15980 20010 16060
rect 20090 15980 20250 16060
rect 19850 15810 20250 15980
rect 20550 16060 20950 16210
rect 20550 15980 20710 16060
rect 20790 15980 20950 16060
rect 20550 15810 20950 15980
rect 21250 16060 21650 16210
rect 21250 15980 21410 16060
rect 21490 15980 21650 16060
rect 21250 15810 21650 15980
rect 21950 16060 22350 16210
rect 21950 15980 22110 16060
rect 22190 15980 22350 16060
rect 21950 15810 22350 15980
rect 22650 16060 23050 16210
rect 22650 15980 22810 16060
rect 22890 15980 23050 16060
rect 22650 15810 23050 15980
rect 23350 16060 23750 16210
rect 23350 15980 23510 16060
rect 23590 15980 23750 16060
rect 23350 15810 23750 15980
rect 24050 16060 24450 16210
rect 24050 15980 24210 16060
rect 24290 15980 24450 16060
rect 24050 15810 24450 15980
rect 24750 16060 25150 16210
rect 24750 15980 24910 16060
rect 24990 15980 25150 16060
rect 24750 15810 25150 15980
rect 25450 16060 25850 16210
rect 25450 15980 25610 16060
rect 25690 15980 25850 16060
rect 25450 15810 25850 15980
rect 19150 15360 19550 15510
rect 19150 15280 19320 15360
rect 19400 15280 19550 15360
rect 19150 15110 19550 15280
rect 19850 15360 20250 15510
rect 19850 15280 20010 15360
rect 20090 15280 20250 15360
rect 19850 15110 20250 15280
rect 20550 15360 20950 15510
rect 20550 15280 20710 15360
rect 20790 15280 20950 15360
rect 20550 15110 20950 15280
rect 21250 15360 21650 15510
rect 21250 15280 21410 15360
rect 21490 15280 21650 15360
rect 21250 15110 21650 15280
rect 21950 15360 22350 15510
rect 21950 15280 22110 15360
rect 22190 15280 22350 15360
rect 21950 15110 22350 15280
rect 22650 15360 23050 15510
rect 22650 15280 22810 15360
rect 22890 15280 23050 15360
rect 22650 15110 23050 15280
rect 23350 15360 23750 15510
rect 23350 15280 23510 15360
rect 23590 15280 23750 15360
rect 23350 15110 23750 15280
rect 24050 15360 24450 15510
rect 24050 15280 24210 15360
rect 24290 15280 24450 15360
rect 24050 15110 24450 15280
rect 24750 15360 25150 15510
rect 24750 15280 24910 15360
rect 24990 15280 25150 15360
rect 24750 15110 25150 15280
rect 25450 15360 25850 15510
rect 25450 15280 25610 15360
rect 25690 15280 25850 15360
rect 25450 15110 25850 15280
<< mimcapcontact >>
rect 19320 18780 19400 18860
rect 20010 18780 20090 18860
rect 20710 18780 20790 18860
rect 21410 18780 21490 18860
rect 22110 18780 22190 18860
rect 22810 18780 22890 18860
rect 23510 18780 23590 18860
rect 24210 18780 24290 18860
rect 24910 18780 24990 18860
rect 25610 18780 25690 18860
rect 19320 18080 19400 18160
rect 20010 18080 20090 18160
rect 20710 18080 20790 18160
rect 21410 18080 21490 18160
rect 22110 18080 22190 18160
rect 22810 18080 22890 18160
rect 23510 18080 23590 18160
rect 24210 18080 24290 18160
rect 24910 18080 24990 18160
rect 25610 18080 25690 18160
rect 19320 17380 19400 17460
rect 20010 17380 20090 17460
rect 20710 17380 20790 17460
rect 21410 17380 21490 17460
rect 22110 17380 22190 17460
rect 22810 17380 22890 17460
rect 23510 17380 23590 17460
rect 24210 17380 24290 17460
rect 24910 17380 24990 17460
rect 25610 17380 25690 17460
rect 19320 16680 19400 16760
rect 20010 16680 20090 16760
rect 20710 16680 20790 16760
rect 21410 16680 21490 16760
rect 22110 16680 22190 16760
rect 22810 16680 22890 16760
rect 23510 16680 23590 16760
rect 24210 16680 24290 16760
rect 24910 16680 24990 16760
rect 25610 16680 25690 16760
rect 19320 15980 19400 16060
rect 20010 15980 20090 16060
rect 20710 15980 20790 16060
rect 21410 15980 21490 16060
rect 22110 15980 22190 16060
rect 22810 15980 22890 16060
rect 23510 15980 23590 16060
rect 24210 15980 24290 16060
rect 24910 15980 24990 16060
rect 25610 15980 25690 16060
rect 19320 15280 19400 15360
rect 20010 15280 20090 15360
rect 20710 15280 20790 15360
rect 21410 15280 21490 15360
rect 22110 15280 22190 15360
rect 22810 15280 22890 15360
rect 23510 15280 23590 15360
rect 24210 15280 24290 15360
rect 24910 15280 24990 15360
rect 25610 15280 25690 15360
<< metal4 >>
rect 19310 18860 25700 18870
rect 19310 18780 19320 18860
rect 19400 18780 20010 18860
rect 20090 18780 20710 18860
rect 20790 18780 21410 18860
rect 21490 18780 22110 18860
rect 22190 18780 22810 18860
rect 22890 18780 23510 18860
rect 23590 18780 24210 18860
rect 24290 18780 24910 18860
rect 24990 18780 25610 18860
rect 25690 18780 25700 18860
rect 19310 18770 25700 18780
rect 25600 18170 25700 18770
rect 18640 18160 25700 18170
rect 18640 18080 18650 18160
rect 18730 18080 19320 18160
rect 19400 18080 20010 18160
rect 20090 18080 20710 18160
rect 20790 18080 21410 18160
rect 21490 18080 22110 18160
rect 22190 18080 22810 18160
rect 22890 18080 23510 18160
rect 23590 18080 24210 18160
rect 24290 18080 24910 18160
rect 24990 18080 25610 18160
rect 25690 18080 25700 18160
rect 18640 18070 25700 18080
rect 19310 17460 25700 17470
rect 19310 17380 19320 17460
rect 19400 17380 20010 17460
rect 20090 17380 20710 17460
rect 20790 17380 21410 17460
rect 21490 17380 22110 17460
rect 22190 17380 22810 17460
rect 22890 17380 23510 17460
rect 23590 17380 24210 17460
rect 24290 17380 24910 17460
rect 24990 17380 25610 17460
rect 25690 17380 25700 17460
rect 19310 17370 25700 17380
rect 25600 16770 25700 17370
rect 18780 16760 25700 16770
rect 18780 16680 18790 16760
rect 18870 16680 19320 16760
rect 19400 16680 20010 16760
rect 20090 16680 20710 16760
rect 20790 16680 21410 16760
rect 21490 16680 22110 16760
rect 22190 16680 22810 16760
rect 22890 16680 23510 16760
rect 23590 16680 24210 16760
rect 24290 16680 24910 16760
rect 24990 16680 25610 16760
rect 25690 16680 25700 16760
rect 18780 16670 25700 16680
rect 19310 16060 25700 16070
rect 19310 15980 19320 16060
rect 19400 15980 20010 16060
rect 20090 15980 20710 16060
rect 20790 15980 21410 16060
rect 21490 15980 22110 16060
rect 22190 15980 22810 16060
rect 22890 15980 23510 16060
rect 23590 15980 24210 16060
rect 24290 15980 24910 16060
rect 24990 15980 25610 16060
rect 25690 15980 25700 16060
rect 19310 15970 25700 15980
rect 25600 15370 25700 15970
rect 18780 15360 25700 15370
rect 18780 15280 18790 15360
rect 18870 15280 19320 15360
rect 19400 15280 20010 15360
rect 20090 15280 20710 15360
rect 20790 15280 21410 15360
rect 21490 15280 22110 15360
rect 22190 15280 22810 15360
rect 22890 15280 23510 15360
rect 23590 15280 24210 15360
rect 24290 15280 24910 15360
rect 24990 15280 25610 15360
rect 25690 15280 25700 15360
rect 18780 15270 25700 15280
<< labels >>
flabel metal2 13290 9690 13290 9690 5 FreeSans 1600 0 0 -800 PFET_GATE
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
