magic
tech sky130A
magscale 1 2
timestamp 1757392821
<< nwell >>
rect 43050 3340 45360 5570
<< pwell >>
rect 43050 1840 45170 3260
<< nmos >>
rect 43278 2840 43310 3040
rect 43798 2840 43830 3040
rect 44318 2840 44350 3040
rect 43280 2360 43310 2660
rect 43800 2360 43830 2660
rect 44320 2360 44350 2660
rect 43280 1980 43310 2180
rect 43800 1980 43830 2180
rect 44320 1980 44350 2180
rect 44920 1980 44950 2180
<< pmos >>
rect 43280 5030 43580 5430
rect 43800 5030 44100 5430
rect 44320 5030 44620 5430
rect 44840 5030 45140 5430
rect 43280 4140 43310 4740
rect 43800 4140 43830 4740
rect 44320 4140 44350 4740
rect 43278 3560 43310 3960
rect 43798 3560 43830 3960
rect 44318 3560 44350 3960
<< ndiff >>
rect 43198 3010 43278 3040
rect 43198 2970 43218 3010
rect 43258 2970 43278 3010
rect 43198 2910 43278 2970
rect 43198 2870 43218 2910
rect 43258 2870 43278 2910
rect 43198 2840 43278 2870
rect 43310 3010 43390 3040
rect 43310 2970 43330 3010
rect 43370 2970 43390 3010
rect 43310 2910 43390 2970
rect 43310 2870 43330 2910
rect 43370 2870 43390 2910
rect 43310 2840 43390 2870
rect 43718 3010 43798 3040
rect 43718 2970 43738 3010
rect 43778 2970 43798 3010
rect 43718 2910 43798 2970
rect 43718 2870 43738 2910
rect 43778 2870 43798 2910
rect 43718 2840 43798 2870
rect 43830 3010 43910 3040
rect 43830 2970 43850 3010
rect 43890 2970 43910 3010
rect 43830 2910 43910 2970
rect 43830 2870 43850 2910
rect 43890 2870 43910 2910
rect 43830 2840 43910 2870
rect 44238 3010 44318 3040
rect 44238 2970 44258 3010
rect 44298 2970 44318 3010
rect 44238 2910 44318 2970
rect 44238 2870 44258 2910
rect 44298 2870 44318 2910
rect 44238 2840 44318 2870
rect 44350 3010 44430 3040
rect 44350 2970 44370 3010
rect 44410 2970 44430 3010
rect 44350 2910 44430 2970
rect 44350 2870 44370 2910
rect 44410 2870 44430 2910
rect 44350 2840 44430 2870
rect 43200 2630 43280 2660
rect 43200 2590 43220 2630
rect 43260 2590 43280 2630
rect 43200 2530 43280 2590
rect 43200 2490 43220 2530
rect 43260 2490 43280 2530
rect 43200 2430 43280 2490
rect 43200 2390 43220 2430
rect 43260 2390 43280 2430
rect 43200 2360 43280 2390
rect 43310 2630 43390 2660
rect 43310 2590 43330 2630
rect 43370 2590 43390 2630
rect 43310 2530 43390 2590
rect 43310 2490 43330 2530
rect 43370 2490 43390 2530
rect 43310 2430 43390 2490
rect 43310 2390 43330 2430
rect 43370 2390 43390 2430
rect 43310 2360 43390 2390
rect 43720 2630 43800 2660
rect 43720 2590 43740 2630
rect 43780 2590 43800 2630
rect 43720 2530 43800 2590
rect 43720 2490 43740 2530
rect 43780 2490 43800 2530
rect 43720 2430 43800 2490
rect 43720 2390 43740 2430
rect 43780 2390 43800 2430
rect 43720 2360 43800 2390
rect 43830 2630 43910 2660
rect 43830 2590 43850 2630
rect 43890 2590 43910 2630
rect 43830 2530 43910 2590
rect 43830 2490 43850 2530
rect 43890 2490 43910 2530
rect 43830 2430 43910 2490
rect 43830 2390 43850 2430
rect 43890 2390 43910 2430
rect 43830 2360 43910 2390
rect 44240 2630 44320 2660
rect 44240 2590 44260 2630
rect 44300 2590 44320 2630
rect 44240 2530 44320 2590
rect 44240 2490 44260 2530
rect 44300 2490 44320 2530
rect 44240 2430 44320 2490
rect 44240 2390 44260 2430
rect 44300 2390 44320 2430
rect 44240 2360 44320 2390
rect 44350 2630 44430 2660
rect 44350 2590 44370 2630
rect 44410 2590 44430 2630
rect 44350 2530 44430 2590
rect 44350 2490 44370 2530
rect 44410 2490 44430 2530
rect 44350 2430 44430 2490
rect 44350 2390 44370 2430
rect 44410 2390 44430 2430
rect 44350 2360 44430 2390
rect 43200 2150 43280 2180
rect 43200 2110 43220 2150
rect 43260 2110 43280 2150
rect 43200 2050 43280 2110
rect 43200 2010 43220 2050
rect 43260 2010 43280 2050
rect 43200 1980 43280 2010
rect 43310 2150 43390 2180
rect 43310 2110 43330 2150
rect 43370 2110 43390 2150
rect 43310 2050 43390 2110
rect 43310 2010 43330 2050
rect 43370 2010 43390 2050
rect 43310 1980 43390 2010
rect 43720 2150 43800 2180
rect 43720 2110 43740 2150
rect 43780 2110 43800 2150
rect 43720 2050 43800 2110
rect 43720 2010 43740 2050
rect 43780 2010 43800 2050
rect 43720 1980 43800 2010
rect 43830 2150 43910 2180
rect 43830 2110 43850 2150
rect 43890 2110 43910 2150
rect 43830 2050 43910 2110
rect 43830 2010 43850 2050
rect 43890 2010 43910 2050
rect 43830 1980 43910 2010
rect 44240 2150 44320 2180
rect 44240 2110 44260 2150
rect 44300 2110 44320 2150
rect 44240 2050 44320 2110
rect 44240 2010 44260 2050
rect 44300 2010 44320 2050
rect 44240 1980 44320 2010
rect 44350 2150 44430 2180
rect 44350 2110 44370 2150
rect 44410 2110 44430 2150
rect 44350 2050 44430 2110
rect 44350 2010 44370 2050
rect 44410 2010 44430 2050
rect 44350 1980 44430 2010
rect 44840 2150 44920 2180
rect 44840 2110 44860 2150
rect 44900 2110 44920 2150
rect 44840 2050 44920 2110
rect 44840 2010 44860 2050
rect 44900 2010 44920 2050
rect 44840 1980 44920 2010
rect 44950 2150 45030 2180
rect 44950 2110 44970 2150
rect 45010 2110 45030 2150
rect 44950 2050 45030 2110
rect 44950 2010 44970 2050
rect 45010 2010 45030 2050
rect 44950 1980 45030 2010
<< pdiff >>
rect 43200 5400 43280 5430
rect 43200 5360 43220 5400
rect 43260 5360 43280 5400
rect 43200 5300 43280 5360
rect 43200 5260 43220 5300
rect 43260 5260 43280 5300
rect 43200 5200 43280 5260
rect 43200 5160 43220 5200
rect 43260 5160 43280 5200
rect 43200 5100 43280 5160
rect 43200 5060 43220 5100
rect 43260 5060 43280 5100
rect 43200 5030 43280 5060
rect 43580 5400 43660 5430
rect 43580 5360 43600 5400
rect 43640 5360 43660 5400
rect 43580 5300 43660 5360
rect 43580 5260 43600 5300
rect 43640 5260 43660 5300
rect 43580 5200 43660 5260
rect 43580 5160 43600 5200
rect 43640 5160 43660 5200
rect 43580 5100 43660 5160
rect 43580 5060 43600 5100
rect 43640 5060 43660 5100
rect 43580 5030 43660 5060
rect 43720 5400 43800 5430
rect 43720 5360 43740 5400
rect 43780 5360 43800 5400
rect 43720 5300 43800 5360
rect 43720 5260 43740 5300
rect 43780 5260 43800 5300
rect 43720 5200 43800 5260
rect 43720 5160 43740 5200
rect 43780 5160 43800 5200
rect 43720 5100 43800 5160
rect 43720 5060 43740 5100
rect 43780 5060 43800 5100
rect 43720 5030 43800 5060
rect 44100 5400 44180 5430
rect 44100 5360 44120 5400
rect 44160 5360 44180 5400
rect 44100 5300 44180 5360
rect 44100 5260 44120 5300
rect 44160 5260 44180 5300
rect 44100 5200 44180 5260
rect 44100 5160 44120 5200
rect 44160 5160 44180 5200
rect 44100 5100 44180 5160
rect 44100 5060 44120 5100
rect 44160 5060 44180 5100
rect 44100 5030 44180 5060
rect 44240 5400 44320 5430
rect 44240 5360 44260 5400
rect 44300 5360 44320 5400
rect 44240 5300 44320 5360
rect 44240 5260 44260 5300
rect 44300 5260 44320 5300
rect 44240 5200 44320 5260
rect 44240 5160 44260 5200
rect 44300 5160 44320 5200
rect 44240 5100 44320 5160
rect 44240 5060 44260 5100
rect 44300 5060 44320 5100
rect 44240 5030 44320 5060
rect 44620 5400 44700 5430
rect 44620 5360 44640 5400
rect 44680 5360 44700 5400
rect 44620 5300 44700 5360
rect 44620 5260 44640 5300
rect 44680 5260 44700 5300
rect 44620 5200 44700 5260
rect 44620 5160 44640 5200
rect 44680 5160 44700 5200
rect 44620 5100 44700 5160
rect 44620 5060 44640 5100
rect 44680 5060 44700 5100
rect 44620 5030 44700 5060
rect 44760 5400 44840 5430
rect 44760 5360 44780 5400
rect 44820 5360 44840 5400
rect 44760 5300 44840 5360
rect 44760 5260 44780 5300
rect 44820 5260 44840 5300
rect 44760 5200 44840 5260
rect 44760 5160 44780 5200
rect 44820 5160 44840 5200
rect 44760 5100 44840 5160
rect 44760 5060 44780 5100
rect 44820 5060 44840 5100
rect 44760 5030 44840 5060
rect 45140 5400 45220 5430
rect 45140 5360 45160 5400
rect 45200 5360 45220 5400
rect 45140 5300 45220 5360
rect 45140 5260 45160 5300
rect 45200 5260 45220 5300
rect 45140 5200 45220 5260
rect 45140 5160 45160 5200
rect 45200 5160 45220 5200
rect 45140 5100 45220 5160
rect 45140 5060 45160 5100
rect 45200 5060 45220 5100
rect 45140 5030 45220 5060
rect 43200 4710 43280 4740
rect 43200 4670 43220 4710
rect 43260 4670 43280 4710
rect 43200 4610 43280 4670
rect 43200 4570 43220 4610
rect 43260 4570 43280 4610
rect 43200 4510 43280 4570
rect 43200 4470 43220 4510
rect 43260 4470 43280 4510
rect 43200 4410 43280 4470
rect 43200 4370 43220 4410
rect 43260 4370 43280 4410
rect 43200 4310 43280 4370
rect 43200 4270 43220 4310
rect 43260 4270 43280 4310
rect 43200 4210 43280 4270
rect 43200 4170 43220 4210
rect 43260 4170 43280 4210
rect 43200 4140 43280 4170
rect 43310 4710 43390 4740
rect 43310 4670 43330 4710
rect 43370 4670 43390 4710
rect 43310 4610 43390 4670
rect 43310 4570 43330 4610
rect 43370 4570 43390 4610
rect 43310 4510 43390 4570
rect 43310 4470 43330 4510
rect 43370 4470 43390 4510
rect 43310 4410 43390 4470
rect 43310 4370 43330 4410
rect 43370 4370 43390 4410
rect 43310 4310 43390 4370
rect 43310 4270 43330 4310
rect 43370 4270 43390 4310
rect 43310 4210 43390 4270
rect 43310 4170 43330 4210
rect 43370 4170 43390 4210
rect 43310 4140 43390 4170
rect 43720 4710 43800 4740
rect 43720 4670 43740 4710
rect 43780 4670 43800 4710
rect 43720 4610 43800 4670
rect 43720 4570 43740 4610
rect 43780 4570 43800 4610
rect 43720 4510 43800 4570
rect 43720 4470 43740 4510
rect 43780 4470 43800 4510
rect 43720 4410 43800 4470
rect 43720 4370 43740 4410
rect 43780 4370 43800 4410
rect 43720 4310 43800 4370
rect 43720 4270 43740 4310
rect 43780 4270 43800 4310
rect 43720 4210 43800 4270
rect 43720 4170 43740 4210
rect 43780 4170 43800 4210
rect 43720 4140 43800 4170
rect 43830 4710 43910 4740
rect 43830 4670 43850 4710
rect 43890 4670 43910 4710
rect 43830 4610 43910 4670
rect 43830 4570 43850 4610
rect 43890 4570 43910 4610
rect 43830 4510 43910 4570
rect 43830 4470 43850 4510
rect 43890 4470 43910 4510
rect 43830 4410 43910 4470
rect 43830 4370 43850 4410
rect 43890 4370 43910 4410
rect 43830 4310 43910 4370
rect 43830 4270 43850 4310
rect 43890 4270 43910 4310
rect 43830 4210 43910 4270
rect 43830 4170 43850 4210
rect 43890 4170 43910 4210
rect 43830 4140 43910 4170
rect 44240 4710 44320 4740
rect 44240 4670 44260 4710
rect 44300 4670 44320 4710
rect 44240 4610 44320 4670
rect 44240 4570 44260 4610
rect 44300 4570 44320 4610
rect 44240 4510 44320 4570
rect 44240 4470 44260 4510
rect 44300 4470 44320 4510
rect 44240 4410 44320 4470
rect 44240 4370 44260 4410
rect 44300 4370 44320 4410
rect 44240 4310 44320 4370
rect 44240 4270 44260 4310
rect 44300 4270 44320 4310
rect 44240 4210 44320 4270
rect 44240 4170 44260 4210
rect 44300 4170 44320 4210
rect 44240 4140 44320 4170
rect 44350 4710 44430 4740
rect 44350 4670 44370 4710
rect 44410 4670 44430 4710
rect 44350 4610 44430 4670
rect 44350 4570 44370 4610
rect 44410 4570 44430 4610
rect 44350 4510 44430 4570
rect 44350 4470 44370 4510
rect 44410 4470 44430 4510
rect 44350 4410 44430 4470
rect 44350 4370 44370 4410
rect 44410 4370 44430 4410
rect 44350 4310 44430 4370
rect 44350 4270 44370 4310
rect 44410 4270 44430 4310
rect 44350 4210 44430 4270
rect 44350 4170 44370 4210
rect 44410 4170 44430 4210
rect 44350 4140 44430 4170
rect 43198 3930 43278 3960
rect 43198 3890 43218 3930
rect 43258 3890 43278 3930
rect 43198 3830 43278 3890
rect 43198 3790 43218 3830
rect 43258 3790 43278 3830
rect 43198 3730 43278 3790
rect 43198 3690 43218 3730
rect 43258 3690 43278 3730
rect 43198 3630 43278 3690
rect 43198 3590 43218 3630
rect 43258 3590 43278 3630
rect 43198 3560 43278 3590
rect 43310 3930 43390 3960
rect 43310 3890 43330 3930
rect 43370 3890 43390 3930
rect 43310 3830 43390 3890
rect 43310 3790 43330 3830
rect 43370 3790 43390 3830
rect 43310 3730 43390 3790
rect 43310 3690 43330 3730
rect 43370 3690 43390 3730
rect 43310 3630 43390 3690
rect 43310 3590 43330 3630
rect 43370 3590 43390 3630
rect 43310 3560 43390 3590
rect 43718 3930 43798 3960
rect 43718 3890 43738 3930
rect 43778 3890 43798 3930
rect 43718 3830 43798 3890
rect 43718 3790 43738 3830
rect 43778 3790 43798 3830
rect 43718 3730 43798 3790
rect 43718 3690 43738 3730
rect 43778 3690 43798 3730
rect 43718 3630 43798 3690
rect 43718 3590 43738 3630
rect 43778 3590 43798 3630
rect 43718 3560 43798 3590
rect 43830 3930 43910 3960
rect 43830 3890 43850 3930
rect 43890 3890 43910 3930
rect 43830 3830 43910 3890
rect 43830 3790 43850 3830
rect 43890 3790 43910 3830
rect 43830 3730 43910 3790
rect 43830 3690 43850 3730
rect 43890 3690 43910 3730
rect 43830 3630 43910 3690
rect 43830 3590 43850 3630
rect 43890 3590 43910 3630
rect 43830 3560 43910 3590
rect 44238 3930 44318 3960
rect 44238 3890 44258 3930
rect 44298 3890 44318 3930
rect 44238 3830 44318 3890
rect 44238 3790 44258 3830
rect 44298 3790 44318 3830
rect 44238 3730 44318 3790
rect 44238 3690 44258 3730
rect 44298 3690 44318 3730
rect 44238 3630 44318 3690
rect 44238 3590 44258 3630
rect 44298 3590 44318 3630
rect 44238 3560 44318 3590
rect 44350 3930 44430 3960
rect 44350 3890 44370 3930
rect 44410 3890 44430 3930
rect 44350 3830 44430 3890
rect 44350 3790 44370 3830
rect 44410 3790 44430 3830
rect 44350 3730 44430 3790
rect 44350 3690 44370 3730
rect 44410 3690 44430 3730
rect 44350 3630 44430 3690
rect 44350 3590 44370 3630
rect 44410 3590 44430 3630
rect 44350 3560 44430 3590
<< ndiffc >>
rect 43218 2970 43258 3010
rect 43218 2870 43258 2910
rect 43330 2970 43370 3010
rect 43330 2870 43370 2910
rect 43738 2970 43778 3010
rect 43738 2870 43778 2910
rect 43850 2970 43890 3010
rect 43850 2870 43890 2910
rect 44258 2970 44298 3010
rect 44258 2870 44298 2910
rect 44370 2970 44410 3010
rect 44370 2870 44410 2910
rect 43220 2590 43260 2630
rect 43220 2490 43260 2530
rect 43220 2390 43260 2430
rect 43330 2590 43370 2630
rect 43330 2490 43370 2530
rect 43330 2390 43370 2430
rect 43740 2590 43780 2630
rect 43740 2490 43780 2530
rect 43740 2390 43780 2430
rect 43850 2590 43890 2630
rect 43850 2490 43890 2530
rect 43850 2390 43890 2430
rect 44260 2590 44300 2630
rect 44260 2490 44300 2530
rect 44260 2390 44300 2430
rect 44370 2590 44410 2630
rect 44370 2490 44410 2530
rect 44370 2390 44410 2430
rect 43220 2110 43260 2150
rect 43220 2010 43260 2050
rect 43330 2110 43370 2150
rect 43330 2010 43370 2050
rect 43740 2110 43780 2150
rect 43740 2010 43780 2050
rect 43850 2110 43890 2150
rect 43850 2010 43890 2050
rect 44260 2110 44300 2150
rect 44260 2010 44300 2050
rect 44370 2110 44410 2150
rect 44370 2010 44410 2050
rect 44860 2110 44900 2150
rect 44860 2010 44900 2050
rect 44970 2110 45010 2150
rect 44970 2010 45010 2050
<< pdiffc >>
rect 43220 5360 43260 5400
rect 43220 5260 43260 5300
rect 43220 5160 43260 5200
rect 43220 5060 43260 5100
rect 43600 5360 43640 5400
rect 43600 5260 43640 5300
rect 43600 5160 43640 5200
rect 43600 5060 43640 5100
rect 43740 5360 43780 5400
rect 43740 5260 43780 5300
rect 43740 5160 43780 5200
rect 43740 5060 43780 5100
rect 44120 5360 44160 5400
rect 44120 5260 44160 5300
rect 44120 5160 44160 5200
rect 44120 5060 44160 5100
rect 44260 5360 44300 5400
rect 44260 5260 44300 5300
rect 44260 5160 44300 5200
rect 44260 5060 44300 5100
rect 44640 5360 44680 5400
rect 44640 5260 44680 5300
rect 44640 5160 44680 5200
rect 44640 5060 44680 5100
rect 44780 5360 44820 5400
rect 44780 5260 44820 5300
rect 44780 5160 44820 5200
rect 44780 5060 44820 5100
rect 45160 5360 45200 5400
rect 45160 5260 45200 5300
rect 45160 5160 45200 5200
rect 45160 5060 45200 5100
rect 43220 4670 43260 4710
rect 43220 4570 43260 4610
rect 43220 4470 43260 4510
rect 43220 4370 43260 4410
rect 43220 4270 43260 4310
rect 43220 4170 43260 4210
rect 43330 4670 43370 4710
rect 43330 4570 43370 4610
rect 43330 4470 43370 4510
rect 43330 4370 43370 4410
rect 43330 4270 43370 4310
rect 43330 4170 43370 4210
rect 43740 4670 43780 4710
rect 43740 4570 43780 4610
rect 43740 4470 43780 4510
rect 43740 4370 43780 4410
rect 43740 4270 43780 4310
rect 43740 4170 43780 4210
rect 43850 4670 43890 4710
rect 43850 4570 43890 4610
rect 43850 4470 43890 4510
rect 43850 4370 43890 4410
rect 43850 4270 43890 4310
rect 43850 4170 43890 4210
rect 44260 4670 44300 4710
rect 44260 4570 44300 4610
rect 44260 4470 44300 4510
rect 44260 4370 44300 4410
rect 44260 4270 44300 4310
rect 44260 4170 44300 4210
rect 44370 4670 44410 4710
rect 44370 4570 44410 4610
rect 44370 4470 44410 4510
rect 44370 4370 44410 4410
rect 44370 4270 44410 4310
rect 44370 4170 44410 4210
rect 43218 3890 43258 3930
rect 43218 3790 43258 3830
rect 43218 3690 43258 3730
rect 43218 3590 43258 3630
rect 43330 3890 43370 3930
rect 43330 3790 43370 3830
rect 43330 3690 43370 3730
rect 43330 3590 43370 3630
rect 43738 3890 43778 3930
rect 43738 3790 43778 3830
rect 43738 3690 43778 3730
rect 43738 3590 43778 3630
rect 43850 3890 43890 3930
rect 43850 3790 43890 3830
rect 43850 3690 43890 3730
rect 43850 3590 43890 3630
rect 44258 3890 44298 3930
rect 44258 3790 44298 3830
rect 44258 3690 44298 3730
rect 44258 3590 44298 3630
rect 44370 3890 44410 3930
rect 44370 3790 44410 3830
rect 44370 3690 44410 3730
rect 44370 3590 44410 3630
<< psubdiff >>
rect 43090 3180 44230 3220
rect 44370 3180 45130 3220
rect 43090 2660 43130 3180
rect 45090 2660 45130 3180
rect 43090 1920 43130 2450
rect 45090 1920 45130 2450
rect 43090 1880 44230 1920
rect 44370 1880 45130 1920
<< nsubdiff >>
rect 43090 5490 44110 5530
rect 44270 5490 45150 5530
rect 45220 5490 45320 5530
rect 43090 5060 43130 5490
rect 45280 5060 45320 5490
rect 43090 3420 43130 4730
rect 45280 3420 45320 4730
rect 43090 3380 44110 3420
rect 44270 3380 45320 3420
<< psubdiffcont >>
rect 44230 3180 44370 3220
rect 43090 2450 43130 2660
rect 45090 2450 45130 2660
rect 44230 1880 44370 1920
<< nsubdiffcont >>
rect 44110 5490 44270 5530
rect 45150 5490 45220 5530
rect 43090 4730 43130 5060
rect 45280 4730 45320 5060
rect 44110 3380 44270 3420
<< poly >>
rect 43280 5430 43580 5460
rect 43800 5430 44100 5460
rect 44320 5430 44620 5460
rect 44840 5430 45140 5460
rect 43280 5000 43580 5030
rect 43800 5000 44100 5030
rect 44320 5000 44620 5030
rect 44840 5000 45140 5030
rect 43390 4980 43470 5000
rect 43390 4940 43410 4980
rect 43450 4940 43470 4980
rect 43390 4920 43470 4940
rect 43910 4980 43990 5000
rect 43910 4940 43930 4980
rect 43970 4940 43990 4980
rect 43910 4920 43990 4940
rect 44430 4980 44510 5000
rect 44430 4940 44450 4980
rect 44490 4940 44510 4980
rect 44430 4920 44510 4940
rect 44960 4980 45020 5000
rect 44960 4940 44970 4980
rect 45010 4940 45020 4980
rect 44960 4920 45020 4940
rect 43280 4740 43310 4770
rect 43800 4740 43830 4770
rect 44320 4740 44350 4770
rect 43280 4110 43310 4140
rect 43800 4110 43830 4140
rect 44320 4110 44350 4140
rect 43280 4092 43338 4110
rect 43280 4058 43292 4092
rect 43326 4058 43338 4092
rect 43280 4040 43338 4058
rect 43800 4092 43858 4110
rect 43800 4058 43812 4092
rect 43846 4058 43858 4092
rect 43800 4040 43858 4058
rect 44320 4092 44378 4110
rect 44320 4058 44332 4092
rect 44366 4058 44378 4092
rect 44320 4040 44378 4058
rect 43278 3960 43310 3990
rect 43798 3960 43830 3990
rect 44318 3960 44350 3990
rect 43278 3530 43310 3560
rect 43798 3530 43830 3560
rect 44318 3530 44350 3560
rect 43252 3512 43310 3530
rect 43252 3478 43264 3512
rect 43298 3478 43310 3512
rect 43252 3460 43310 3478
rect 43772 3512 43830 3530
rect 43772 3478 43784 3512
rect 43818 3478 43830 3512
rect 43772 3460 43830 3478
rect 44292 3512 44350 3530
rect 44292 3478 44304 3512
rect 44338 3478 44350 3512
rect 44292 3460 44350 3478
rect 43252 3122 43310 3140
rect 43252 3088 43264 3122
rect 43298 3088 43310 3122
rect 43252 3070 43310 3088
rect 43772 3122 43830 3140
rect 43772 3088 43784 3122
rect 43818 3088 43830 3122
rect 43772 3070 43830 3088
rect 44292 3122 44350 3140
rect 44292 3088 44304 3122
rect 44338 3088 44350 3122
rect 44292 3070 44350 3088
rect 43278 3040 43310 3070
rect 43798 3040 43830 3070
rect 44318 3040 44350 3070
rect 43278 2810 43310 2840
rect 43798 2810 43830 2840
rect 44318 2810 44350 2840
rect 43280 2742 43338 2760
rect 43280 2708 43292 2742
rect 43326 2708 43338 2742
rect 43280 2690 43338 2708
rect 43800 2742 43858 2760
rect 43800 2708 43812 2742
rect 43846 2708 43858 2742
rect 43800 2690 43858 2708
rect 44320 2742 44378 2760
rect 44320 2708 44332 2742
rect 44366 2708 44378 2742
rect 44320 2690 44378 2708
rect 43280 2660 43310 2690
rect 43800 2660 43830 2690
rect 44320 2660 44350 2690
rect 43280 2330 43310 2360
rect 43800 2330 43830 2360
rect 44320 2330 44350 2360
rect 43266 2262 43324 2280
rect 43266 2228 43278 2262
rect 43312 2228 43324 2262
rect 43266 2210 43324 2228
rect 43786 2262 43844 2280
rect 43786 2228 43798 2262
rect 43832 2228 43844 2262
rect 43786 2210 43844 2228
rect 44306 2262 44364 2280
rect 44306 2228 44318 2262
rect 44352 2228 44364 2262
rect 44306 2210 44364 2228
rect 44874 2262 44950 2280
rect 44874 2228 44886 2262
rect 44920 2228 44950 2262
rect 44874 2210 44950 2228
rect 43280 2180 43310 2210
rect 43800 2180 43830 2210
rect 44320 2180 44350 2210
rect 44920 2180 44950 2210
rect 43280 1950 43310 1980
rect 43800 1950 43830 1980
rect 44320 1950 44350 1980
rect 44920 1950 44950 1980
<< polycont >>
rect 43410 4940 43450 4980
rect 43930 4940 43970 4980
rect 44450 4940 44490 4980
rect 44970 4940 45010 4980
rect 43292 4058 43326 4092
rect 43812 4058 43846 4092
rect 44332 4058 44366 4092
rect 43264 3478 43298 3512
rect 43784 3478 43818 3512
rect 44304 3478 44338 3512
rect 43264 3088 43298 3122
rect 43784 3088 43818 3122
rect 44304 3088 44338 3122
rect 43292 2708 43326 2742
rect 43812 2708 43846 2742
rect 44332 2708 44366 2742
rect 43278 2228 43312 2262
rect 43798 2228 43832 2262
rect 44318 2228 44352 2262
rect 44886 2228 44920 2262
<< locali >>
rect 43580 5530 43660 5550
rect 44100 5530 44180 5550
rect 44620 5530 44700 5550
rect 45140 5530 45220 5550
rect 43090 5490 43600 5530
rect 43640 5490 44110 5530
rect 44270 5490 44640 5530
rect 44680 5490 45150 5530
rect 45220 5490 45320 5530
rect 43090 5060 43130 5490
rect 43580 5470 43660 5490
rect 44100 5470 44180 5490
rect 44620 5470 44700 5490
rect 45140 5470 45220 5490
rect 43210 5400 43270 5420
rect 43210 5360 43220 5400
rect 43260 5360 43270 5400
rect 43210 5300 43270 5360
rect 43210 5260 43220 5300
rect 43260 5260 43270 5300
rect 43210 5200 43270 5260
rect 43210 5160 43220 5200
rect 43260 5160 43270 5200
rect 43210 5100 43270 5160
rect 43210 5060 43220 5100
rect 43260 5060 43270 5100
rect 43210 5040 43270 5060
rect 43590 5400 43650 5420
rect 43590 5360 43600 5400
rect 43640 5360 43650 5400
rect 43590 5300 43650 5360
rect 43590 5260 43600 5300
rect 43640 5260 43650 5300
rect 43590 5200 43650 5260
rect 43590 5160 43600 5200
rect 43640 5160 43650 5200
rect 43590 5100 43650 5160
rect 43590 5060 43600 5100
rect 43640 5060 43650 5100
rect 43590 5040 43650 5060
rect 43730 5400 43790 5420
rect 43730 5360 43740 5400
rect 43780 5360 43790 5400
rect 43730 5300 43790 5360
rect 43730 5260 43740 5300
rect 43780 5260 43790 5300
rect 43730 5200 43790 5260
rect 43730 5160 43740 5200
rect 43780 5160 43790 5200
rect 43730 5100 43790 5160
rect 43730 5060 43740 5100
rect 43780 5060 43790 5100
rect 43730 5040 43790 5060
rect 44110 5400 44170 5420
rect 44110 5360 44120 5400
rect 44160 5360 44170 5400
rect 44110 5300 44170 5360
rect 44110 5260 44120 5300
rect 44160 5260 44170 5300
rect 44110 5200 44170 5260
rect 44110 5160 44120 5200
rect 44160 5160 44170 5200
rect 44110 5100 44170 5160
rect 44110 5060 44120 5100
rect 44160 5060 44170 5100
rect 44110 5040 44170 5060
rect 44250 5400 44310 5420
rect 44250 5360 44260 5400
rect 44300 5360 44310 5400
rect 44250 5300 44310 5360
rect 44250 5260 44260 5300
rect 44300 5260 44310 5300
rect 44250 5200 44310 5260
rect 44250 5160 44260 5200
rect 44300 5160 44310 5200
rect 44250 5100 44310 5160
rect 44250 5060 44260 5100
rect 44300 5060 44310 5100
rect 44250 5040 44310 5060
rect 44630 5400 44690 5420
rect 44630 5360 44640 5400
rect 44680 5360 44690 5400
rect 44630 5300 44690 5360
rect 44630 5260 44640 5300
rect 44680 5260 44690 5300
rect 44630 5200 44690 5260
rect 44630 5160 44640 5200
rect 44680 5160 44690 5200
rect 44630 5100 44690 5160
rect 44630 5060 44640 5100
rect 44680 5060 44690 5100
rect 44630 5040 44690 5060
rect 44770 5400 44830 5420
rect 44770 5360 44780 5400
rect 44820 5360 44830 5400
rect 44770 5300 44830 5360
rect 44770 5260 44780 5300
rect 44820 5260 44830 5300
rect 44770 5200 44830 5260
rect 44770 5160 44780 5200
rect 44820 5160 44830 5200
rect 44770 5100 44830 5160
rect 44770 5060 44780 5100
rect 44820 5060 44830 5100
rect 44770 5040 44830 5060
rect 45150 5400 45210 5420
rect 45150 5360 45160 5400
rect 45200 5360 45210 5400
rect 45150 5300 45210 5360
rect 45150 5260 45160 5300
rect 45200 5260 45210 5300
rect 45150 5200 45210 5260
rect 45150 5160 45160 5200
rect 45200 5160 45210 5200
rect 45150 5100 45210 5160
rect 45150 5060 45160 5100
rect 45200 5060 45210 5100
rect 45150 5040 45210 5060
rect 45280 5060 45320 5490
rect 43390 4980 43470 5000
rect 43390 4940 43410 4980
rect 43450 4940 43470 4980
rect 43390 4920 43470 4940
rect 43910 4980 43990 5000
rect 43910 4940 43930 4980
rect 43970 4940 43990 4980
rect 43910 4920 43990 4940
rect 44430 4980 44510 5000
rect 44430 4940 44450 4980
rect 44490 4940 44510 4980
rect 44430 4920 44510 4940
rect 44960 4980 45020 5000
rect 44960 4940 44970 4980
rect 45010 4940 45020 4980
rect 44960 4920 45020 4940
rect 43090 3420 43130 4730
rect 43210 4710 43270 4730
rect 43210 4670 43220 4710
rect 43260 4670 43270 4710
rect 43210 4610 43270 4670
rect 43210 4570 43220 4610
rect 43260 4570 43270 4610
rect 43210 4510 43270 4570
rect 43210 4470 43220 4510
rect 43260 4470 43270 4510
rect 43210 4410 43270 4470
rect 43210 4370 43220 4410
rect 43260 4370 43270 4410
rect 43210 4310 43270 4370
rect 43210 4270 43220 4310
rect 43260 4270 43270 4310
rect 43210 4210 43270 4270
rect 43210 4170 43220 4210
rect 43260 4170 43270 4210
rect 43210 4150 43270 4170
rect 43320 4710 43380 4730
rect 43320 4670 43330 4710
rect 43370 4670 43380 4710
rect 43320 4610 43380 4670
rect 43320 4570 43330 4610
rect 43370 4570 43380 4610
rect 43320 4510 43380 4570
rect 43320 4470 43330 4510
rect 43370 4470 43380 4510
rect 43320 4410 43380 4470
rect 43320 4370 43330 4410
rect 43370 4370 43380 4410
rect 43320 4310 43380 4370
rect 43320 4270 43330 4310
rect 43370 4270 43380 4310
rect 43320 4210 43380 4270
rect 43320 4170 43330 4210
rect 43370 4170 43380 4210
rect 43320 4150 43380 4170
rect 43730 4710 43790 4730
rect 43730 4670 43740 4710
rect 43780 4670 43790 4710
rect 43730 4610 43790 4670
rect 43730 4570 43740 4610
rect 43780 4570 43790 4610
rect 43730 4510 43790 4570
rect 43730 4470 43740 4510
rect 43780 4470 43790 4510
rect 43730 4410 43790 4470
rect 43730 4370 43740 4410
rect 43780 4370 43790 4410
rect 43730 4310 43790 4370
rect 43730 4270 43740 4310
rect 43780 4270 43790 4310
rect 43730 4210 43790 4270
rect 43730 4170 43740 4210
rect 43780 4170 43790 4210
rect 43730 4150 43790 4170
rect 43840 4710 43900 4730
rect 43840 4670 43850 4710
rect 43890 4670 43900 4710
rect 43840 4610 43900 4670
rect 43840 4570 43850 4610
rect 43890 4570 43900 4610
rect 43840 4510 43900 4570
rect 43840 4470 43850 4510
rect 43890 4470 43900 4510
rect 43840 4410 43900 4470
rect 43840 4370 43850 4410
rect 43890 4370 43900 4410
rect 43840 4310 43900 4370
rect 43840 4270 43850 4310
rect 43890 4270 43900 4310
rect 43840 4210 43900 4270
rect 43840 4170 43850 4210
rect 43890 4170 43900 4210
rect 43840 4150 43900 4170
rect 44250 4710 44310 4730
rect 44250 4670 44260 4710
rect 44300 4670 44310 4710
rect 44250 4610 44310 4670
rect 44250 4570 44260 4610
rect 44300 4570 44310 4610
rect 44250 4510 44310 4570
rect 44250 4470 44260 4510
rect 44300 4470 44310 4510
rect 44250 4410 44310 4470
rect 44250 4370 44260 4410
rect 44300 4370 44310 4410
rect 44250 4310 44310 4370
rect 44250 4270 44260 4310
rect 44300 4270 44310 4310
rect 44250 4210 44310 4270
rect 44250 4170 44260 4210
rect 44300 4170 44310 4210
rect 44250 4150 44310 4170
rect 44360 4710 44420 4730
rect 44360 4670 44370 4710
rect 44410 4670 44420 4710
rect 44360 4610 44420 4670
rect 44360 4570 44370 4610
rect 44410 4570 44420 4610
rect 44360 4510 44420 4570
rect 44360 4470 44370 4510
rect 44410 4470 44420 4510
rect 44360 4410 44420 4470
rect 44360 4370 44370 4410
rect 44410 4370 44420 4410
rect 44360 4310 44420 4370
rect 44360 4270 44370 4310
rect 44410 4270 44420 4310
rect 44360 4210 44420 4270
rect 44360 4170 44370 4210
rect 44410 4170 44420 4210
rect 44360 4150 44420 4170
rect 43280 4092 43338 4110
rect 43280 4058 43292 4092
rect 43326 4058 43338 4092
rect 43280 4040 43338 4058
rect 43800 4092 43858 4110
rect 43800 4058 43812 4092
rect 43846 4058 43858 4092
rect 43800 4040 43858 4058
rect 44320 4092 44378 4110
rect 44320 4058 44332 4092
rect 44366 4058 44378 4092
rect 44320 4040 44378 4058
rect 43208 3930 43268 3950
rect 43208 3890 43218 3930
rect 43258 3890 43268 3930
rect 43208 3830 43268 3890
rect 43208 3790 43218 3830
rect 43258 3790 43268 3830
rect 43208 3730 43268 3790
rect 43208 3690 43218 3730
rect 43258 3690 43268 3730
rect 43208 3630 43268 3690
rect 43208 3590 43218 3630
rect 43258 3590 43268 3630
rect 43208 3570 43268 3590
rect 43320 3930 43380 3950
rect 43320 3890 43330 3930
rect 43370 3890 43380 3930
rect 43320 3830 43380 3890
rect 43320 3790 43330 3830
rect 43370 3790 43380 3830
rect 43320 3730 43380 3790
rect 43320 3690 43330 3730
rect 43370 3690 43380 3730
rect 43320 3630 43380 3690
rect 43320 3590 43330 3630
rect 43370 3590 43380 3630
rect 43320 3570 43380 3590
rect 43728 3930 43788 3950
rect 43728 3890 43738 3930
rect 43778 3890 43788 3930
rect 43728 3830 43788 3890
rect 43728 3790 43738 3830
rect 43778 3790 43788 3830
rect 43728 3730 43788 3790
rect 43728 3690 43738 3730
rect 43778 3690 43788 3730
rect 43728 3630 43788 3690
rect 43728 3590 43738 3630
rect 43778 3590 43788 3630
rect 43728 3570 43788 3590
rect 43840 3930 43900 3950
rect 43840 3890 43850 3930
rect 43890 3890 43900 3930
rect 43840 3830 43900 3890
rect 43840 3790 43850 3830
rect 43890 3790 43900 3830
rect 43840 3730 43900 3790
rect 43840 3690 43850 3730
rect 43890 3690 43900 3730
rect 43840 3630 43900 3690
rect 43840 3590 43850 3630
rect 43890 3590 43900 3630
rect 43840 3570 43900 3590
rect 44248 3930 44308 3950
rect 44248 3890 44258 3930
rect 44298 3890 44308 3930
rect 44248 3830 44308 3890
rect 44248 3790 44258 3830
rect 44298 3790 44308 3830
rect 44248 3730 44308 3790
rect 44248 3690 44258 3730
rect 44298 3690 44308 3730
rect 44248 3630 44308 3690
rect 44248 3590 44258 3630
rect 44298 3590 44308 3630
rect 44248 3570 44308 3590
rect 44360 3930 44420 3950
rect 44360 3890 44370 3930
rect 44410 3890 44420 3930
rect 44360 3830 44420 3890
rect 44360 3790 44370 3830
rect 44410 3790 44420 3830
rect 44360 3730 44420 3790
rect 44360 3690 44370 3730
rect 44410 3690 44420 3730
rect 44360 3630 44420 3690
rect 44360 3590 44370 3630
rect 44410 3590 44420 3630
rect 44360 3570 44420 3590
rect 43252 3512 43310 3530
rect 43252 3478 43264 3512
rect 43298 3478 43310 3512
rect 43252 3460 43310 3478
rect 43772 3512 43830 3530
rect 43772 3478 43784 3512
rect 43818 3478 43830 3512
rect 43772 3460 43830 3478
rect 44292 3512 44350 3530
rect 44292 3478 44304 3512
rect 44338 3478 44350 3512
rect 44292 3460 44350 3478
rect 45280 3420 45320 4730
rect 43090 3380 44110 3420
rect 44270 3380 45320 3420
rect 43090 3180 44230 3220
rect 44370 3180 45130 3220
rect 43090 2660 43130 3180
rect 43252 3122 43310 3140
rect 43252 3088 43264 3122
rect 43298 3088 43310 3122
rect 43252 3070 43310 3088
rect 43772 3122 43830 3140
rect 43772 3088 43784 3122
rect 43818 3088 43830 3122
rect 43772 3070 43830 3088
rect 44292 3122 44350 3140
rect 44292 3088 44304 3122
rect 44338 3088 44350 3122
rect 44292 3070 44350 3088
rect 43208 3010 43268 3030
rect 43208 2970 43218 3010
rect 43258 2970 43268 3010
rect 43208 2910 43268 2970
rect 43208 2870 43218 2910
rect 43258 2870 43268 2910
rect 43208 2850 43268 2870
rect 43320 3010 43380 3030
rect 43320 2970 43330 3010
rect 43370 2970 43380 3010
rect 43320 2910 43380 2970
rect 43320 2870 43330 2910
rect 43370 2870 43380 2910
rect 43320 2850 43380 2870
rect 43728 3010 43788 3030
rect 43728 2970 43738 3010
rect 43778 2970 43788 3010
rect 43728 2910 43788 2970
rect 43728 2870 43738 2910
rect 43778 2870 43788 2910
rect 43728 2850 43788 2870
rect 43840 3010 43900 3030
rect 43840 2970 43850 3010
rect 43890 2970 43900 3010
rect 43840 2910 43900 2970
rect 43840 2870 43850 2910
rect 43890 2870 43900 2910
rect 43840 2850 43900 2870
rect 44248 3010 44308 3030
rect 44248 2970 44258 3010
rect 44298 2970 44308 3010
rect 44248 2910 44308 2970
rect 44248 2870 44258 2910
rect 44298 2870 44308 2910
rect 44248 2850 44308 2870
rect 44360 3010 44420 3030
rect 44360 2970 44370 3010
rect 44410 2970 44420 3010
rect 44360 2910 44420 2970
rect 44360 2870 44370 2910
rect 44410 2870 44420 2910
rect 44360 2850 44420 2870
rect 43280 2742 43338 2760
rect 43280 2708 43292 2742
rect 43326 2708 43338 2742
rect 43280 2690 43338 2708
rect 43800 2742 43858 2760
rect 43800 2708 43812 2742
rect 43846 2708 43858 2742
rect 43800 2690 43858 2708
rect 44320 2742 44378 2760
rect 44320 2708 44332 2742
rect 44366 2708 44378 2742
rect 44320 2690 44378 2708
rect 45090 2660 45130 3180
rect 43090 1920 43130 2450
rect 43210 2630 43270 2650
rect 43210 2590 43220 2630
rect 43260 2590 43270 2630
rect 43210 2530 43270 2590
rect 43210 2490 43220 2530
rect 43260 2490 43270 2530
rect 43210 2430 43270 2490
rect 43210 2390 43220 2430
rect 43260 2390 43270 2430
rect 43210 2370 43270 2390
rect 43320 2630 43380 2650
rect 43320 2590 43330 2630
rect 43370 2590 43380 2630
rect 43320 2530 43380 2590
rect 43320 2490 43330 2530
rect 43370 2490 43380 2530
rect 43320 2430 43380 2490
rect 43320 2390 43330 2430
rect 43370 2390 43380 2430
rect 43320 2370 43380 2390
rect 43730 2630 43790 2650
rect 43730 2590 43740 2630
rect 43780 2590 43790 2630
rect 43730 2530 43790 2590
rect 43730 2490 43740 2530
rect 43780 2490 43790 2530
rect 43730 2430 43790 2490
rect 43730 2390 43740 2430
rect 43780 2390 43790 2430
rect 43730 2370 43790 2390
rect 43840 2630 43900 2650
rect 43840 2590 43850 2630
rect 43890 2590 43900 2630
rect 43840 2530 43900 2590
rect 43840 2490 43850 2530
rect 43890 2490 43900 2530
rect 43840 2430 43900 2490
rect 43840 2390 43850 2430
rect 43890 2390 43900 2430
rect 43840 2370 43900 2390
rect 44250 2630 44310 2650
rect 44250 2590 44260 2630
rect 44300 2590 44310 2630
rect 44250 2530 44310 2590
rect 44250 2490 44260 2530
rect 44300 2490 44310 2530
rect 44250 2430 44310 2490
rect 44250 2390 44260 2430
rect 44300 2390 44310 2430
rect 44250 2370 44310 2390
rect 44360 2630 44420 2650
rect 44360 2590 44370 2630
rect 44410 2590 44420 2630
rect 44360 2530 44420 2590
rect 44360 2490 44370 2530
rect 44410 2490 44420 2530
rect 44360 2430 44420 2490
rect 44360 2390 44370 2430
rect 44410 2390 44420 2430
rect 44360 2370 44420 2390
rect 43266 2262 43324 2280
rect 43266 2228 43278 2262
rect 43312 2228 43324 2262
rect 43266 2210 43324 2228
rect 43786 2262 43844 2280
rect 43786 2228 43798 2262
rect 43832 2228 43844 2262
rect 43786 2210 43844 2228
rect 44306 2262 44364 2280
rect 44306 2228 44318 2262
rect 44352 2228 44364 2262
rect 44306 2210 44364 2228
rect 44874 2262 44932 2280
rect 44874 2228 44886 2262
rect 44920 2228 44932 2262
rect 44874 2210 44932 2228
rect 43210 2150 43270 2170
rect 43210 2110 43220 2150
rect 43260 2110 43270 2150
rect 43210 2050 43270 2110
rect 43210 2010 43220 2050
rect 43260 2010 43270 2050
rect 43210 1990 43270 2010
rect 43320 2150 43380 2170
rect 43320 2110 43330 2150
rect 43370 2110 43380 2150
rect 43320 2050 43380 2110
rect 43320 2010 43330 2050
rect 43370 2010 43380 2050
rect 43320 1990 43380 2010
rect 43730 2150 43790 2170
rect 43730 2110 43740 2150
rect 43780 2110 43790 2150
rect 43730 2050 43790 2110
rect 43730 2010 43740 2050
rect 43780 2010 43790 2050
rect 43730 1990 43790 2010
rect 43840 2150 43900 2170
rect 43840 2110 43850 2150
rect 43890 2110 43900 2150
rect 43840 2050 43900 2110
rect 43840 2010 43850 2050
rect 43890 2010 43900 2050
rect 43840 1990 43900 2010
rect 44250 2150 44310 2170
rect 44250 2110 44260 2150
rect 44300 2110 44310 2150
rect 44250 2050 44310 2110
rect 44250 2010 44260 2050
rect 44300 2010 44310 2050
rect 44250 1990 44310 2010
rect 44360 2150 44420 2170
rect 44360 2110 44370 2150
rect 44410 2110 44420 2150
rect 44360 2050 44420 2110
rect 44360 2010 44370 2050
rect 44410 2010 44420 2050
rect 44360 1990 44420 2010
rect 44850 2150 44910 2170
rect 44850 2110 44860 2150
rect 44900 2110 44910 2150
rect 44850 2050 44910 2110
rect 44850 2010 44860 2050
rect 44900 2010 44910 2050
rect 44850 1990 44910 2010
rect 44960 2150 45020 2170
rect 44960 2110 44970 2150
rect 45010 2110 45020 2150
rect 44960 2050 45020 2110
rect 44960 2010 44970 2050
rect 45010 2010 45020 2050
rect 44960 1990 45020 2010
rect 43310 1920 43390 1940
rect 43830 1920 43910 1940
rect 44350 1920 44430 1940
rect 44840 1920 44920 1940
rect 45090 1920 45130 2450
rect 43090 1880 43330 1920
rect 43370 1880 43850 1920
rect 43890 1880 44230 1920
rect 44410 1880 44860 1920
rect 44900 1880 45130 1920
rect 43310 1860 43390 1880
rect 43830 1860 43910 1880
rect 44350 1860 44430 1880
rect 44840 1860 44920 1880
<< viali >>
rect 43600 5490 43640 5530
rect 44120 5490 44160 5530
rect 44640 5490 44680 5530
rect 45160 5490 45200 5530
rect 43220 5360 43260 5400
rect 43220 5260 43260 5300
rect 43220 5160 43260 5200
rect 43220 5060 43260 5100
rect 43600 5360 43640 5400
rect 43600 5260 43640 5300
rect 43600 5160 43640 5200
rect 43600 5060 43640 5100
rect 43740 5360 43780 5400
rect 43740 5260 43780 5300
rect 43740 5160 43780 5200
rect 43740 5060 43780 5100
rect 44120 5360 44160 5400
rect 44120 5260 44160 5300
rect 44120 5160 44160 5200
rect 44120 5060 44160 5100
rect 44260 5360 44300 5400
rect 44260 5260 44300 5300
rect 44260 5160 44300 5200
rect 44260 5060 44300 5100
rect 44640 5360 44680 5400
rect 44640 5260 44680 5300
rect 44640 5160 44680 5200
rect 44640 5060 44680 5100
rect 44780 5360 44820 5400
rect 44780 5260 44820 5300
rect 44780 5160 44820 5200
rect 44780 5060 44820 5100
rect 45160 5360 45200 5400
rect 45160 5260 45200 5300
rect 45160 5160 45200 5200
rect 45160 5060 45200 5100
rect 43410 4940 43450 4980
rect 43930 4940 43970 4980
rect 44450 4940 44490 4980
rect 44970 4940 45010 4980
rect 43220 4670 43260 4710
rect 43220 4570 43260 4610
rect 43220 4470 43260 4510
rect 43220 4370 43260 4410
rect 43220 4270 43260 4310
rect 43220 4170 43260 4210
rect 43330 4670 43370 4710
rect 43330 4570 43370 4610
rect 43330 4470 43370 4510
rect 43330 4370 43370 4410
rect 43330 4270 43370 4310
rect 43330 4170 43370 4210
rect 43740 4670 43780 4710
rect 43740 4570 43780 4610
rect 43740 4470 43780 4510
rect 43740 4370 43780 4410
rect 43740 4270 43780 4310
rect 43740 4170 43780 4210
rect 43850 4670 43890 4710
rect 43850 4570 43890 4610
rect 43850 4470 43890 4510
rect 43850 4370 43890 4410
rect 43850 4270 43890 4310
rect 43850 4170 43890 4210
rect 44260 4670 44300 4710
rect 44260 4570 44300 4610
rect 44260 4470 44300 4510
rect 44260 4370 44300 4410
rect 44260 4270 44300 4310
rect 44260 4170 44300 4210
rect 44370 4670 44410 4710
rect 44370 4570 44410 4610
rect 44370 4470 44410 4510
rect 44370 4370 44410 4410
rect 44370 4270 44410 4310
rect 44370 4170 44410 4210
rect 43292 4058 43326 4092
rect 43812 4058 43846 4092
rect 44332 4058 44366 4092
rect 43218 3890 43258 3930
rect 43218 3790 43258 3830
rect 43218 3690 43258 3730
rect 43218 3590 43258 3630
rect 43330 3890 43370 3930
rect 43330 3790 43370 3830
rect 43330 3690 43370 3730
rect 43330 3590 43370 3630
rect 43738 3890 43778 3930
rect 43738 3790 43778 3830
rect 43738 3690 43778 3730
rect 43738 3590 43778 3630
rect 43850 3890 43890 3930
rect 43850 3790 43890 3830
rect 43850 3690 43890 3730
rect 43850 3590 43890 3630
rect 44258 3890 44298 3930
rect 44258 3790 44298 3830
rect 44258 3690 44298 3730
rect 44258 3590 44298 3630
rect 44370 3890 44410 3930
rect 44370 3790 44410 3830
rect 44370 3690 44410 3730
rect 44370 3590 44410 3630
rect 43264 3478 43298 3512
rect 43784 3478 43818 3512
rect 44304 3478 44338 3512
rect 43264 3088 43298 3122
rect 43784 3088 43818 3122
rect 44304 3088 44338 3122
rect 43218 2970 43258 3010
rect 43218 2870 43258 2910
rect 43330 2970 43370 3010
rect 43330 2870 43370 2910
rect 43738 2970 43778 3010
rect 43738 2870 43778 2910
rect 43850 2970 43890 3010
rect 43850 2870 43890 2910
rect 44258 2970 44298 3010
rect 44258 2870 44298 2910
rect 44370 2970 44410 3010
rect 44370 2870 44410 2910
rect 43292 2708 43326 2742
rect 43812 2708 43846 2742
rect 44332 2708 44366 2742
rect 43220 2590 43260 2630
rect 43220 2490 43260 2530
rect 43220 2390 43260 2430
rect 43330 2590 43370 2630
rect 43330 2490 43370 2530
rect 43330 2390 43370 2430
rect 43740 2590 43780 2630
rect 43740 2490 43780 2530
rect 43740 2390 43780 2430
rect 43850 2590 43890 2630
rect 43850 2490 43890 2530
rect 43850 2390 43890 2430
rect 44260 2590 44300 2630
rect 44260 2490 44300 2530
rect 44260 2390 44300 2430
rect 44370 2590 44410 2630
rect 44370 2490 44410 2530
rect 44370 2390 44410 2430
rect 43278 2228 43312 2262
rect 43798 2228 43832 2262
rect 44318 2228 44352 2262
rect 44886 2228 44920 2262
rect 43220 2110 43260 2150
rect 43220 2010 43260 2050
rect 43330 2110 43370 2150
rect 43330 2010 43370 2050
rect 43740 2110 43780 2150
rect 43740 2010 43780 2050
rect 43850 2110 43890 2150
rect 43850 2010 43890 2050
rect 44260 2110 44300 2150
rect 44260 2010 44300 2050
rect 44370 2110 44410 2150
rect 44370 2010 44410 2050
rect 44860 2110 44900 2150
rect 44860 2010 44900 2050
rect 44970 2110 45010 2150
rect 44970 2010 45010 2050
rect 43330 1880 43370 1920
rect 43850 1880 43890 1920
rect 44370 1880 44410 1920
rect 44860 1880 44900 1920
<< metal1 >>
rect 43580 5640 43660 5650
rect 43580 5580 43590 5640
rect 43650 5580 43660 5640
rect 43580 5530 43660 5580
rect 43580 5490 43600 5530
rect 43640 5490 43660 5530
rect 43580 5470 43660 5490
rect 44100 5640 44180 5650
rect 44100 5580 44110 5640
rect 44170 5580 44180 5640
rect 44100 5530 44180 5580
rect 44100 5490 44120 5530
rect 44160 5490 44180 5530
rect 44100 5470 44180 5490
rect 44620 5640 44700 5650
rect 44620 5580 44630 5640
rect 44690 5580 44700 5640
rect 44620 5530 44700 5580
rect 44620 5490 44640 5530
rect 44680 5490 44700 5530
rect 44620 5470 44700 5490
rect 45140 5640 45220 5650
rect 45140 5580 45150 5640
rect 45210 5580 45220 5640
rect 45140 5530 45220 5580
rect 45140 5490 45160 5530
rect 45200 5490 45220 5530
rect 45140 5470 45220 5490
rect 43210 5400 43270 5420
rect 43210 5360 43220 5400
rect 43260 5360 43270 5400
rect 43210 5300 43270 5360
rect 43210 5260 43220 5300
rect 43260 5260 43270 5300
rect 43210 5200 43270 5260
rect 43210 5160 43220 5200
rect 43260 5160 43270 5200
rect 43210 5100 43270 5160
rect 43210 5060 43220 5100
rect 43260 5060 43270 5100
rect 43210 4710 43270 5060
rect 43590 5400 43650 5470
rect 43590 5360 43600 5400
rect 43640 5360 43650 5400
rect 43590 5300 43650 5360
rect 43590 5260 43600 5300
rect 43640 5260 43650 5300
rect 43590 5200 43650 5260
rect 43590 5160 43600 5200
rect 43640 5160 43650 5200
rect 43590 5100 43650 5160
rect 43590 5060 43600 5100
rect 43640 5060 43650 5100
rect 43390 4990 43470 5000
rect 43390 4930 43400 4990
rect 43460 4930 43470 4990
rect 43390 4920 43470 4930
rect 43590 4820 43650 5060
rect 43730 5400 43790 5420
rect 43730 5360 43740 5400
rect 43780 5360 43790 5400
rect 43730 5300 43790 5360
rect 43730 5260 43740 5300
rect 43780 5260 43790 5300
rect 43730 5200 43790 5260
rect 43730 5160 43740 5200
rect 43780 5160 43790 5200
rect 43730 5100 43790 5160
rect 43730 5060 43740 5100
rect 43780 5060 43790 5100
rect 43310 4810 43390 4820
rect 43310 4750 43320 4810
rect 43380 4750 43390 4810
rect 43310 4740 43390 4750
rect 43580 4810 43660 4820
rect 43580 4750 43590 4810
rect 43650 4750 43660 4810
rect 43580 4740 43660 4750
rect 43210 4670 43220 4710
rect 43260 4670 43270 4710
rect 43210 4610 43270 4670
rect 43210 4570 43220 4610
rect 43260 4570 43270 4610
rect 43210 4510 43270 4570
rect 43210 4470 43220 4510
rect 43260 4470 43270 4510
rect 43210 4410 43270 4470
rect 43210 4370 43220 4410
rect 43260 4370 43270 4410
rect 43210 4310 43270 4370
rect 43210 4270 43220 4310
rect 43260 4270 43270 4310
rect 43210 4210 43270 4270
rect 43210 4170 43220 4210
rect 43260 4170 43270 4210
rect 43210 4150 43270 4170
rect 43320 4710 43380 4740
rect 43320 4670 43330 4710
rect 43370 4670 43380 4710
rect 43320 4610 43380 4670
rect 43320 4570 43330 4610
rect 43370 4570 43380 4610
rect 43320 4510 43380 4570
rect 43320 4470 43330 4510
rect 43370 4470 43380 4510
rect 43320 4410 43380 4470
rect 43320 4370 43330 4410
rect 43370 4370 43380 4410
rect 43320 4310 43380 4370
rect 43320 4270 43330 4310
rect 43370 4270 43380 4310
rect 43320 4220 43380 4270
rect 43730 4710 43790 5060
rect 44110 5400 44170 5470
rect 44110 5360 44120 5400
rect 44160 5360 44170 5400
rect 44110 5300 44170 5360
rect 44110 5260 44120 5300
rect 44160 5260 44170 5300
rect 44110 5200 44170 5260
rect 44110 5160 44120 5200
rect 44160 5160 44170 5200
rect 44110 5100 44170 5160
rect 44110 5060 44120 5100
rect 44160 5060 44170 5100
rect 43910 4990 43990 5000
rect 43910 4930 43920 4990
rect 43980 4930 43990 4990
rect 43910 4920 43990 4930
rect 44110 4820 44170 5060
rect 44250 5400 44310 5420
rect 44250 5360 44260 5400
rect 44300 5360 44310 5400
rect 44250 5300 44310 5360
rect 44250 5260 44260 5300
rect 44300 5260 44310 5300
rect 44250 5200 44310 5260
rect 44250 5160 44260 5200
rect 44300 5160 44310 5200
rect 44250 5100 44310 5160
rect 44250 5060 44260 5100
rect 44300 5060 44310 5100
rect 43830 4810 43910 4820
rect 43830 4750 43840 4810
rect 43900 4750 43910 4810
rect 43830 4740 43910 4750
rect 44100 4810 44180 4820
rect 44100 4750 44110 4810
rect 44170 4750 44180 4810
rect 44100 4740 44180 4750
rect 43730 4670 43740 4710
rect 43780 4670 43790 4710
rect 43730 4610 43790 4670
rect 43730 4570 43740 4610
rect 43780 4570 43790 4610
rect 43730 4510 43790 4570
rect 43730 4470 43740 4510
rect 43780 4470 43790 4510
rect 43730 4410 43790 4470
rect 43730 4370 43740 4410
rect 43780 4370 43790 4410
rect 43730 4310 43790 4370
rect 43730 4270 43740 4310
rect 43780 4270 43790 4310
rect 43320 4150 43380 4160
rect 43410 4220 43490 4230
rect 43410 4160 43420 4220
rect 43480 4160 43490 4220
rect 43410 4150 43490 4160
rect 43210 3950 43250 4150
rect 43280 4100 43338 4110
rect 43280 4048 43284 4100
rect 43336 4048 43338 4100
rect 43280 4040 43338 4048
rect 43208 3930 43268 3950
rect 43208 3890 43218 3930
rect 43258 3890 43268 3930
rect 43208 3830 43268 3890
rect 43208 3790 43218 3830
rect 43258 3790 43268 3830
rect 43208 3730 43268 3790
rect 43208 3690 43218 3730
rect 43258 3690 43268 3730
rect 43208 3630 43268 3690
rect 43208 3590 43218 3630
rect 43258 3590 43268 3630
rect 43208 3570 43268 3590
rect 43320 3930 43380 3950
rect 43320 3890 43330 3930
rect 43370 3890 43380 3930
rect 43320 3830 43380 3890
rect 43320 3790 43330 3830
rect 43370 3790 43380 3830
rect 43320 3730 43380 3790
rect 43320 3690 43330 3730
rect 43370 3690 43380 3730
rect 43320 3630 43380 3690
rect 43320 3590 43330 3630
rect 43370 3590 43380 3630
rect 43320 3560 43380 3590
rect 43252 3512 43310 3530
rect 43252 3478 43264 3512
rect 43298 3478 43310 3512
rect 43252 3460 43310 3478
rect 43260 3420 43310 3460
rect 42810 3410 43050 3420
rect 42810 3350 42820 3410
rect 42880 3350 42900 3410
rect 42960 3350 42980 3410
rect 43040 3350 43050 3410
rect 42810 3330 43050 3350
rect 42810 3270 42820 3330
rect 42880 3270 42900 3330
rect 42960 3270 42980 3330
rect 43040 3270 43050 3330
rect 42810 3250 43050 3270
rect 42810 3190 42820 3250
rect 42880 3190 42900 3250
rect 42960 3190 42980 3250
rect 43040 3190 43050 3250
rect 42810 1830 43050 3190
rect 43250 3410 43310 3420
rect 43250 3330 43310 3350
rect 43250 3250 43310 3270
rect 43250 3180 43310 3190
rect 43260 3140 43310 3180
rect 43252 3122 43310 3140
rect 43252 3088 43264 3122
rect 43298 3088 43310 3122
rect 43252 3070 43310 3088
rect 43340 3420 43380 3560
rect 43340 3410 43400 3420
rect 43340 3330 43400 3350
rect 43340 3250 43400 3270
rect 43340 3180 43400 3190
rect 43340 3030 43380 3180
rect 43170 3010 43268 3030
rect 43170 2970 43218 3010
rect 43258 2970 43268 3010
rect 43170 2910 43268 2970
rect 43170 2870 43218 2910
rect 43258 2870 43268 2910
rect 43170 2850 43268 2870
rect 43320 3010 43380 3030
rect 43320 2970 43330 3010
rect 43370 2970 43380 3010
rect 43320 2910 43380 2970
rect 43320 2870 43330 2910
rect 43370 2870 43380 2910
rect 43320 2850 43380 2870
rect 43170 2800 43212 2850
rect 43170 2650 43210 2800
rect 43430 2770 43490 4150
rect 43730 4210 43790 4270
rect 43730 4170 43740 4210
rect 43780 4170 43790 4210
rect 43730 4150 43790 4170
rect 43840 4710 43900 4740
rect 43840 4670 43850 4710
rect 43890 4670 43900 4710
rect 43840 4610 43900 4670
rect 43840 4570 43850 4610
rect 43890 4570 43900 4610
rect 43840 4510 43900 4570
rect 43840 4470 43850 4510
rect 43890 4470 43900 4510
rect 43840 4410 43900 4470
rect 43840 4370 43850 4410
rect 43890 4370 43900 4410
rect 43840 4310 43900 4370
rect 43840 4270 43850 4310
rect 43890 4270 43900 4310
rect 43840 4220 43900 4270
rect 44250 4710 44310 5060
rect 44630 5400 44690 5470
rect 44630 5360 44640 5400
rect 44680 5360 44690 5400
rect 44630 5300 44690 5360
rect 44630 5260 44640 5300
rect 44680 5260 44690 5300
rect 44630 5200 44690 5260
rect 44630 5160 44640 5200
rect 44680 5160 44690 5200
rect 44630 5100 44690 5160
rect 44630 5060 44640 5100
rect 44680 5060 44690 5100
rect 44430 4990 44510 5000
rect 44430 4930 44440 4990
rect 44500 4930 44510 4990
rect 44430 4920 44510 4930
rect 44630 4820 44690 5060
rect 44770 5400 44830 5420
rect 44770 5360 44780 5400
rect 44820 5360 44830 5400
rect 44770 5300 44830 5360
rect 44770 5260 44780 5300
rect 44820 5260 44830 5300
rect 44770 5200 44830 5260
rect 44770 5160 44780 5200
rect 44820 5160 44830 5200
rect 44770 5100 44830 5160
rect 44770 5060 44780 5100
rect 44820 5060 44830 5100
rect 44770 4990 44830 5060
rect 45150 5400 45210 5470
rect 45150 5360 45160 5400
rect 45200 5360 45210 5400
rect 45150 5300 45210 5360
rect 45150 5260 45160 5300
rect 45200 5260 45210 5300
rect 45150 5200 45210 5260
rect 45150 5160 45160 5200
rect 45200 5160 45210 5200
rect 45150 5100 45210 5160
rect 45150 5060 45160 5100
rect 45200 5060 45210 5100
rect 45150 5040 45210 5060
rect 44770 4920 44830 4930
rect 44960 4990 45020 5000
rect 44350 4810 44430 4820
rect 44350 4750 44360 4810
rect 44420 4750 44430 4810
rect 44350 4740 44430 4750
rect 44620 4810 44700 4820
rect 44620 4750 44630 4810
rect 44690 4750 44700 4810
rect 44620 4740 44700 4750
rect 44250 4670 44260 4710
rect 44300 4670 44310 4710
rect 44250 4610 44310 4670
rect 44250 4570 44260 4610
rect 44300 4570 44310 4610
rect 44250 4510 44310 4570
rect 44250 4470 44260 4510
rect 44300 4470 44310 4510
rect 44250 4410 44310 4470
rect 44250 4370 44260 4410
rect 44300 4370 44310 4410
rect 44250 4310 44310 4370
rect 44250 4270 44260 4310
rect 44300 4270 44310 4310
rect 43840 4150 43900 4160
rect 43930 4220 44010 4230
rect 43930 4160 43940 4220
rect 44000 4160 44010 4220
rect 43930 4150 44010 4160
rect 43410 2760 43490 2770
rect 43280 2750 43338 2760
rect 43280 2698 43284 2750
rect 43336 2698 43338 2750
rect 43280 2690 43338 2698
rect 43410 2700 43420 2760
rect 43480 2700 43490 2760
rect 43410 2690 43490 2700
rect 43520 4100 43600 4110
rect 43520 4040 43530 4100
rect 43590 4040 43600 4100
rect 43170 2630 43270 2650
rect 43170 2590 43220 2630
rect 43260 2590 43270 2630
rect 43170 2530 43270 2590
rect 43170 2490 43220 2530
rect 43260 2490 43270 2530
rect 43170 2430 43270 2490
rect 43170 2390 43220 2430
rect 43260 2390 43270 2430
rect 43170 2370 43270 2390
rect 43320 2640 43420 2650
rect 43380 2580 43420 2640
rect 43320 2530 43420 2580
rect 43520 2640 43600 4040
rect 43730 3950 43770 4150
rect 43800 4100 43858 4110
rect 43800 4048 43804 4100
rect 43856 4048 43858 4100
rect 43800 4040 43858 4048
rect 43728 3930 43788 3950
rect 43728 3890 43738 3930
rect 43778 3890 43788 3930
rect 43728 3830 43788 3890
rect 43728 3790 43738 3830
rect 43778 3790 43788 3830
rect 43728 3730 43788 3790
rect 43728 3690 43738 3730
rect 43778 3690 43788 3730
rect 43728 3630 43788 3690
rect 43728 3590 43738 3630
rect 43778 3590 43788 3630
rect 43728 3570 43788 3590
rect 43840 3930 43900 3950
rect 43840 3890 43850 3930
rect 43890 3890 43900 3930
rect 43840 3830 43900 3890
rect 43840 3790 43850 3830
rect 43890 3790 43900 3830
rect 43840 3730 43900 3790
rect 43840 3690 43850 3730
rect 43890 3690 43900 3730
rect 43840 3630 43900 3690
rect 43840 3590 43850 3630
rect 43890 3590 43900 3630
rect 43840 3560 43900 3590
rect 43772 3512 43830 3530
rect 43772 3478 43784 3512
rect 43818 3478 43830 3512
rect 43772 3460 43830 3478
rect 43780 3420 43830 3460
rect 43770 3410 43830 3420
rect 43770 3330 43830 3350
rect 43770 3250 43830 3270
rect 43770 3180 43830 3190
rect 43780 3140 43830 3180
rect 43772 3122 43830 3140
rect 43772 3088 43784 3122
rect 43818 3088 43830 3122
rect 43772 3070 43830 3088
rect 43860 3420 43900 3560
rect 43860 3410 43920 3420
rect 43860 3330 43920 3350
rect 43860 3250 43920 3270
rect 43860 3180 43920 3190
rect 43860 3030 43900 3180
rect 43520 2580 43530 2640
rect 43590 2580 43600 2640
rect 43520 2570 43600 2580
rect 43690 3010 43788 3030
rect 43690 2970 43738 3010
rect 43778 2970 43788 3010
rect 43690 2910 43788 2970
rect 43690 2870 43738 2910
rect 43778 2870 43788 2910
rect 43690 2850 43788 2870
rect 43840 3010 43900 3030
rect 43840 2970 43850 3010
rect 43890 2970 43900 3010
rect 43840 2910 43900 2970
rect 43840 2870 43850 2910
rect 43890 2870 43900 2910
rect 43840 2850 43900 2870
rect 43690 2800 43732 2850
rect 43690 2650 43730 2800
rect 43950 2770 44010 4150
rect 44250 4210 44310 4270
rect 44250 4170 44260 4210
rect 44300 4170 44310 4210
rect 44250 4150 44310 4170
rect 44360 4710 44420 4740
rect 44360 4670 44370 4710
rect 44410 4670 44420 4710
rect 44360 4610 44420 4670
rect 44360 4570 44370 4610
rect 44410 4570 44420 4610
rect 44360 4510 44420 4570
rect 44360 4470 44370 4510
rect 44410 4470 44420 4510
rect 44360 4410 44420 4470
rect 44360 4370 44370 4410
rect 44410 4370 44420 4410
rect 44360 4310 44420 4370
rect 44360 4270 44370 4310
rect 44410 4270 44420 4310
rect 44360 4220 44420 4270
rect 44360 4150 44420 4160
rect 44450 4220 44530 4230
rect 44450 4160 44460 4220
rect 44520 4160 44530 4220
rect 44450 4150 44530 4160
rect 43930 2760 44010 2770
rect 43800 2750 43858 2760
rect 43800 2698 43804 2750
rect 43856 2698 43858 2750
rect 43800 2690 43858 2698
rect 43930 2700 43940 2760
rect 44000 2700 44010 2760
rect 43930 2690 44010 2700
rect 44040 4100 44120 4110
rect 44040 4040 44050 4100
rect 44110 4040 44120 4100
rect 43690 2630 43790 2650
rect 43690 2590 43740 2630
rect 43780 2590 43790 2630
rect 43320 2490 43330 2530
rect 43370 2490 43420 2530
rect 43320 2430 43420 2490
rect 43320 2390 43330 2430
rect 43370 2390 43420 2430
rect 43320 2370 43420 2390
rect 43170 2170 43210 2370
rect 43266 2270 43324 2280
rect 43266 2218 43270 2270
rect 43322 2218 43324 2270
rect 43266 2210 43324 2218
rect 43380 2170 43420 2370
rect 43170 2150 43270 2170
rect 43170 2110 43220 2150
rect 43260 2110 43270 2150
rect 43170 2050 43270 2110
rect 43170 2010 43220 2050
rect 43260 2010 43270 2050
rect 43170 1990 43270 2010
rect 43320 2150 43420 2170
rect 43320 2110 43330 2150
rect 43370 2110 43420 2150
rect 43320 2050 43420 2110
rect 43320 2010 43330 2050
rect 43370 2010 43420 2050
rect 43320 1990 43420 2010
rect 43690 2530 43790 2590
rect 43690 2490 43740 2530
rect 43780 2490 43790 2530
rect 43690 2430 43790 2490
rect 43690 2390 43740 2430
rect 43780 2390 43790 2430
rect 43690 2370 43790 2390
rect 43840 2640 43940 2650
rect 43900 2580 43940 2640
rect 43840 2530 43940 2580
rect 44040 2640 44120 4040
rect 44250 3950 44290 4150
rect 44320 4100 44378 4110
rect 44320 4048 44324 4100
rect 44376 4048 44378 4100
rect 44320 4040 44378 4048
rect 44248 3930 44308 3950
rect 44248 3890 44258 3930
rect 44298 3890 44308 3930
rect 44248 3830 44308 3890
rect 44248 3790 44258 3830
rect 44298 3790 44308 3830
rect 44248 3730 44308 3790
rect 44248 3690 44258 3730
rect 44298 3690 44308 3730
rect 44248 3630 44308 3690
rect 44248 3590 44258 3630
rect 44298 3590 44308 3630
rect 44248 3570 44308 3590
rect 44360 3930 44420 3950
rect 44360 3890 44370 3930
rect 44410 3890 44420 3930
rect 44360 3830 44420 3890
rect 44360 3790 44370 3830
rect 44410 3790 44420 3830
rect 44360 3730 44420 3790
rect 44360 3690 44370 3730
rect 44410 3690 44420 3730
rect 44360 3630 44420 3690
rect 44360 3590 44370 3630
rect 44410 3590 44420 3630
rect 44360 3560 44420 3590
rect 44292 3512 44350 3530
rect 44292 3478 44304 3512
rect 44338 3478 44350 3512
rect 44292 3460 44350 3478
rect 44300 3420 44350 3460
rect 44290 3410 44350 3420
rect 44290 3330 44350 3350
rect 44290 3250 44350 3270
rect 44290 3180 44350 3190
rect 44300 3140 44350 3180
rect 44292 3122 44350 3140
rect 44292 3088 44304 3122
rect 44338 3088 44350 3122
rect 44292 3070 44350 3088
rect 44380 3420 44420 3560
rect 44380 3410 44440 3420
rect 44380 3330 44440 3350
rect 44380 3250 44440 3270
rect 44380 3180 44440 3190
rect 44380 3030 44420 3180
rect 44040 2580 44050 2640
rect 44110 2580 44120 2640
rect 44040 2570 44120 2580
rect 44210 3010 44308 3030
rect 44210 2970 44258 3010
rect 44298 2970 44308 3010
rect 44210 2910 44308 2970
rect 44210 2870 44258 2910
rect 44298 2870 44308 2910
rect 44210 2850 44308 2870
rect 44360 3010 44420 3030
rect 44360 2970 44370 3010
rect 44410 2970 44420 3010
rect 44360 2910 44420 2970
rect 44360 2870 44370 2910
rect 44410 2870 44420 2910
rect 44360 2850 44420 2870
rect 44210 2800 44252 2850
rect 44210 2650 44250 2800
rect 44470 2770 44530 4150
rect 44450 2760 44530 2770
rect 44320 2750 44378 2760
rect 44320 2698 44324 2750
rect 44376 2698 44378 2750
rect 44320 2690 44378 2698
rect 44450 2700 44460 2760
rect 44520 2700 44530 2760
rect 44450 2690 44530 2700
rect 44560 4100 44640 4110
rect 44560 4040 44570 4100
rect 44630 4040 44640 4100
rect 44210 2630 44310 2650
rect 44210 2590 44260 2630
rect 44300 2590 44310 2630
rect 43840 2490 43850 2530
rect 43890 2490 43940 2530
rect 43840 2430 43940 2490
rect 43840 2390 43850 2430
rect 43890 2390 43940 2430
rect 43840 2370 43940 2390
rect 43690 2170 43730 2370
rect 43786 2270 43844 2280
rect 43786 2218 43790 2270
rect 43842 2218 43844 2270
rect 43786 2210 43844 2218
rect 43900 2170 43940 2370
rect 43690 2150 43790 2170
rect 43690 2110 43740 2150
rect 43780 2110 43790 2150
rect 43690 2050 43790 2110
rect 43690 2010 43740 2050
rect 43780 2010 43790 2050
rect 43690 1990 43790 2010
rect 43840 2150 43940 2170
rect 43840 2110 43850 2150
rect 43890 2110 43940 2150
rect 43840 2050 43940 2110
rect 43840 2010 43850 2050
rect 43890 2010 43940 2050
rect 43840 1990 43940 2010
rect 44210 2530 44310 2590
rect 44210 2490 44260 2530
rect 44300 2490 44310 2530
rect 44210 2430 44310 2490
rect 44210 2390 44260 2430
rect 44300 2390 44310 2430
rect 44210 2370 44310 2390
rect 44360 2640 44460 2650
rect 44420 2580 44460 2640
rect 44360 2530 44460 2580
rect 44560 2640 44640 4040
rect 44560 2580 44570 2640
rect 44630 2580 44640 2640
rect 44560 2570 44640 2580
rect 44360 2490 44370 2530
rect 44410 2490 44460 2530
rect 44360 2430 44460 2490
rect 44360 2390 44370 2430
rect 44410 2390 44460 2430
rect 44360 2370 44460 2390
rect 44210 2170 44250 2370
rect 44306 2270 44364 2280
rect 44306 2218 44310 2270
rect 44362 2218 44364 2270
rect 44306 2210 44364 2218
rect 44420 2170 44460 2370
rect 44874 2270 44932 2280
rect 44874 2218 44876 2270
rect 44928 2218 44932 2270
rect 44874 2210 44932 2218
rect 44210 2150 44310 2170
rect 44210 2110 44260 2150
rect 44300 2110 44310 2150
rect 44210 2050 44310 2110
rect 44210 2010 44260 2050
rect 44300 2010 44310 2050
rect 44210 1990 44310 2010
rect 44360 2150 44460 2170
rect 44360 2110 44370 2150
rect 44410 2110 44460 2150
rect 44360 2050 44460 2110
rect 44360 2010 44370 2050
rect 44410 2010 44460 2050
rect 44360 1990 44460 2010
rect 44850 2150 44910 2170
rect 44850 2110 44860 2150
rect 44900 2110 44910 2150
rect 44850 2050 44910 2110
rect 44850 2010 44860 2050
rect 44900 2010 44910 2050
rect 43320 1940 43380 1990
rect 43840 1940 43900 1990
rect 44360 1940 44420 1990
rect 44850 1940 44910 2010
rect 44960 2150 45020 4930
rect 44960 2110 44970 2150
rect 45010 2110 45020 2150
rect 44960 2050 45020 2110
rect 44960 2010 44970 2050
rect 45010 2010 45020 2050
rect 44960 1990 45020 2010
rect 45170 3410 45410 3420
rect 45170 3350 45180 3410
rect 45240 3350 45260 3410
rect 45320 3350 45340 3410
rect 45400 3350 45410 3410
rect 45170 3330 45410 3350
rect 45170 3270 45180 3330
rect 45240 3270 45260 3330
rect 45320 3270 45340 3330
rect 45400 3270 45410 3330
rect 45170 3250 45410 3270
rect 45170 3190 45180 3250
rect 45240 3190 45260 3250
rect 45320 3190 45340 3250
rect 45400 3190 45410 3250
rect 42810 1770 42820 1830
rect 42880 1770 42900 1830
rect 42960 1770 42980 1830
rect 43040 1770 43050 1830
rect 42810 1750 43050 1770
rect 42810 1690 42820 1750
rect 42880 1690 42900 1750
rect 42960 1690 42980 1750
rect 43040 1690 43050 1750
rect 42810 1670 43050 1690
rect 42810 1610 42820 1670
rect 42880 1610 42900 1670
rect 42960 1610 42980 1670
rect 43040 1610 43050 1670
rect 42810 1600 43050 1610
rect 43310 1920 43390 1940
rect 43310 1880 43330 1920
rect 43370 1880 43390 1920
rect 43310 1560 43390 1880
rect 43310 1500 43320 1560
rect 43380 1500 43390 1560
rect 43310 1490 43390 1500
rect 43830 1920 43910 1940
rect 43830 1880 43850 1920
rect 43890 1880 43910 1920
rect 43830 1560 43910 1880
rect 43830 1500 43840 1560
rect 43900 1500 43910 1560
rect 43830 1490 43910 1500
rect 44350 1920 44430 1940
rect 44350 1880 44370 1920
rect 44410 1880 44430 1920
rect 44350 1560 44430 1880
rect 44350 1500 44360 1560
rect 44420 1500 44430 1560
rect 44350 1490 44430 1500
rect 44840 1920 44920 1940
rect 44840 1880 44860 1920
rect 44900 1880 44920 1920
rect 44840 1560 44920 1880
rect 45170 1830 45410 3190
rect 45170 1770 45180 1830
rect 45240 1770 45260 1830
rect 45320 1770 45340 1830
rect 45400 1770 45410 1830
rect 45170 1750 45410 1770
rect 45170 1690 45180 1750
rect 45240 1690 45260 1750
rect 45320 1690 45340 1750
rect 45400 1690 45410 1750
rect 45170 1670 45410 1690
rect 45170 1610 45180 1670
rect 45240 1610 45260 1670
rect 45320 1610 45340 1670
rect 45400 1610 45410 1670
rect 45170 1600 45410 1610
rect 44840 1500 44850 1560
rect 44910 1500 44920 1560
rect 44840 1490 44920 1500
<< via1 >>
rect 43590 5580 43650 5640
rect 44110 5580 44170 5640
rect 44630 5580 44690 5640
rect 45150 5580 45210 5640
rect 43400 4980 43460 4990
rect 43400 4940 43410 4980
rect 43410 4940 43450 4980
rect 43450 4940 43460 4980
rect 43400 4930 43460 4940
rect 43320 4750 43380 4810
rect 43590 4750 43650 4810
rect 43920 4980 43980 4990
rect 43920 4940 43930 4980
rect 43930 4940 43970 4980
rect 43970 4940 43980 4980
rect 43920 4930 43980 4940
rect 43840 4750 43900 4810
rect 44110 4750 44170 4810
rect 43320 4210 43380 4220
rect 43320 4170 43330 4210
rect 43330 4170 43370 4210
rect 43370 4170 43380 4210
rect 43320 4160 43380 4170
rect 43420 4160 43480 4220
rect 43284 4092 43336 4100
rect 43284 4058 43292 4092
rect 43292 4058 43326 4092
rect 43326 4058 43336 4092
rect 43284 4048 43336 4058
rect 42820 3350 42880 3410
rect 42900 3350 42960 3410
rect 42980 3350 43040 3410
rect 42820 3270 42880 3330
rect 42900 3270 42960 3330
rect 42980 3270 43040 3330
rect 42820 3190 42880 3250
rect 42900 3190 42960 3250
rect 42980 3190 43040 3250
rect 43250 3350 43310 3410
rect 43250 3270 43310 3330
rect 43250 3190 43310 3250
rect 43340 3350 43400 3410
rect 43340 3270 43400 3330
rect 43340 3190 43400 3250
rect 44440 4980 44500 4990
rect 44440 4940 44450 4980
rect 44450 4940 44490 4980
rect 44490 4940 44500 4980
rect 44440 4930 44500 4940
rect 44770 4930 44830 4990
rect 44960 4980 45020 4990
rect 44960 4940 44970 4980
rect 44970 4940 45010 4980
rect 45010 4940 45020 4980
rect 44960 4930 45020 4940
rect 44360 4750 44420 4810
rect 44630 4750 44690 4810
rect 43840 4210 43900 4220
rect 43840 4170 43850 4210
rect 43850 4170 43890 4210
rect 43890 4170 43900 4210
rect 43840 4160 43900 4170
rect 43940 4160 44000 4220
rect 43284 2742 43336 2750
rect 43284 2708 43292 2742
rect 43292 2708 43326 2742
rect 43326 2708 43336 2742
rect 43284 2698 43336 2708
rect 43420 2700 43480 2760
rect 43530 4040 43590 4100
rect 43320 2630 43380 2640
rect 43320 2590 43330 2630
rect 43330 2590 43370 2630
rect 43370 2590 43380 2630
rect 43320 2580 43380 2590
rect 43804 4092 43856 4100
rect 43804 4058 43812 4092
rect 43812 4058 43846 4092
rect 43846 4058 43856 4092
rect 43804 4048 43856 4058
rect 43770 3350 43830 3410
rect 43770 3270 43830 3330
rect 43770 3190 43830 3250
rect 43860 3350 43920 3410
rect 43860 3270 43920 3330
rect 43860 3190 43920 3250
rect 43530 2580 43590 2640
rect 44360 4210 44420 4220
rect 44360 4170 44370 4210
rect 44370 4170 44410 4210
rect 44410 4170 44420 4210
rect 44360 4160 44420 4170
rect 44460 4160 44520 4220
rect 43804 2742 43856 2750
rect 43804 2708 43812 2742
rect 43812 2708 43846 2742
rect 43846 2708 43856 2742
rect 43804 2698 43856 2708
rect 43940 2700 44000 2760
rect 44050 4040 44110 4100
rect 43270 2262 43322 2270
rect 43270 2228 43278 2262
rect 43278 2228 43312 2262
rect 43312 2228 43322 2262
rect 43270 2218 43322 2228
rect 43840 2630 43900 2640
rect 43840 2590 43850 2630
rect 43850 2590 43890 2630
rect 43890 2590 43900 2630
rect 43840 2580 43900 2590
rect 44324 4092 44376 4100
rect 44324 4058 44332 4092
rect 44332 4058 44366 4092
rect 44366 4058 44376 4092
rect 44324 4048 44376 4058
rect 44290 3350 44350 3410
rect 44290 3270 44350 3330
rect 44290 3190 44350 3250
rect 44380 3350 44440 3410
rect 44380 3270 44440 3330
rect 44380 3190 44440 3250
rect 44050 2580 44110 2640
rect 44324 2742 44376 2750
rect 44324 2708 44332 2742
rect 44332 2708 44366 2742
rect 44366 2708 44376 2742
rect 44324 2698 44376 2708
rect 44460 2700 44520 2760
rect 44570 4040 44630 4100
rect 43790 2262 43842 2270
rect 43790 2228 43798 2262
rect 43798 2228 43832 2262
rect 43832 2228 43842 2262
rect 43790 2218 43842 2228
rect 44360 2630 44420 2640
rect 44360 2590 44370 2630
rect 44370 2590 44410 2630
rect 44410 2590 44420 2630
rect 44360 2580 44420 2590
rect 44570 2580 44630 2640
rect 44310 2262 44362 2270
rect 44310 2228 44318 2262
rect 44318 2228 44352 2262
rect 44352 2228 44362 2262
rect 44310 2218 44362 2228
rect 44876 2262 44928 2270
rect 44876 2228 44886 2262
rect 44886 2228 44920 2262
rect 44920 2228 44928 2262
rect 44876 2218 44928 2228
rect 45180 3350 45240 3410
rect 45260 3350 45320 3410
rect 45340 3350 45400 3410
rect 45180 3270 45240 3330
rect 45260 3270 45320 3330
rect 45340 3270 45400 3330
rect 45180 3190 45240 3250
rect 45260 3190 45320 3250
rect 45340 3190 45400 3250
rect 42820 1770 42880 1830
rect 42900 1770 42960 1830
rect 42980 1770 43040 1830
rect 42820 1690 42880 1750
rect 42900 1690 42960 1750
rect 42980 1690 43040 1750
rect 42820 1610 42880 1670
rect 42900 1610 42960 1670
rect 42980 1610 43040 1670
rect 43320 1500 43380 1560
rect 43840 1500 43900 1560
rect 44360 1500 44420 1560
rect 45180 1770 45240 1830
rect 45260 1770 45320 1830
rect 45340 1770 45400 1830
rect 45180 1690 45240 1750
rect 45260 1690 45320 1750
rect 45340 1690 45400 1750
rect 45180 1610 45240 1670
rect 45260 1610 45320 1670
rect 45340 1610 45400 1670
rect 44850 1500 44910 1560
<< metal2 >>
rect 43580 5640 45220 5650
rect 43580 5580 43590 5640
rect 43650 5580 44110 5640
rect 44170 5580 44630 5640
rect 44690 5580 45150 5640
rect 45210 5580 45220 5640
rect 43580 5570 45220 5580
rect 43390 4990 45020 5000
rect 43390 4930 43400 4990
rect 43460 4930 43920 4990
rect 43980 4930 44440 4990
rect 44500 4930 44770 4990
rect 44830 4930 44960 4990
rect 43390 4920 45020 4930
rect 43310 4810 43660 4820
rect 43310 4750 43320 4810
rect 43380 4750 43590 4810
rect 43650 4750 43660 4810
rect 43310 4740 43660 4750
rect 43830 4810 44180 4820
rect 43830 4750 43840 4810
rect 43900 4750 44110 4810
rect 44170 4750 44180 4810
rect 43830 4740 44180 4750
rect 44350 4810 44700 4820
rect 44350 4750 44360 4810
rect 44420 4750 44630 4810
rect 44690 4750 44700 4810
rect 44350 4740 44700 4750
rect 43320 4220 43490 4230
rect 43380 4160 43420 4220
rect 43480 4160 43490 4220
rect 43320 4150 43490 4160
rect 43840 4220 44010 4230
rect 43900 4160 43940 4220
rect 44000 4160 44010 4220
rect 43840 4150 44010 4160
rect 44360 4220 44530 4230
rect 44420 4160 44460 4220
rect 44520 4160 44530 4220
rect 44360 4150 44530 4160
rect 43280 4100 43600 4110
rect 43280 4048 43284 4100
rect 43336 4048 43530 4100
rect 43280 4040 43530 4048
rect 43590 4040 43600 4100
rect 43800 4100 44120 4110
rect 43800 4048 43804 4100
rect 43856 4048 44050 4100
rect 43800 4040 44050 4048
rect 44110 4040 44120 4100
rect 44320 4100 44640 4110
rect 44320 4048 44324 4100
rect 44376 4048 44570 4100
rect 44320 4040 44570 4048
rect 44630 4040 44640 4100
rect 43520 4030 43600 4040
rect 44040 4030 44120 4040
rect 44560 4030 44640 4040
rect 42810 3410 43310 3420
rect 42810 3350 42820 3410
rect 42880 3350 42900 3410
rect 42960 3350 42980 3410
rect 43040 3350 43250 3410
rect 42810 3330 43310 3350
rect 42810 3270 42820 3330
rect 42880 3270 42900 3330
rect 42960 3270 42980 3330
rect 43040 3270 43250 3330
rect 42810 3250 43310 3270
rect 42810 3190 42820 3250
rect 42880 3190 42900 3250
rect 42960 3190 42980 3250
rect 43040 3190 43250 3250
rect 42810 3180 43310 3190
rect 43340 3410 43830 3420
rect 43400 3350 43770 3410
rect 43340 3330 43830 3350
rect 43400 3270 43770 3330
rect 43340 3250 43830 3270
rect 43400 3190 43770 3250
rect 43340 3180 43830 3190
rect 43860 3410 44350 3420
rect 43920 3350 44290 3410
rect 43860 3330 44350 3350
rect 43920 3270 44290 3330
rect 43860 3250 44350 3270
rect 43920 3190 44290 3250
rect 43860 3180 44350 3190
rect 44380 3410 45410 3420
rect 44440 3350 45180 3410
rect 45240 3350 45260 3410
rect 45320 3350 45340 3410
rect 45400 3350 45410 3410
rect 44380 3330 45410 3350
rect 44440 3270 45180 3330
rect 45240 3270 45260 3330
rect 45320 3270 45340 3330
rect 45400 3270 45410 3330
rect 44380 3250 45410 3270
rect 44440 3190 45180 3250
rect 45240 3190 45260 3250
rect 45320 3190 45340 3250
rect 45400 3190 45410 3250
rect 44380 3180 45410 3190
rect 43410 2760 43490 2770
rect 43930 2760 44010 2770
rect 44450 2760 44530 2770
rect 43280 2750 43420 2760
rect 43280 2698 43284 2750
rect 43336 2700 43420 2750
rect 43480 2700 43490 2760
rect 43336 2698 43490 2700
rect 43280 2690 43490 2698
rect 43800 2750 43940 2760
rect 43800 2698 43804 2750
rect 43856 2700 43940 2750
rect 44000 2700 44010 2760
rect 43856 2698 44010 2700
rect 43800 2690 44010 2698
rect 44320 2750 44460 2760
rect 44320 2698 44324 2750
rect 44376 2700 44460 2750
rect 44520 2700 44530 2760
rect 44376 2698 44530 2700
rect 44320 2690 44530 2698
rect 43320 2640 43600 2650
rect 43380 2580 43530 2640
rect 43590 2580 43600 2640
rect 43320 2570 43600 2580
rect 43840 2640 44120 2650
rect 43900 2580 44050 2640
rect 44110 2580 44120 2640
rect 43840 2570 44120 2580
rect 44360 2640 44640 2650
rect 44420 2580 44570 2640
rect 44630 2580 44640 2640
rect 44360 2570 44640 2580
rect 43265 2270 44950 2280
rect 43265 2218 43270 2270
rect 43322 2218 43790 2270
rect 43842 2218 44310 2270
rect 44362 2218 44876 2270
rect 44928 2218 44950 2270
rect 43265 2210 44950 2218
rect 42810 1830 45410 1840
rect 42810 1770 42820 1830
rect 42880 1770 42900 1830
rect 42960 1770 42980 1830
rect 43040 1770 45180 1830
rect 45240 1770 45260 1830
rect 45320 1770 45340 1830
rect 45400 1770 45410 1830
rect 42810 1750 45410 1770
rect 42810 1690 42820 1750
rect 42880 1690 42900 1750
rect 42960 1690 42980 1750
rect 43040 1690 45180 1750
rect 45240 1690 45260 1750
rect 45320 1690 45340 1750
rect 45400 1690 45410 1750
rect 42810 1670 45410 1690
rect 42810 1610 42820 1670
rect 42880 1610 42900 1670
rect 42960 1610 42980 1670
rect 43040 1610 45180 1670
rect 45240 1610 45260 1670
rect 45320 1610 45340 1670
rect 45400 1610 45410 1670
rect 42810 1600 45410 1610
rect 43310 1560 44920 1570
rect 43310 1500 43320 1560
rect 43380 1500 43840 1560
rect 43900 1500 44360 1560
rect 44420 1500 44850 1560
rect 44910 1500 44920 1560
rect 43310 1490 44920 1500
<< end >>
