magic
tech sky130A
timestamp 1757393171
<< nwell >>
rect 21130 1695 26385 1800
<< nmos >>
rect 21235 1555 21250 1605
rect 21290 1555 21305 1605
rect 21345 1555 21360 1605
rect 21400 1555 21415 1605
rect 21525 1555 21540 1605
rect 21580 1555 21595 1605
rect 21750 1555 21765 1605
rect 21805 1555 21820 1605
rect 21860 1555 21875 1605
rect 21915 1555 21930 1605
rect 22080 1555 22095 1605
rect 22135 1555 22150 1605
rect 22190 1555 22205 1605
rect 22245 1555 22260 1605
rect 22440 1555 22455 1605
rect 22495 1555 22510 1605
rect 22550 1555 22565 1605
rect 22605 1555 22620 1605
rect 22730 1555 22745 1605
rect 22785 1555 22800 1605
rect 23010 1555 23025 1605
rect 23190 1555 23205 1605
rect 23315 1555 23330 1605
rect 23370 1555 23385 1605
rect 23425 1555 23440 1605
rect 23480 1555 23495 1605
rect 23645 1555 23660 1605
rect 23700 1555 23715 1605
rect 23755 1555 23770 1605
rect 23920 1555 23935 1605
rect 23975 1555 23990 1605
rect 24030 1555 24045 1605
rect 24085 1555 24100 1605
rect 24250 1555 24265 1605
rect 24305 1555 24320 1605
rect 24360 1555 24375 1605
rect 24570 1510 24585 1560
rect 24625 1510 24640 1560
rect 24680 1510 24695 1560
rect 24735 1510 24750 1560
rect 24900 1510 24915 1560
rect 24955 1510 24970 1560
rect 25010 1510 25025 1560
rect 25220 1510 25235 1560
rect 25275 1510 25290 1560
rect 25330 1510 25345 1560
rect 25385 1510 25400 1560
rect 25550 1510 25565 1560
rect 25605 1510 25620 1560
rect 25660 1510 25675 1560
rect 25870 1510 25885 1560
rect 25925 1510 25940 1560
rect 25980 1510 25995 1560
rect 26035 1510 26050 1560
rect 26200 1510 26215 1560
rect 26255 1510 26270 1560
rect 26310 1510 26325 1560
<< pmos >>
rect 21315 1715 21330 1765
rect 21525 1715 21540 1765
rect 21580 1715 21595 1765
rect 21860 1715 21875 1765
rect 21915 1715 21930 1765
rect 22080 1715 22095 1765
rect 22135 1715 22150 1765
rect 22190 1715 22205 1765
rect 22520 1715 22535 1765
rect 22730 1715 22745 1765
rect 22785 1715 22800 1765
rect 22955 1715 22970 1765
rect 23010 1715 23025 1765
rect 23135 1715 23150 1765
rect 23190 1715 23205 1765
rect 23425 1715 23440 1765
rect 23480 1715 23495 1765
rect 23645 1715 23660 1765
rect 23700 1715 23715 1765
rect 23955 1715 23970 1765
rect 24125 1715 24140 1765
rect 24180 1715 24195 1765
rect 24305 1715 24320 1765
rect 24360 1715 24375 1765
rect 24605 1715 24620 1765
rect 24775 1715 24790 1765
rect 24830 1715 24845 1765
rect 24955 1715 24970 1765
rect 25010 1715 25025 1765
rect 25255 1715 25270 1765
rect 25425 1715 25440 1765
rect 25480 1715 25495 1765
rect 25605 1715 25620 1765
rect 25660 1715 25675 1765
rect 25905 1715 25920 1765
rect 26075 1715 26090 1765
rect 26130 1715 26145 1765
rect 26255 1715 26270 1765
rect 26310 1715 26325 1765
<< ndiff >>
rect 21195 1590 21235 1605
rect 21195 1570 21205 1590
rect 21225 1570 21235 1590
rect 21195 1555 21235 1570
rect 21250 1590 21290 1605
rect 21250 1570 21260 1590
rect 21280 1570 21290 1590
rect 21250 1555 21290 1570
rect 21305 1590 21345 1605
rect 21305 1570 21315 1590
rect 21335 1570 21345 1590
rect 21305 1555 21345 1570
rect 21360 1590 21400 1605
rect 21360 1570 21370 1590
rect 21390 1570 21400 1590
rect 21360 1555 21400 1570
rect 21415 1590 21455 1605
rect 21415 1570 21425 1590
rect 21445 1570 21455 1590
rect 21415 1555 21455 1570
rect 21485 1590 21525 1605
rect 21485 1570 21495 1590
rect 21515 1570 21525 1590
rect 21485 1555 21525 1570
rect 21540 1590 21580 1605
rect 21540 1570 21550 1590
rect 21570 1570 21580 1590
rect 21540 1555 21580 1570
rect 21595 1590 21635 1605
rect 21595 1570 21605 1590
rect 21625 1570 21635 1590
rect 21595 1555 21635 1570
rect 21710 1590 21750 1605
rect 21710 1570 21720 1590
rect 21740 1570 21750 1590
rect 21710 1555 21750 1570
rect 21765 1590 21805 1605
rect 21765 1570 21775 1590
rect 21795 1570 21805 1590
rect 21765 1555 21805 1570
rect 21820 1590 21860 1605
rect 21820 1570 21830 1590
rect 21850 1570 21860 1590
rect 21820 1555 21860 1570
rect 21875 1590 21915 1605
rect 21875 1570 21885 1590
rect 21905 1570 21915 1590
rect 21875 1555 21915 1570
rect 21930 1590 21970 1605
rect 21930 1570 21940 1590
rect 21960 1570 21970 1590
rect 21930 1555 21970 1570
rect 22040 1590 22080 1605
rect 22040 1570 22050 1590
rect 22070 1570 22080 1590
rect 22040 1555 22080 1570
rect 22095 1590 22135 1605
rect 22095 1570 22105 1590
rect 22125 1570 22135 1590
rect 22095 1555 22135 1570
rect 22150 1590 22190 1605
rect 22150 1570 22160 1590
rect 22180 1570 22190 1590
rect 22150 1555 22190 1570
rect 22205 1590 22245 1605
rect 22205 1570 22215 1590
rect 22235 1570 22245 1590
rect 22205 1555 22245 1570
rect 22260 1590 22300 1605
rect 22260 1570 22270 1590
rect 22290 1570 22300 1590
rect 22260 1555 22300 1570
rect 22400 1590 22440 1605
rect 22400 1570 22410 1590
rect 22430 1570 22440 1590
rect 22400 1555 22440 1570
rect 22455 1590 22495 1605
rect 22455 1570 22465 1590
rect 22485 1570 22495 1590
rect 22455 1555 22495 1570
rect 22510 1590 22550 1605
rect 22510 1570 22520 1590
rect 22540 1570 22550 1590
rect 22510 1555 22550 1570
rect 22565 1590 22605 1605
rect 22565 1570 22575 1590
rect 22595 1570 22605 1590
rect 22565 1555 22605 1570
rect 22620 1590 22660 1605
rect 22620 1570 22630 1590
rect 22650 1570 22660 1590
rect 22620 1555 22660 1570
rect 22690 1590 22730 1605
rect 22690 1570 22700 1590
rect 22720 1570 22730 1590
rect 22690 1555 22730 1570
rect 22745 1590 22785 1605
rect 22745 1570 22755 1590
rect 22775 1570 22785 1590
rect 22745 1555 22785 1570
rect 22800 1590 22840 1605
rect 22800 1570 22810 1590
rect 22830 1570 22840 1590
rect 22800 1555 22840 1570
rect 22970 1590 23010 1605
rect 22970 1570 22980 1590
rect 23000 1570 23010 1590
rect 22970 1555 23010 1570
rect 23025 1590 23065 1605
rect 23025 1570 23035 1590
rect 23055 1570 23065 1590
rect 23025 1555 23065 1570
rect 23150 1590 23190 1605
rect 23150 1570 23160 1590
rect 23180 1570 23190 1590
rect 23150 1555 23190 1570
rect 23205 1590 23245 1605
rect 23205 1570 23215 1590
rect 23235 1570 23245 1590
rect 23205 1555 23245 1570
rect 23275 1590 23315 1605
rect 23275 1570 23285 1590
rect 23305 1570 23315 1590
rect 23275 1555 23315 1570
rect 23330 1590 23370 1605
rect 23330 1570 23340 1590
rect 23360 1570 23370 1590
rect 23330 1555 23370 1570
rect 23385 1590 23425 1605
rect 23385 1570 23395 1590
rect 23415 1570 23425 1590
rect 23385 1555 23425 1570
rect 23440 1590 23480 1605
rect 23440 1570 23450 1590
rect 23470 1570 23480 1590
rect 23440 1555 23480 1570
rect 23495 1590 23535 1605
rect 23495 1570 23505 1590
rect 23525 1570 23535 1590
rect 23495 1555 23535 1570
rect 23605 1590 23645 1605
rect 23605 1570 23615 1590
rect 23635 1570 23645 1590
rect 23605 1555 23645 1570
rect 23660 1590 23700 1605
rect 23660 1570 23670 1590
rect 23690 1570 23700 1590
rect 23660 1555 23700 1570
rect 23715 1590 23755 1605
rect 23715 1570 23725 1590
rect 23745 1570 23755 1590
rect 23715 1555 23755 1570
rect 23770 1590 23810 1605
rect 23770 1570 23780 1590
rect 23800 1570 23810 1590
rect 23770 1555 23810 1570
rect 23880 1590 23920 1605
rect 23880 1570 23890 1590
rect 23910 1570 23920 1590
rect 23880 1555 23920 1570
rect 23935 1590 23975 1605
rect 23935 1570 23945 1590
rect 23965 1570 23975 1590
rect 23935 1555 23975 1570
rect 23990 1590 24030 1605
rect 23990 1570 24000 1590
rect 24020 1570 24030 1590
rect 23990 1555 24030 1570
rect 24045 1590 24085 1605
rect 24045 1570 24055 1590
rect 24075 1570 24085 1590
rect 24045 1555 24085 1570
rect 24100 1590 24140 1605
rect 24100 1570 24110 1590
rect 24130 1570 24140 1590
rect 24100 1555 24140 1570
rect 24210 1590 24250 1605
rect 24210 1570 24220 1590
rect 24240 1570 24250 1590
rect 24210 1555 24250 1570
rect 24265 1590 24305 1605
rect 24265 1570 24275 1590
rect 24295 1570 24305 1590
rect 24265 1555 24305 1570
rect 24320 1590 24360 1605
rect 24320 1570 24330 1590
rect 24350 1570 24360 1590
rect 24320 1555 24360 1570
rect 24375 1590 24415 1605
rect 24375 1570 24385 1590
rect 24405 1570 24415 1590
rect 24375 1555 24415 1570
rect 24530 1545 24570 1560
rect 24530 1525 24540 1545
rect 24560 1525 24570 1545
rect 24530 1510 24570 1525
rect 24585 1545 24625 1560
rect 24585 1525 24595 1545
rect 24615 1525 24625 1545
rect 24585 1510 24625 1525
rect 24640 1545 24680 1560
rect 24640 1525 24650 1545
rect 24670 1525 24680 1545
rect 24640 1510 24680 1525
rect 24695 1545 24735 1560
rect 24695 1525 24705 1545
rect 24725 1525 24735 1545
rect 24695 1510 24735 1525
rect 24750 1545 24790 1560
rect 24750 1525 24760 1545
rect 24780 1525 24790 1545
rect 24750 1510 24790 1525
rect 24860 1545 24900 1560
rect 24860 1525 24870 1545
rect 24890 1525 24900 1545
rect 24860 1510 24900 1525
rect 24915 1545 24955 1560
rect 24915 1525 24925 1545
rect 24945 1525 24955 1545
rect 24915 1510 24955 1525
rect 24970 1545 25010 1560
rect 24970 1525 24980 1545
rect 25000 1525 25010 1545
rect 24970 1510 25010 1525
rect 25025 1545 25065 1560
rect 25025 1525 25035 1545
rect 25055 1525 25065 1545
rect 25025 1510 25065 1525
rect 25180 1545 25220 1560
rect 25180 1525 25190 1545
rect 25210 1525 25220 1545
rect 25180 1510 25220 1525
rect 25235 1545 25275 1560
rect 25235 1525 25245 1545
rect 25265 1525 25275 1545
rect 25235 1510 25275 1525
rect 25290 1545 25330 1560
rect 25290 1525 25300 1545
rect 25320 1525 25330 1545
rect 25290 1510 25330 1525
rect 25345 1545 25385 1560
rect 25345 1525 25355 1545
rect 25375 1525 25385 1545
rect 25345 1510 25385 1525
rect 25400 1545 25440 1560
rect 25400 1525 25410 1545
rect 25430 1525 25440 1545
rect 25400 1510 25440 1525
rect 25510 1545 25550 1560
rect 25510 1525 25520 1545
rect 25540 1525 25550 1545
rect 25510 1510 25550 1525
rect 25565 1545 25605 1560
rect 25565 1525 25575 1545
rect 25595 1525 25605 1545
rect 25565 1510 25605 1525
rect 25620 1545 25660 1560
rect 25620 1525 25630 1545
rect 25650 1525 25660 1545
rect 25620 1510 25660 1525
rect 25675 1545 25715 1560
rect 25675 1525 25685 1545
rect 25705 1525 25715 1545
rect 25675 1510 25715 1525
rect 25830 1545 25870 1560
rect 25830 1525 25840 1545
rect 25860 1525 25870 1545
rect 25830 1510 25870 1525
rect 25885 1545 25925 1560
rect 25885 1525 25895 1545
rect 25915 1525 25925 1545
rect 25885 1510 25925 1525
rect 25940 1545 25980 1560
rect 25940 1525 25950 1545
rect 25970 1525 25980 1545
rect 25940 1510 25980 1525
rect 25995 1545 26035 1560
rect 25995 1525 26005 1545
rect 26025 1525 26035 1545
rect 25995 1510 26035 1525
rect 26050 1545 26090 1560
rect 26050 1525 26060 1545
rect 26080 1525 26090 1545
rect 26050 1510 26090 1525
rect 26160 1545 26200 1560
rect 26160 1525 26170 1545
rect 26190 1525 26200 1545
rect 26160 1510 26200 1525
rect 26215 1545 26255 1560
rect 26215 1525 26225 1545
rect 26245 1525 26255 1545
rect 26215 1510 26255 1525
rect 26270 1545 26310 1560
rect 26270 1525 26280 1545
rect 26300 1525 26310 1545
rect 26270 1510 26310 1525
rect 26325 1545 26365 1560
rect 26325 1525 26335 1545
rect 26355 1525 26365 1545
rect 26325 1510 26365 1525
<< pdiff >>
rect 21275 1750 21315 1765
rect 21275 1730 21285 1750
rect 21305 1730 21315 1750
rect 21275 1715 21315 1730
rect 21330 1750 21370 1765
rect 21330 1730 21340 1750
rect 21360 1730 21370 1750
rect 21330 1715 21370 1730
rect 21485 1750 21525 1765
rect 21485 1730 21495 1750
rect 21515 1730 21525 1750
rect 21485 1715 21525 1730
rect 21540 1750 21580 1765
rect 21540 1730 21550 1750
rect 21570 1730 21580 1750
rect 21540 1715 21580 1730
rect 21595 1750 21635 1765
rect 21595 1730 21605 1750
rect 21625 1730 21635 1750
rect 21595 1715 21635 1730
rect 21820 1750 21860 1765
rect 21820 1730 21830 1750
rect 21850 1730 21860 1750
rect 21820 1715 21860 1730
rect 21875 1750 21915 1765
rect 21875 1730 21885 1750
rect 21905 1730 21915 1750
rect 21875 1715 21915 1730
rect 21930 1750 21970 1765
rect 21930 1730 21940 1750
rect 21960 1730 21970 1750
rect 21930 1715 21970 1730
rect 22040 1750 22080 1765
rect 22040 1730 22050 1750
rect 22070 1730 22080 1750
rect 22040 1715 22080 1730
rect 22095 1750 22135 1765
rect 22095 1730 22105 1750
rect 22125 1730 22135 1750
rect 22095 1715 22135 1730
rect 22150 1750 22190 1765
rect 22150 1730 22160 1750
rect 22180 1730 22190 1750
rect 22150 1715 22190 1730
rect 22205 1750 22245 1765
rect 22205 1730 22215 1750
rect 22235 1730 22245 1750
rect 22205 1715 22245 1730
rect 22480 1750 22520 1765
rect 22480 1730 22490 1750
rect 22510 1730 22520 1750
rect 22480 1715 22520 1730
rect 22535 1750 22575 1765
rect 22535 1730 22545 1750
rect 22565 1730 22575 1750
rect 22535 1715 22575 1730
rect 22690 1750 22730 1765
rect 22690 1730 22700 1750
rect 22720 1730 22730 1750
rect 22690 1715 22730 1730
rect 22745 1750 22785 1765
rect 22745 1730 22755 1750
rect 22775 1730 22785 1750
rect 22745 1715 22785 1730
rect 22800 1750 22840 1765
rect 22800 1730 22810 1750
rect 22830 1730 22840 1750
rect 22800 1715 22840 1730
rect 22915 1750 22955 1765
rect 22915 1730 22925 1750
rect 22945 1730 22955 1750
rect 22915 1715 22955 1730
rect 22970 1750 23010 1765
rect 22970 1730 22980 1750
rect 23000 1730 23010 1750
rect 22970 1715 23010 1730
rect 23025 1750 23065 1765
rect 23025 1730 23035 1750
rect 23055 1730 23065 1750
rect 23025 1715 23065 1730
rect 23095 1750 23135 1765
rect 23095 1730 23105 1750
rect 23125 1730 23135 1750
rect 23095 1715 23135 1730
rect 23150 1750 23190 1765
rect 23150 1730 23160 1750
rect 23180 1730 23190 1750
rect 23150 1715 23190 1730
rect 23205 1750 23245 1765
rect 23205 1730 23215 1750
rect 23235 1730 23245 1750
rect 23205 1715 23245 1730
rect 23385 1750 23425 1765
rect 23385 1730 23395 1750
rect 23415 1730 23425 1750
rect 23385 1715 23425 1730
rect 23440 1750 23480 1765
rect 23440 1730 23450 1750
rect 23470 1730 23480 1750
rect 23440 1715 23480 1730
rect 23495 1750 23535 1765
rect 23495 1730 23505 1750
rect 23525 1730 23535 1750
rect 23495 1715 23535 1730
rect 23605 1750 23645 1765
rect 23605 1730 23615 1750
rect 23635 1730 23645 1750
rect 23605 1715 23645 1730
rect 23660 1750 23700 1765
rect 23660 1730 23670 1750
rect 23690 1730 23700 1750
rect 23660 1715 23700 1730
rect 23715 1750 23755 1765
rect 23715 1730 23725 1750
rect 23745 1730 23755 1750
rect 23715 1715 23755 1730
rect 23915 1750 23955 1765
rect 23915 1730 23925 1750
rect 23945 1730 23955 1750
rect 23915 1715 23955 1730
rect 23970 1750 24010 1765
rect 23970 1730 23980 1750
rect 24000 1730 24010 1750
rect 23970 1715 24010 1730
rect 24085 1750 24125 1765
rect 24085 1730 24095 1750
rect 24115 1730 24125 1750
rect 24085 1715 24125 1730
rect 24140 1750 24180 1765
rect 24140 1730 24150 1750
rect 24170 1730 24180 1750
rect 24140 1715 24180 1730
rect 24195 1750 24235 1765
rect 24195 1730 24205 1750
rect 24225 1730 24235 1750
rect 24195 1715 24235 1730
rect 24265 1750 24305 1765
rect 24265 1730 24275 1750
rect 24295 1730 24305 1750
rect 24265 1715 24305 1730
rect 24320 1750 24360 1765
rect 24320 1730 24330 1750
rect 24350 1730 24360 1750
rect 24320 1715 24360 1730
rect 24375 1750 24415 1765
rect 24375 1730 24385 1750
rect 24405 1730 24415 1750
rect 24375 1715 24415 1730
rect 24565 1750 24605 1765
rect 24565 1730 24575 1750
rect 24595 1730 24605 1750
rect 24565 1715 24605 1730
rect 24620 1750 24660 1765
rect 24620 1730 24630 1750
rect 24650 1730 24660 1750
rect 24620 1715 24660 1730
rect 24735 1750 24775 1765
rect 24735 1730 24745 1750
rect 24765 1730 24775 1750
rect 24735 1715 24775 1730
rect 24790 1750 24830 1765
rect 24790 1730 24800 1750
rect 24820 1730 24830 1750
rect 24790 1715 24830 1730
rect 24845 1750 24885 1765
rect 24845 1730 24855 1750
rect 24875 1730 24885 1750
rect 24845 1715 24885 1730
rect 24915 1750 24955 1765
rect 24915 1730 24925 1750
rect 24945 1730 24955 1750
rect 24915 1715 24955 1730
rect 24970 1750 25010 1765
rect 24970 1730 24980 1750
rect 25000 1730 25010 1750
rect 24970 1715 25010 1730
rect 25025 1750 25065 1765
rect 25025 1730 25035 1750
rect 25055 1730 25065 1750
rect 25025 1715 25065 1730
rect 25215 1750 25255 1765
rect 25215 1730 25225 1750
rect 25245 1730 25255 1750
rect 25215 1715 25255 1730
rect 25270 1750 25310 1765
rect 25270 1730 25280 1750
rect 25300 1730 25310 1750
rect 25270 1715 25310 1730
rect 25385 1750 25425 1765
rect 25385 1730 25395 1750
rect 25415 1730 25425 1750
rect 25385 1715 25425 1730
rect 25440 1750 25480 1765
rect 25440 1730 25450 1750
rect 25470 1730 25480 1750
rect 25440 1715 25480 1730
rect 25495 1750 25535 1765
rect 25495 1730 25505 1750
rect 25525 1730 25535 1750
rect 25495 1715 25535 1730
rect 25565 1750 25605 1765
rect 25565 1730 25575 1750
rect 25595 1730 25605 1750
rect 25565 1715 25605 1730
rect 25620 1750 25660 1765
rect 25620 1730 25630 1750
rect 25650 1730 25660 1750
rect 25620 1715 25660 1730
rect 25675 1750 25715 1765
rect 25675 1730 25685 1750
rect 25705 1730 25715 1750
rect 25675 1715 25715 1730
rect 25865 1750 25905 1765
rect 25865 1730 25875 1750
rect 25895 1730 25905 1750
rect 25865 1715 25905 1730
rect 25920 1750 25960 1765
rect 25920 1730 25930 1750
rect 25950 1730 25960 1750
rect 25920 1715 25960 1730
rect 26035 1750 26075 1765
rect 26035 1730 26045 1750
rect 26065 1730 26075 1750
rect 26035 1715 26075 1730
rect 26090 1750 26130 1765
rect 26090 1730 26100 1750
rect 26120 1730 26130 1750
rect 26090 1715 26130 1730
rect 26145 1750 26185 1765
rect 26145 1730 26155 1750
rect 26175 1730 26185 1750
rect 26145 1715 26185 1730
rect 26215 1750 26255 1765
rect 26215 1730 26225 1750
rect 26245 1730 26255 1750
rect 26215 1715 26255 1730
rect 26270 1750 26310 1765
rect 26270 1730 26280 1750
rect 26300 1730 26310 1750
rect 26270 1715 26310 1730
rect 26325 1750 26365 1765
rect 26325 1730 26335 1750
rect 26355 1730 26365 1750
rect 26325 1715 26365 1730
<< ndiffc >>
rect 21205 1570 21225 1590
rect 21260 1570 21280 1590
rect 21315 1570 21335 1590
rect 21370 1570 21390 1590
rect 21425 1570 21445 1590
rect 21495 1570 21515 1590
rect 21550 1570 21570 1590
rect 21605 1570 21625 1590
rect 21720 1570 21740 1590
rect 21775 1570 21795 1590
rect 21830 1570 21850 1590
rect 21885 1570 21905 1590
rect 21940 1570 21960 1590
rect 22050 1570 22070 1590
rect 22105 1570 22125 1590
rect 22160 1570 22180 1590
rect 22215 1570 22235 1590
rect 22270 1570 22290 1590
rect 22410 1570 22430 1590
rect 22465 1570 22485 1590
rect 22520 1570 22540 1590
rect 22575 1570 22595 1590
rect 22630 1570 22650 1590
rect 22700 1570 22720 1590
rect 22755 1570 22775 1590
rect 22810 1570 22830 1590
rect 22980 1570 23000 1590
rect 23035 1570 23055 1590
rect 23160 1570 23180 1590
rect 23215 1570 23235 1590
rect 23285 1570 23305 1590
rect 23340 1570 23360 1590
rect 23395 1570 23415 1590
rect 23450 1570 23470 1590
rect 23505 1570 23525 1590
rect 23615 1570 23635 1590
rect 23670 1570 23690 1590
rect 23725 1570 23745 1590
rect 23780 1570 23800 1590
rect 23890 1570 23910 1590
rect 23945 1570 23965 1590
rect 24000 1570 24020 1590
rect 24055 1570 24075 1590
rect 24110 1570 24130 1590
rect 24220 1570 24240 1590
rect 24275 1570 24295 1590
rect 24330 1570 24350 1590
rect 24385 1570 24405 1590
rect 24540 1525 24560 1545
rect 24595 1525 24615 1545
rect 24650 1525 24670 1545
rect 24705 1525 24725 1545
rect 24760 1525 24780 1545
rect 24870 1525 24890 1545
rect 24925 1525 24945 1545
rect 24980 1525 25000 1545
rect 25035 1525 25055 1545
rect 25190 1525 25210 1545
rect 25245 1525 25265 1545
rect 25300 1525 25320 1545
rect 25355 1525 25375 1545
rect 25410 1525 25430 1545
rect 25520 1525 25540 1545
rect 25575 1525 25595 1545
rect 25630 1525 25650 1545
rect 25685 1525 25705 1545
rect 25840 1525 25860 1545
rect 25895 1525 25915 1545
rect 25950 1525 25970 1545
rect 26005 1525 26025 1545
rect 26060 1525 26080 1545
rect 26170 1525 26190 1545
rect 26225 1525 26245 1545
rect 26280 1525 26300 1545
rect 26335 1525 26355 1545
<< pdiffc >>
rect 21285 1730 21305 1750
rect 21340 1730 21360 1750
rect 21495 1730 21515 1750
rect 21550 1730 21570 1750
rect 21605 1730 21625 1750
rect 21830 1730 21850 1750
rect 21885 1730 21905 1750
rect 21940 1730 21960 1750
rect 22050 1730 22070 1750
rect 22105 1730 22125 1750
rect 22160 1730 22180 1750
rect 22215 1730 22235 1750
rect 22490 1730 22510 1750
rect 22545 1730 22565 1750
rect 22700 1730 22720 1750
rect 22755 1730 22775 1750
rect 22810 1730 22830 1750
rect 22925 1730 22945 1750
rect 22980 1730 23000 1750
rect 23035 1730 23055 1750
rect 23105 1730 23125 1750
rect 23160 1730 23180 1750
rect 23215 1730 23235 1750
rect 23395 1730 23415 1750
rect 23450 1730 23470 1750
rect 23505 1730 23525 1750
rect 23615 1730 23635 1750
rect 23670 1730 23690 1750
rect 23725 1730 23745 1750
rect 23925 1730 23945 1750
rect 23980 1730 24000 1750
rect 24095 1730 24115 1750
rect 24150 1730 24170 1750
rect 24205 1730 24225 1750
rect 24275 1730 24295 1750
rect 24330 1730 24350 1750
rect 24385 1730 24405 1750
rect 24575 1730 24595 1750
rect 24630 1730 24650 1750
rect 24745 1730 24765 1750
rect 24800 1730 24820 1750
rect 24855 1730 24875 1750
rect 24925 1730 24945 1750
rect 24980 1730 25000 1750
rect 25035 1730 25055 1750
rect 25225 1730 25245 1750
rect 25280 1730 25300 1750
rect 25395 1730 25415 1750
rect 25450 1730 25470 1750
rect 25505 1730 25525 1750
rect 25575 1730 25595 1750
rect 25630 1730 25650 1750
rect 25685 1730 25705 1750
rect 25875 1730 25895 1750
rect 25930 1730 25950 1750
rect 26045 1730 26065 1750
rect 26100 1730 26120 1750
rect 26155 1730 26175 1750
rect 26225 1730 26245 1750
rect 26280 1730 26300 1750
rect 26335 1730 26355 1750
<< psubdiff >>
rect 22330 1545 22370 1560
rect 22840 1590 22880 1605
rect 22840 1570 22850 1590
rect 22870 1570 22880 1590
rect 22840 1555 22880 1570
rect 23565 1590 23605 1605
rect 23565 1570 23575 1590
rect 23595 1570 23605 1590
rect 23565 1555 23605 1570
rect 22330 1525 22340 1545
rect 22360 1525 22370 1545
rect 24460 1545 24500 1560
rect 22330 1510 22370 1525
rect 24460 1525 24470 1545
rect 24490 1525 24500 1545
rect 24460 1510 24500 1525
rect 25110 1545 25150 1560
rect 25110 1525 25120 1545
rect 25140 1525 25150 1545
rect 25110 1510 25150 1525
rect 25760 1545 25800 1560
rect 25760 1525 25770 1545
rect 25790 1525 25800 1545
rect 25760 1510 25800 1525
<< nsubdiff >>
rect 21370 1750 21410 1765
rect 21370 1730 21380 1750
rect 21400 1730 21410 1750
rect 21370 1715 21410 1730
rect 22575 1750 22615 1765
rect 22575 1730 22585 1750
rect 22605 1730 22615 1750
rect 22575 1715 22615 1730
rect 24010 1750 24050 1765
rect 24010 1730 24020 1750
rect 24040 1730 24050 1750
rect 24010 1715 24050 1730
rect 24660 1750 24700 1765
rect 24660 1730 24670 1750
rect 24690 1730 24700 1750
rect 24660 1715 24700 1730
rect 25310 1750 25350 1765
rect 25310 1730 25320 1750
rect 25340 1730 25350 1750
rect 25310 1715 25350 1730
rect 25960 1750 26000 1765
rect 25960 1730 25970 1750
rect 25990 1730 26000 1750
rect 25960 1715 26000 1730
<< psubdiffcont >>
rect 22850 1570 22870 1590
rect 23575 1570 23595 1590
rect 22340 1525 22360 1545
rect 24470 1525 24490 1545
rect 25120 1525 25140 1545
rect 25770 1525 25790 1545
<< nsubdiffcont >>
rect 21380 1730 21400 1750
rect 22585 1730 22605 1750
rect 24020 1730 24040 1750
rect 24670 1730 24690 1750
rect 25320 1730 25340 1750
rect 25970 1730 25990 1750
<< poly >>
rect 21490 1810 21540 1820
rect 22050 1810 22095 1820
rect 21490 1790 21500 1810
rect 21520 1790 21540 1810
rect 21490 1780 21540 1790
rect 21645 1800 21685 1810
rect 21645 1780 21655 1800
rect 21675 1780 21685 1800
rect 22050 1790 22060 1810
rect 22080 1790 22095 1810
rect 22050 1780 22095 1790
rect 22120 1810 22150 1820
rect 22120 1790 22125 1810
rect 22145 1790 22150 1810
rect 22120 1780 22150 1790
rect 22700 1810 22745 1820
rect 22700 1790 22710 1810
rect 22730 1790 22745 1810
rect 22700 1780 22745 1790
rect 23580 1815 23620 1820
rect 23580 1795 23590 1815
rect 23610 1800 23620 1815
rect 24830 1810 24885 1820
rect 23610 1795 23660 1800
rect 23580 1785 23660 1795
rect 24830 1790 24855 1810
rect 24875 1790 24885 1810
rect 25480 1810 25535 1820
rect 25480 1790 25505 1810
rect 25525 1790 25535 1810
rect 26130 1810 26185 1820
rect 26130 1790 26155 1810
rect 26175 1790 26185 1810
rect 21315 1765 21330 1780
rect 21525 1765 21540 1780
rect 21580 1765 21595 1780
rect 21645 1770 21685 1780
rect 21150 1750 21190 1760
rect 21150 1730 21160 1750
rect 21180 1730 21190 1750
rect 21150 1720 21190 1730
rect 21225 1650 21265 1660
rect 21225 1630 21235 1650
rect 21255 1630 21265 1650
rect 21315 1630 21330 1715
rect 21525 1700 21540 1715
rect 21580 1685 21595 1715
rect 21645 1685 21660 1770
rect 21860 1765 21875 1780
rect 21915 1765 21930 1780
rect 22080 1765 22095 1780
rect 22135 1765 22150 1780
rect 22190 1765 22205 1780
rect 22520 1765 22535 1780
rect 22730 1765 22745 1780
rect 22785 1765 22800 1780
rect 22955 1765 22970 1780
rect 23010 1765 23025 1780
rect 23135 1765 23150 1780
rect 23190 1765 23205 1780
rect 23425 1765 23440 1780
rect 23480 1765 23495 1780
rect 23645 1765 23660 1785
rect 23700 1765 23715 1780
rect 23955 1765 23970 1780
rect 24125 1765 24140 1780
rect 24180 1765 24195 1780
rect 24305 1775 24375 1790
rect 24830 1780 24885 1790
rect 24305 1765 24320 1775
rect 24360 1765 24375 1775
rect 24605 1765 24620 1780
rect 24775 1765 24790 1780
rect 24830 1765 24845 1780
rect 24955 1775 25025 1790
rect 25480 1780 25535 1790
rect 24955 1765 24970 1775
rect 25010 1765 25025 1775
rect 25255 1765 25270 1780
rect 25425 1765 25440 1780
rect 25480 1765 25495 1780
rect 25605 1775 25675 1790
rect 26130 1780 26185 1790
rect 25605 1765 25620 1775
rect 25660 1765 25675 1775
rect 25905 1765 25920 1780
rect 26075 1765 26090 1780
rect 26130 1765 26145 1780
rect 26255 1775 26325 1790
rect 26255 1765 26270 1775
rect 26310 1765 26325 1775
rect 21580 1670 21660 1685
rect 21785 1690 21825 1700
rect 21785 1675 21795 1690
rect 21515 1650 21555 1660
rect 21515 1630 21525 1650
rect 21545 1630 21555 1650
rect 21225 1620 21265 1630
rect 21290 1620 21555 1630
rect 21235 1605 21250 1620
rect 21290 1615 21540 1620
rect 21290 1605 21305 1615
rect 21345 1605 21360 1615
rect 21400 1605 21415 1615
rect 21525 1605 21540 1615
rect 21580 1605 21595 1670
rect 21235 1540 21250 1555
rect 21290 1540 21305 1555
rect 21345 1540 21360 1555
rect 21400 1540 21415 1555
rect 21525 1540 21540 1555
rect 21580 1540 21595 1555
rect 21645 1550 21660 1670
rect 21750 1670 21795 1675
rect 21815 1670 21825 1690
rect 21750 1660 21825 1670
rect 21685 1650 21725 1660
rect 21685 1630 21695 1650
rect 21715 1630 21725 1650
rect 21685 1620 21725 1630
rect 21750 1605 21765 1660
rect 21860 1635 21875 1715
rect 21915 1700 21930 1715
rect 21985 1710 22025 1720
rect 21985 1700 21995 1710
rect 21915 1690 21995 1700
rect 22015 1690 22025 1710
rect 21915 1685 22025 1690
rect 21985 1680 22025 1685
rect 21975 1650 22015 1655
rect 21975 1635 21985 1650
rect 21805 1630 21985 1635
rect 22005 1630 22015 1650
rect 21805 1620 22015 1630
rect 21805 1605 21820 1620
rect 21860 1605 21875 1620
rect 21915 1605 21930 1620
rect 22080 1605 22095 1715
rect 22135 1605 22150 1715
rect 22190 1605 22205 1715
rect 22520 1695 22535 1715
rect 22730 1700 22745 1715
rect 22355 1680 22535 1695
rect 22235 1650 22275 1655
rect 22235 1630 22245 1650
rect 22265 1635 22275 1650
rect 22355 1635 22370 1680
rect 22265 1630 22370 1635
rect 22235 1620 22370 1630
rect 22430 1650 22470 1655
rect 22430 1630 22440 1650
rect 22460 1630 22470 1650
rect 22520 1630 22535 1680
rect 22785 1695 22800 1715
rect 22855 1710 22895 1720
rect 22855 1695 22865 1710
rect 22785 1690 22865 1695
rect 22885 1690 22895 1710
rect 22955 1705 22970 1715
rect 23010 1705 23025 1715
rect 22955 1690 23025 1705
rect 23135 1705 23150 1715
rect 23190 1705 23205 1715
rect 23135 1690 23205 1705
rect 22785 1680 22895 1690
rect 22720 1650 22760 1660
rect 22720 1630 22730 1650
rect 22750 1630 22760 1650
rect 22430 1620 22470 1630
rect 22495 1620 22760 1630
rect 22245 1605 22260 1620
rect 22440 1605 22455 1620
rect 22495 1615 22745 1620
rect 22495 1605 22510 1615
rect 22550 1605 22565 1615
rect 22605 1605 22620 1615
rect 22730 1605 22745 1615
rect 22785 1605 22800 1680
rect 22825 1650 22865 1655
rect 22945 1650 22985 1660
rect 22825 1630 22835 1650
rect 22855 1635 22955 1650
rect 22855 1630 22865 1635
rect 22825 1620 22865 1630
rect 22945 1630 22955 1635
rect 22975 1630 22985 1650
rect 22945 1620 22985 1630
rect 23010 1605 23025 1690
rect 23190 1670 23205 1690
rect 23350 1690 23390 1700
rect 23250 1675 23290 1685
rect 23350 1675 23360 1690
rect 23250 1670 23260 1675
rect 23115 1655 23155 1665
rect 23115 1635 23125 1655
rect 23145 1635 23155 1655
rect 23115 1625 23155 1635
rect 23190 1655 23260 1670
rect 23280 1655 23290 1675
rect 23190 1605 23205 1655
rect 23250 1645 23290 1655
rect 23315 1670 23360 1675
rect 23380 1670 23390 1690
rect 23315 1660 23390 1670
rect 23315 1605 23330 1660
rect 23425 1635 23440 1715
rect 23480 1700 23495 1715
rect 23550 1710 23590 1720
rect 23845 1750 23885 1760
rect 23845 1735 23855 1750
rect 23765 1730 23855 1735
rect 23875 1730 23885 1750
rect 23765 1720 23885 1730
rect 23550 1700 23560 1710
rect 23480 1690 23560 1700
rect 23580 1690 23590 1710
rect 23480 1685 23590 1690
rect 23550 1680 23590 1685
rect 23565 1650 23605 1655
rect 23565 1635 23575 1650
rect 23370 1630 23575 1635
rect 23595 1630 23605 1650
rect 23370 1620 23605 1630
rect 23370 1605 23385 1620
rect 23425 1605 23440 1620
rect 23480 1605 23495 1620
rect 23645 1605 23660 1715
rect 23700 1695 23715 1715
rect 23765 1695 23780 1720
rect 23955 1695 23970 1715
rect 24125 1700 24140 1715
rect 24180 1705 24195 1715
rect 23700 1680 23780 1695
rect 23835 1680 23990 1695
rect 23700 1605 23715 1680
rect 23745 1650 23785 1655
rect 23745 1630 23755 1650
rect 23775 1635 23785 1650
rect 23835 1635 23850 1680
rect 23775 1630 23850 1635
rect 23745 1620 23850 1630
rect 23910 1650 23950 1655
rect 23910 1630 23920 1650
rect 23940 1630 23950 1650
rect 23910 1620 23950 1630
rect 23975 1630 23990 1680
rect 24115 1690 24155 1700
rect 24180 1690 24280 1705
rect 24305 1700 24320 1715
rect 24115 1670 24125 1690
rect 24145 1670 24155 1690
rect 24115 1660 24155 1670
rect 24265 1675 24280 1690
rect 24265 1660 24320 1675
rect 24200 1650 24240 1660
rect 24200 1630 24210 1650
rect 24230 1630 24240 1650
rect 23755 1605 23770 1620
rect 23920 1605 23935 1620
rect 23975 1615 24265 1630
rect 23975 1605 23990 1615
rect 24030 1605 24045 1615
rect 24085 1605 24100 1615
rect 24250 1605 24265 1615
rect 24305 1605 24320 1660
rect 24360 1660 24375 1715
rect 24605 1700 24620 1715
rect 24775 1700 24790 1715
rect 24605 1685 24640 1700
rect 24435 1660 24475 1670
rect 24360 1645 24445 1660
rect 24360 1605 24375 1645
rect 24435 1640 24445 1645
rect 24465 1640 24475 1660
rect 24435 1630 24475 1640
rect 24560 1605 24600 1615
rect 21645 1540 21685 1550
rect 21750 1540 21765 1555
rect 21805 1540 21820 1555
rect 21860 1540 21875 1555
rect 21915 1540 21930 1555
rect 22080 1540 22095 1555
rect 22135 1540 22150 1555
rect 22190 1540 22205 1555
rect 22245 1540 22260 1555
rect 24560 1585 24570 1605
rect 24590 1585 24600 1605
rect 24560 1575 24600 1585
rect 24625 1585 24640 1685
rect 24765 1690 24805 1700
rect 24765 1670 24775 1690
rect 24795 1670 24805 1690
rect 24765 1660 24805 1670
rect 24830 1660 24845 1715
rect 24955 1700 24970 1715
rect 25010 1660 25025 1715
rect 25255 1700 25270 1715
rect 25425 1700 25440 1715
rect 25255 1685 25290 1700
rect 25085 1660 25125 1670
rect 24830 1645 24970 1660
rect 24850 1605 24890 1615
rect 24850 1585 24860 1605
rect 24880 1585 24890 1605
rect 24570 1560 24585 1575
rect 24625 1570 24915 1585
rect 24625 1560 24640 1570
rect 24680 1560 24695 1570
rect 24735 1560 24750 1570
rect 24900 1560 24915 1570
rect 24955 1560 24970 1645
rect 25010 1645 25095 1660
rect 25010 1560 25025 1645
rect 25085 1640 25095 1645
rect 25115 1640 25125 1660
rect 25085 1630 25125 1640
rect 25210 1605 25250 1615
rect 25210 1585 25220 1605
rect 25240 1585 25250 1605
rect 25210 1575 25250 1585
rect 25275 1585 25290 1685
rect 25415 1690 25455 1700
rect 25415 1670 25425 1690
rect 25445 1670 25455 1690
rect 25415 1660 25455 1670
rect 25480 1660 25495 1715
rect 25605 1700 25620 1715
rect 25660 1660 25675 1715
rect 25905 1700 25920 1715
rect 26075 1700 26090 1715
rect 25905 1685 25940 1700
rect 25735 1660 25775 1670
rect 25480 1645 25620 1660
rect 25500 1605 25540 1615
rect 25500 1585 25510 1605
rect 25530 1585 25540 1605
rect 25220 1560 25235 1575
rect 25275 1570 25565 1585
rect 25275 1560 25290 1570
rect 25330 1560 25345 1570
rect 25385 1560 25400 1570
rect 25550 1560 25565 1570
rect 25605 1560 25620 1645
rect 25660 1645 25745 1660
rect 25660 1560 25675 1645
rect 25735 1640 25745 1645
rect 25765 1640 25775 1660
rect 25735 1630 25775 1640
rect 25860 1605 25900 1615
rect 25860 1585 25870 1605
rect 25890 1585 25900 1605
rect 25860 1575 25900 1585
rect 25925 1585 25940 1685
rect 26065 1690 26105 1700
rect 26065 1670 26075 1690
rect 26095 1670 26105 1690
rect 26065 1660 26105 1670
rect 26130 1660 26145 1715
rect 26255 1700 26270 1715
rect 26310 1660 26325 1715
rect 26376 1661 26405 1670
rect 26376 1660 26382 1661
rect 26130 1645 26270 1660
rect 26150 1605 26190 1615
rect 26150 1585 26160 1605
rect 26180 1585 26190 1605
rect 25870 1560 25885 1575
rect 25925 1570 26215 1585
rect 25925 1560 25940 1570
rect 25980 1560 25995 1570
rect 26035 1560 26050 1570
rect 26200 1560 26215 1570
rect 26255 1560 26270 1645
rect 26310 1645 26382 1660
rect 26310 1560 26325 1645
rect 26376 1644 26382 1645
rect 26399 1644 26405 1661
rect 26376 1630 26405 1644
rect 21150 1530 21190 1540
rect 21150 1510 21160 1530
rect 21180 1510 21190 1530
rect 21645 1520 21655 1540
rect 21675 1520 21685 1540
rect 21645 1510 21685 1520
rect 22180 1535 22220 1540
rect 22180 1515 22190 1535
rect 22210 1515 22220 1535
rect 21150 1500 21190 1510
rect 22180 1505 22220 1515
rect 22440 1540 22455 1555
rect 22495 1540 22510 1555
rect 22550 1540 22565 1555
rect 22605 1540 22620 1555
rect 22730 1540 22745 1555
rect 22785 1540 22800 1555
rect 23010 1540 23025 1555
rect 23190 1540 23205 1555
rect 23315 1540 23330 1555
rect 23370 1540 23385 1555
rect 23425 1540 23440 1555
rect 23480 1540 23495 1555
rect 23645 1540 23660 1555
rect 23700 1540 23715 1555
rect 23755 1540 23770 1555
rect 23920 1540 23935 1555
rect 23975 1540 23990 1555
rect 24030 1540 24045 1555
rect 24085 1540 24100 1555
rect 24250 1540 24265 1555
rect 24305 1540 24320 1555
rect 24360 1540 24375 1555
rect 22980 1535 23025 1540
rect 22980 1515 22990 1535
rect 23010 1515 23025 1535
rect 22980 1505 23025 1515
rect 24287 1530 24320 1540
rect 24287 1510 24292 1530
rect 24312 1510 24320 1530
rect 24287 1500 24320 1510
rect 24570 1495 24585 1510
rect 24625 1495 24640 1510
rect 24680 1495 24695 1510
rect 24735 1495 24750 1510
rect 24900 1495 24915 1510
rect 24955 1495 24970 1510
rect 25010 1495 25025 1510
rect 25220 1495 25235 1510
rect 25275 1495 25290 1510
rect 25330 1495 25345 1510
rect 25385 1495 25400 1510
rect 25550 1495 25565 1510
rect 25605 1495 25620 1510
rect 25660 1495 25675 1510
rect 25870 1495 25885 1510
rect 25925 1495 25940 1510
rect 25980 1495 25995 1510
rect 26035 1495 26050 1510
rect 26200 1495 26215 1510
rect 26255 1495 26270 1510
rect 26310 1495 26325 1510
<< polycont >>
rect 21500 1790 21520 1810
rect 21655 1780 21675 1800
rect 22060 1790 22080 1810
rect 22125 1790 22145 1810
rect 22710 1790 22730 1810
rect 23590 1795 23610 1815
rect 24855 1790 24875 1810
rect 25505 1790 25525 1810
rect 26155 1790 26175 1810
rect 21160 1730 21180 1750
rect 21235 1630 21255 1650
rect 21525 1630 21545 1650
rect 21795 1670 21815 1690
rect 21695 1630 21715 1650
rect 21995 1690 22015 1710
rect 21985 1630 22005 1650
rect 22245 1630 22265 1650
rect 22440 1630 22460 1650
rect 22865 1690 22885 1710
rect 22730 1630 22750 1650
rect 22835 1630 22855 1650
rect 22955 1630 22975 1650
rect 23125 1635 23145 1655
rect 23260 1655 23280 1675
rect 23360 1670 23380 1690
rect 23855 1730 23875 1750
rect 23560 1690 23580 1710
rect 23575 1630 23595 1650
rect 23755 1630 23775 1650
rect 23920 1630 23940 1650
rect 24125 1670 24145 1690
rect 24210 1630 24230 1650
rect 24445 1640 24465 1660
rect 24570 1585 24590 1605
rect 24775 1670 24795 1690
rect 24860 1585 24880 1605
rect 25095 1640 25115 1660
rect 25220 1585 25240 1605
rect 25425 1670 25445 1690
rect 25510 1585 25530 1605
rect 25745 1640 25765 1660
rect 25870 1585 25890 1605
rect 26075 1670 26095 1690
rect 26160 1585 26180 1605
rect 26382 1644 26399 1661
rect 21160 1510 21180 1530
rect 21655 1520 21675 1540
rect 22190 1515 22210 1535
rect 22990 1515 23010 1535
rect 24292 1510 24312 1530
<< locali >>
rect 21330 1865 21370 1875
rect 21330 1845 21340 1865
rect 21360 1845 21370 1865
rect 21330 1835 21370 1845
rect 21540 1865 21580 1875
rect 21540 1845 21550 1865
rect 21570 1845 21580 1865
rect 21540 1835 21580 1845
rect 21875 1865 21915 1875
rect 21875 1845 21885 1865
rect 21905 1845 21915 1865
rect 21875 1835 21915 1845
rect 22160 1865 22200 1875
rect 22160 1845 22170 1865
rect 22190 1845 22200 1865
rect 22160 1835 22200 1845
rect 22535 1865 22575 1875
rect 22535 1845 22545 1865
rect 22565 1845 22575 1865
rect 22535 1835 22575 1845
rect 22750 1865 22790 1875
rect 22750 1845 22760 1865
rect 22780 1845 22790 1865
rect 22750 1835 22790 1845
rect 22970 1865 23010 1875
rect 22970 1845 22980 1865
rect 23000 1845 23010 1865
rect 22970 1835 23010 1845
rect 23095 1865 23135 1875
rect 23095 1845 23105 1865
rect 23125 1845 23135 1865
rect 23095 1835 23135 1845
rect 23205 1865 23245 1875
rect 23205 1845 23215 1865
rect 23235 1845 23245 1865
rect 23205 1835 23245 1845
rect 23440 1865 23480 1875
rect 23440 1845 23450 1865
rect 23470 1845 23480 1865
rect 23440 1835 23480 1845
rect 23660 1865 23700 1875
rect 23660 1845 23670 1865
rect 23690 1845 23700 1865
rect 23660 1835 23700 1845
rect 23970 1865 24010 1875
rect 23970 1845 23980 1865
rect 24000 1845 24010 1865
rect 23970 1835 24010 1845
rect 24140 1865 24180 1875
rect 24140 1845 24150 1865
rect 24170 1845 24180 1865
rect 24140 1835 24180 1845
rect 24320 1865 24360 1875
rect 24320 1845 24330 1865
rect 24350 1845 24360 1865
rect 24320 1835 24360 1845
rect 24620 1865 24660 1875
rect 24620 1845 24630 1865
rect 24650 1845 24660 1865
rect 24620 1835 24660 1845
rect 24790 1865 24830 1875
rect 24790 1845 24800 1865
rect 24820 1845 24830 1865
rect 24790 1835 24830 1845
rect 24970 1865 25010 1875
rect 24970 1845 24980 1865
rect 25000 1845 25010 1865
rect 24970 1835 25010 1845
rect 25270 1865 25310 1875
rect 25270 1845 25280 1865
rect 25300 1845 25310 1865
rect 25270 1835 25310 1845
rect 25440 1865 25480 1875
rect 25440 1845 25450 1865
rect 25470 1845 25480 1865
rect 25440 1835 25480 1845
rect 25620 1865 25660 1875
rect 25620 1845 25630 1865
rect 25650 1845 25660 1865
rect 25620 1835 25660 1845
rect 25920 1865 25960 1875
rect 25920 1845 25930 1865
rect 25950 1845 25960 1865
rect 25920 1835 25960 1845
rect 26090 1865 26130 1875
rect 26090 1845 26100 1865
rect 26120 1845 26130 1865
rect 26090 1835 26130 1845
rect 26270 1865 26310 1875
rect 26270 1845 26280 1865
rect 26300 1845 26310 1865
rect 26270 1835 26310 1845
rect 21340 1760 21360 1835
rect 21490 1810 21530 1820
rect 21490 1790 21500 1810
rect 21520 1790 21530 1810
rect 21490 1780 21530 1790
rect 21550 1760 21570 1835
rect 21590 1810 21625 1820
rect 21590 1790 21595 1810
rect 21615 1790 21625 1810
rect 21590 1780 21625 1790
rect 21605 1760 21625 1780
rect 21645 1800 21685 1810
rect 21645 1780 21655 1800
rect 21675 1780 21685 1800
rect 21645 1770 21685 1780
rect 21885 1760 21905 1835
rect 22050 1810 22090 1820
rect 22050 1790 22060 1810
rect 22080 1790 22090 1810
rect 22050 1780 22090 1790
rect 22120 1810 22150 1820
rect 22120 1790 22125 1810
rect 22145 1790 22150 1810
rect 22120 1780 22150 1790
rect 22170 1760 22190 1835
rect 22545 1760 22565 1835
rect 22700 1810 22740 1820
rect 22700 1790 22710 1810
rect 22730 1790 22740 1810
rect 22700 1780 22740 1790
rect 22760 1760 22780 1835
rect 22810 1810 22850 1820
rect 22810 1790 22820 1810
rect 22840 1790 22850 1810
rect 22810 1780 22850 1790
rect 22810 1760 22830 1780
rect 22980 1760 23000 1835
rect 23105 1760 23125 1835
rect 23215 1760 23235 1835
rect 23375 1815 23415 1820
rect 23375 1795 23385 1815
rect 23405 1795 23415 1815
rect 23375 1785 23415 1795
rect 23395 1760 23415 1785
rect 23450 1760 23470 1835
rect 23580 1815 23620 1820
rect 23580 1795 23590 1815
rect 23610 1795 23620 1815
rect 23580 1785 23620 1795
rect 23670 1760 23690 1835
rect 23980 1760 24000 1835
rect 24150 1760 24170 1835
rect 24330 1760 24350 1835
rect 24555 1810 24595 1820
rect 24555 1790 24565 1810
rect 24585 1790 24595 1810
rect 24555 1780 24595 1790
rect 24575 1760 24595 1780
rect 24630 1760 24650 1835
rect 24800 1760 24820 1835
rect 24845 1810 24885 1820
rect 24845 1790 24855 1810
rect 24875 1790 24885 1810
rect 24845 1780 24885 1790
rect 24980 1760 25000 1835
rect 25205 1810 25245 1820
rect 25205 1790 25215 1810
rect 25235 1790 25245 1810
rect 25205 1780 25245 1790
rect 25225 1760 25245 1780
rect 25280 1760 25300 1835
rect 25450 1760 25470 1835
rect 25495 1810 25535 1820
rect 25495 1790 25505 1810
rect 25525 1790 25535 1810
rect 25495 1780 25535 1790
rect 25630 1760 25650 1835
rect 25855 1810 25895 1820
rect 25855 1790 25865 1810
rect 25885 1790 25895 1810
rect 25855 1780 25895 1790
rect 25875 1760 25895 1780
rect 25930 1760 25950 1835
rect 26100 1760 26120 1835
rect 26145 1810 26185 1820
rect 26145 1790 26155 1810
rect 26175 1790 26185 1810
rect 26145 1780 26185 1790
rect 26280 1760 26300 1835
rect 21150 1750 21190 1760
rect 21280 1750 21310 1760
rect 21150 1730 21160 1750
rect 21180 1730 21285 1750
rect 21305 1730 21310 1750
rect 21150 1720 21190 1730
rect 21280 1720 21310 1730
rect 21335 1750 21405 1760
rect 21490 1750 21520 1760
rect 21335 1730 21340 1750
rect 21360 1730 21380 1750
rect 21400 1730 21405 1750
rect 21335 1720 21405 1730
rect 21425 1730 21495 1750
rect 21515 1730 21520 1750
rect 21160 1675 21180 1720
rect 21120 1665 21180 1675
rect 21120 1645 21130 1665
rect 21150 1645 21180 1665
rect 21120 1635 21180 1645
rect 21160 1600 21180 1635
rect 21225 1650 21265 1660
rect 21225 1630 21235 1650
rect 21255 1640 21265 1650
rect 21425 1640 21445 1730
rect 21490 1720 21520 1730
rect 21545 1750 21575 1760
rect 21545 1730 21550 1750
rect 21570 1730 21575 1750
rect 21545 1720 21575 1730
rect 21600 1750 21630 1760
rect 21825 1750 21855 1760
rect 21600 1730 21605 1750
rect 21625 1730 21630 1750
rect 21600 1720 21630 1730
rect 21715 1730 21830 1750
rect 21850 1730 21855 1750
rect 21605 1700 21625 1720
rect 21255 1630 21445 1640
rect 21225 1620 21445 1630
rect 21315 1600 21335 1620
rect 21425 1600 21445 1620
rect 21470 1680 21625 1700
rect 21470 1600 21490 1680
rect 21715 1660 21735 1730
rect 21825 1720 21855 1730
rect 21880 1750 21910 1760
rect 21880 1730 21885 1750
rect 21905 1730 21910 1750
rect 21880 1720 21910 1730
rect 21935 1750 21965 1760
rect 21935 1730 21940 1750
rect 21960 1730 21965 1750
rect 21935 1720 21965 1730
rect 22045 1750 22075 1760
rect 22045 1730 22050 1750
rect 22070 1730 22075 1750
rect 22045 1720 22075 1730
rect 22100 1750 22130 1760
rect 22100 1730 22105 1750
rect 22125 1730 22130 1750
rect 22100 1720 22130 1730
rect 22155 1750 22190 1760
rect 22155 1730 22160 1750
rect 22180 1730 22190 1750
rect 22155 1720 22190 1730
rect 22210 1750 22240 1760
rect 22210 1730 22215 1750
rect 22235 1730 22240 1750
rect 22210 1720 22240 1730
rect 22365 1750 22405 1760
rect 22485 1750 22515 1760
rect 22365 1730 22375 1750
rect 22395 1730 22490 1750
rect 22510 1730 22515 1750
rect 22365 1720 22405 1730
rect 22485 1720 22515 1730
rect 22540 1750 22610 1760
rect 22695 1750 22725 1760
rect 22540 1730 22545 1750
rect 22565 1730 22585 1750
rect 22605 1730 22610 1750
rect 22540 1720 22610 1730
rect 22630 1730 22700 1750
rect 22720 1730 22725 1750
rect 21785 1690 21825 1700
rect 21785 1670 21795 1690
rect 21815 1670 21825 1690
rect 21785 1660 21825 1670
rect 21515 1650 21555 1660
rect 21685 1650 21735 1660
rect 21515 1630 21525 1650
rect 21545 1630 21695 1650
rect 21715 1630 21735 1650
rect 21515 1620 21555 1630
rect 21685 1620 21735 1630
rect 21805 1640 21825 1660
rect 21935 1640 21955 1720
rect 21985 1710 22025 1720
rect 21985 1690 21995 1710
rect 22015 1700 22025 1710
rect 22050 1700 22070 1720
rect 22215 1700 22235 1720
rect 22015 1690 22315 1700
rect 21985 1680 22315 1690
rect 21805 1620 21955 1640
rect 21975 1650 22015 1655
rect 21975 1630 21985 1650
rect 22005 1630 22015 1650
rect 22235 1650 22275 1655
rect 21975 1620 22015 1630
rect 22050 1620 22180 1640
rect 22235 1630 22245 1650
rect 22265 1630 22275 1650
rect 22235 1620 22275 1630
rect 21715 1600 21735 1620
rect 21825 1600 21845 1620
rect 21935 1600 21955 1620
rect 22050 1600 22070 1620
rect 22160 1600 22180 1620
rect 22295 1600 22315 1680
rect 21160 1590 21230 1600
rect 21160 1570 21205 1590
rect 21225 1570 21230 1590
rect 21160 1560 21230 1570
rect 21255 1590 21285 1600
rect 21255 1570 21260 1590
rect 21280 1570 21285 1590
rect 21255 1560 21285 1570
rect 21310 1590 21340 1600
rect 21310 1570 21315 1590
rect 21335 1570 21340 1590
rect 21310 1560 21340 1570
rect 21365 1590 21395 1600
rect 21365 1570 21370 1590
rect 21390 1570 21395 1590
rect 21365 1560 21395 1570
rect 21420 1590 21450 1600
rect 21420 1570 21425 1590
rect 21445 1570 21450 1590
rect 21470 1590 21520 1600
rect 21470 1570 21495 1590
rect 21515 1570 21520 1590
rect 21420 1560 21450 1570
rect 21490 1560 21520 1570
rect 21545 1590 21575 1600
rect 21545 1570 21550 1590
rect 21570 1570 21575 1590
rect 21545 1560 21575 1570
rect 21600 1590 21630 1600
rect 21600 1570 21605 1590
rect 21625 1570 21630 1590
rect 21600 1560 21630 1570
rect 21715 1590 21745 1600
rect 21715 1570 21720 1590
rect 21740 1570 21745 1590
rect 21715 1560 21745 1570
rect 21770 1590 21800 1600
rect 21770 1570 21775 1590
rect 21795 1570 21800 1590
rect 21770 1560 21800 1570
rect 21825 1590 21855 1600
rect 21825 1570 21830 1590
rect 21850 1570 21855 1590
rect 21825 1560 21855 1570
rect 21880 1590 21910 1600
rect 21880 1570 21885 1590
rect 21905 1570 21910 1590
rect 21880 1560 21910 1570
rect 21935 1590 21965 1600
rect 21935 1570 21940 1590
rect 21960 1570 21965 1590
rect 21935 1560 21965 1570
rect 22045 1590 22075 1600
rect 22045 1570 22050 1590
rect 22070 1570 22075 1590
rect 22045 1560 22075 1570
rect 22100 1590 22130 1600
rect 22100 1570 22105 1590
rect 22125 1570 22130 1590
rect 22100 1560 22130 1570
rect 22155 1590 22185 1600
rect 22155 1570 22160 1590
rect 22180 1570 22185 1590
rect 22155 1560 22185 1570
rect 22210 1590 22240 1600
rect 22210 1570 22215 1590
rect 22235 1570 22240 1590
rect 22210 1560 22240 1570
rect 22265 1590 22315 1600
rect 22265 1570 22270 1590
rect 22290 1570 22315 1590
rect 22385 1600 22405 1720
rect 22430 1650 22470 1655
rect 22430 1630 22440 1650
rect 22460 1640 22470 1650
rect 22630 1640 22650 1730
rect 22695 1720 22725 1730
rect 22750 1750 22780 1760
rect 22750 1730 22755 1750
rect 22775 1730 22780 1750
rect 22750 1720 22780 1730
rect 22805 1750 22835 1760
rect 22805 1730 22810 1750
rect 22830 1730 22835 1750
rect 22805 1720 22835 1730
rect 22920 1750 22950 1760
rect 22920 1730 22925 1750
rect 22945 1730 22950 1750
rect 22920 1720 22950 1730
rect 22975 1750 23005 1760
rect 22975 1730 22980 1750
rect 23000 1730 23005 1750
rect 22975 1720 23005 1730
rect 23030 1750 23060 1760
rect 23030 1730 23035 1750
rect 23055 1730 23060 1750
rect 23030 1720 23060 1730
rect 23100 1750 23130 1760
rect 23100 1730 23105 1750
rect 23125 1730 23130 1750
rect 23100 1720 23130 1730
rect 23155 1750 23185 1760
rect 23155 1730 23160 1750
rect 23180 1730 23185 1750
rect 23155 1720 23185 1730
rect 23210 1750 23240 1760
rect 23390 1750 23420 1760
rect 23210 1730 23215 1750
rect 23235 1730 23240 1750
rect 23210 1720 23240 1730
rect 23280 1730 23395 1750
rect 23415 1730 23420 1750
rect 22810 1700 22830 1720
rect 22460 1630 22650 1640
rect 22430 1620 22650 1630
rect 22520 1600 22540 1620
rect 22630 1600 22650 1620
rect 22675 1680 22830 1700
rect 22855 1710 22895 1720
rect 22855 1690 22865 1710
rect 22885 1700 22895 1710
rect 22925 1700 22945 1720
rect 23035 1700 23055 1720
rect 22885 1690 23055 1700
rect 22855 1680 23055 1690
rect 22675 1600 22695 1680
rect 22720 1650 22760 1660
rect 22825 1650 22865 1655
rect 22720 1630 22730 1650
rect 22750 1630 22835 1650
rect 22855 1630 22865 1650
rect 22720 1620 22760 1630
rect 22825 1620 22865 1630
rect 22385 1590 22435 1600
rect 22385 1570 22410 1590
rect 22430 1570 22435 1590
rect 22265 1560 22295 1570
rect 22405 1560 22435 1570
rect 22460 1590 22490 1600
rect 22460 1570 22465 1590
rect 22485 1570 22490 1590
rect 22460 1560 22490 1570
rect 22515 1590 22545 1600
rect 22515 1570 22520 1590
rect 22540 1570 22545 1590
rect 22515 1560 22545 1570
rect 22570 1590 22600 1600
rect 22570 1570 22575 1590
rect 22595 1570 22600 1590
rect 22570 1560 22600 1570
rect 22625 1590 22655 1600
rect 22625 1570 22630 1590
rect 22650 1570 22655 1590
rect 22675 1590 22725 1600
rect 22675 1570 22700 1590
rect 22720 1570 22725 1590
rect 22625 1560 22655 1570
rect 22695 1560 22725 1570
rect 22750 1590 22780 1600
rect 22750 1570 22755 1590
rect 22775 1570 22780 1590
rect 22750 1560 22780 1570
rect 22805 1590 22875 1600
rect 22805 1570 22810 1590
rect 22830 1570 22850 1590
rect 22870 1570 22875 1590
rect 22895 1590 22915 1680
rect 23160 1665 23180 1720
rect 23280 1685 23300 1730
rect 23390 1720 23420 1730
rect 23445 1750 23475 1760
rect 23445 1730 23450 1750
rect 23470 1730 23475 1750
rect 23445 1720 23475 1730
rect 23500 1750 23530 1760
rect 23500 1730 23505 1750
rect 23525 1730 23530 1750
rect 23500 1720 23530 1730
rect 23610 1750 23640 1760
rect 23610 1730 23615 1750
rect 23635 1730 23640 1750
rect 23610 1720 23640 1730
rect 23665 1750 23695 1760
rect 23665 1730 23670 1750
rect 23690 1730 23695 1750
rect 23665 1720 23695 1730
rect 23720 1750 23750 1760
rect 23845 1750 23885 1760
rect 23920 1750 23950 1760
rect 23720 1730 23725 1750
rect 23745 1730 23825 1750
rect 23720 1720 23750 1730
rect 23115 1660 23180 1665
rect 22945 1655 23180 1660
rect 22945 1650 23125 1655
rect 22945 1630 22955 1650
rect 22975 1640 23125 1650
rect 22975 1630 22985 1640
rect 22945 1620 22985 1630
rect 23115 1635 23125 1640
rect 23145 1635 23180 1655
rect 23250 1675 23300 1685
rect 23250 1655 23260 1675
rect 23280 1655 23300 1675
rect 23350 1690 23390 1700
rect 23350 1670 23360 1690
rect 23380 1670 23390 1690
rect 23350 1660 23390 1670
rect 23250 1645 23300 1655
rect 23115 1625 23180 1635
rect 23160 1600 23180 1625
rect 23280 1600 23300 1645
rect 23370 1640 23390 1660
rect 23500 1640 23520 1720
rect 23550 1710 23590 1720
rect 23550 1690 23560 1710
rect 23580 1700 23590 1710
rect 23615 1700 23635 1720
rect 23725 1700 23745 1720
rect 23580 1690 23745 1700
rect 23550 1680 23745 1690
rect 23370 1620 23520 1640
rect 23565 1650 23605 1655
rect 23745 1650 23785 1655
rect 23565 1630 23575 1650
rect 23595 1630 23755 1650
rect 23775 1630 23785 1650
rect 23565 1620 23605 1630
rect 23745 1620 23785 1630
rect 23390 1600 23410 1620
rect 23500 1600 23520 1620
rect 23805 1600 23825 1730
rect 23845 1730 23855 1750
rect 23875 1730 23925 1750
rect 23945 1730 23950 1750
rect 23845 1720 23885 1730
rect 23920 1720 23950 1730
rect 23975 1750 24045 1760
rect 23975 1730 23980 1750
rect 24000 1730 24020 1750
rect 24040 1730 24045 1750
rect 23975 1720 24045 1730
rect 24075 1750 24120 1760
rect 24075 1730 24095 1750
rect 24115 1730 24120 1750
rect 24075 1720 24120 1730
rect 24145 1750 24175 1760
rect 24145 1730 24150 1750
rect 24170 1730 24175 1750
rect 24145 1720 24175 1730
rect 24200 1750 24230 1760
rect 24200 1730 24205 1750
rect 24225 1730 24230 1750
rect 24200 1720 24230 1730
rect 24270 1750 24300 1760
rect 24270 1730 24275 1750
rect 24295 1730 24300 1750
rect 24270 1720 24300 1730
rect 24325 1750 24355 1760
rect 24325 1730 24330 1750
rect 24350 1730 24355 1750
rect 24325 1720 24355 1730
rect 24380 1750 24410 1760
rect 24570 1750 24600 1760
rect 24380 1730 24385 1750
rect 24405 1730 24410 1750
rect 24380 1720 24410 1730
rect 24515 1730 24575 1750
rect 24595 1730 24600 1750
rect 22975 1590 23005 1600
rect 22895 1570 22980 1590
rect 23000 1570 23005 1590
rect 22805 1560 22875 1570
rect 22975 1560 23005 1570
rect 23030 1590 23060 1600
rect 23030 1570 23035 1590
rect 23055 1570 23060 1590
rect 23030 1560 23060 1570
rect 23155 1590 23185 1600
rect 23155 1570 23160 1590
rect 23180 1570 23185 1590
rect 23155 1560 23185 1570
rect 23210 1590 23240 1600
rect 23210 1570 23215 1590
rect 23235 1570 23240 1590
rect 23210 1560 23240 1570
rect 23280 1590 23310 1600
rect 23280 1570 23285 1590
rect 23305 1570 23310 1590
rect 23280 1560 23310 1570
rect 23335 1590 23365 1600
rect 23335 1570 23340 1590
rect 23360 1570 23365 1590
rect 23335 1560 23365 1570
rect 23390 1590 23420 1600
rect 23390 1570 23395 1590
rect 23415 1570 23420 1590
rect 23390 1560 23420 1570
rect 23445 1590 23475 1600
rect 23445 1570 23450 1590
rect 23470 1570 23475 1590
rect 23445 1560 23475 1570
rect 23500 1590 23530 1600
rect 23500 1570 23505 1590
rect 23525 1570 23530 1590
rect 23500 1560 23530 1570
rect 23570 1590 23640 1600
rect 23570 1570 23575 1590
rect 23595 1570 23615 1590
rect 23635 1570 23640 1590
rect 23570 1560 23640 1570
rect 23665 1590 23695 1600
rect 23665 1570 23670 1590
rect 23690 1570 23695 1590
rect 23665 1560 23695 1570
rect 23720 1590 23750 1600
rect 23720 1570 23725 1590
rect 23745 1570 23750 1590
rect 23720 1560 23750 1570
rect 23775 1590 23825 1600
rect 23775 1570 23780 1590
rect 23800 1570 23825 1590
rect 23865 1600 23885 1720
rect 23910 1650 23950 1655
rect 23910 1630 23920 1650
rect 23940 1640 23950 1650
rect 24075 1640 24095 1720
rect 24205 1700 24225 1720
rect 24115 1690 24225 1700
rect 24115 1670 24125 1690
rect 24145 1680 24225 1690
rect 24145 1670 24175 1680
rect 24115 1660 24175 1670
rect 23940 1630 24130 1640
rect 23910 1620 24130 1630
rect 24000 1600 24020 1620
rect 24110 1600 24130 1620
rect 24155 1600 24175 1660
rect 24200 1650 24240 1660
rect 24200 1630 24210 1650
rect 24230 1640 24240 1650
rect 24275 1640 24295 1720
rect 24385 1640 24405 1720
rect 24515 1670 24535 1730
rect 24570 1720 24600 1730
rect 24625 1750 24695 1760
rect 24625 1730 24630 1750
rect 24650 1730 24670 1750
rect 24690 1730 24695 1750
rect 24625 1720 24695 1730
rect 24725 1750 24770 1760
rect 24725 1730 24745 1750
rect 24765 1730 24770 1750
rect 24725 1720 24770 1730
rect 24795 1750 24825 1760
rect 24795 1730 24800 1750
rect 24820 1730 24825 1750
rect 24795 1720 24825 1730
rect 24850 1750 24880 1760
rect 24850 1730 24855 1750
rect 24875 1730 24880 1750
rect 24850 1720 24880 1730
rect 24920 1750 24950 1760
rect 24920 1730 24925 1750
rect 24945 1730 24950 1750
rect 24920 1720 24950 1730
rect 24975 1750 25005 1760
rect 24975 1730 24980 1750
rect 25000 1730 25005 1750
rect 24975 1720 25005 1730
rect 25030 1750 25060 1760
rect 25220 1750 25250 1760
rect 25030 1730 25035 1750
rect 25055 1730 25060 1750
rect 25030 1720 25060 1730
rect 25165 1730 25225 1750
rect 25245 1730 25250 1750
rect 24230 1630 24405 1640
rect 24435 1660 24535 1670
rect 24435 1640 24445 1660
rect 24465 1650 24535 1660
rect 24465 1640 24475 1650
rect 24435 1630 24475 1640
rect 24200 1620 24405 1630
rect 24385 1600 24405 1620
rect 23865 1590 23915 1600
rect 23865 1570 23890 1590
rect 23910 1570 23915 1590
rect 23775 1560 23805 1570
rect 23885 1560 23915 1570
rect 23940 1590 23970 1600
rect 23940 1570 23945 1590
rect 23965 1570 23970 1590
rect 23940 1560 23970 1570
rect 23995 1590 24025 1600
rect 23995 1570 24000 1590
rect 24020 1570 24025 1590
rect 23995 1560 24025 1570
rect 24050 1590 24080 1600
rect 24050 1570 24055 1590
rect 24075 1570 24080 1590
rect 24050 1560 24080 1570
rect 24105 1590 24135 1600
rect 24105 1570 24110 1590
rect 24130 1570 24135 1590
rect 24155 1590 24245 1600
rect 24155 1580 24220 1590
rect 24105 1560 24135 1570
rect 24215 1570 24220 1580
rect 24240 1570 24245 1590
rect 24215 1560 24245 1570
rect 24270 1590 24300 1600
rect 24270 1570 24275 1590
rect 24295 1570 24300 1590
rect 24270 1560 24300 1570
rect 24325 1590 24360 1600
rect 24325 1570 24330 1590
rect 24350 1570 24360 1590
rect 24325 1560 24360 1570
rect 24380 1590 24410 1600
rect 24380 1570 24385 1590
rect 24405 1570 24410 1590
rect 24380 1560 24410 1570
rect 21160 1540 21180 1560
rect 21150 1530 21190 1540
rect 21150 1510 21160 1530
rect 21180 1510 21190 1530
rect 21150 1500 21190 1510
rect 21260 1485 21280 1560
rect 21370 1485 21390 1560
rect 21605 1485 21625 1560
rect 21645 1540 21685 1550
rect 21720 1540 21740 1560
rect 21645 1520 21655 1540
rect 21675 1520 21685 1540
rect 21645 1510 21685 1520
rect 21710 1535 21750 1540
rect 21710 1515 21720 1535
rect 21740 1515 21750 1535
rect 21710 1505 21750 1515
rect 21775 1485 21795 1560
rect 21885 1485 21905 1560
rect 22105 1485 22125 1560
rect 22335 1545 22365 1555
rect 22180 1535 22220 1540
rect 22180 1515 22190 1535
rect 22210 1515 22220 1535
rect 22335 1525 22340 1545
rect 22360 1525 22365 1545
rect 22335 1515 22365 1525
rect 22180 1505 22220 1515
rect 22340 1485 22360 1515
rect 22465 1485 22485 1560
rect 22575 1485 22595 1560
rect 22810 1485 22830 1560
rect 22980 1535 23020 1540
rect 22980 1515 22990 1535
rect 23010 1515 23020 1535
rect 22980 1505 23020 1515
rect 23040 1485 23060 1560
rect 23215 1485 23235 1560
rect 23340 1485 23360 1560
rect 23450 1485 23470 1560
rect 23615 1485 23635 1560
rect 23945 1485 23965 1560
rect 24055 1485 24075 1560
rect 24287 1530 24320 1540
rect 24287 1510 24292 1530
rect 24312 1510 24320 1530
rect 24287 1500 24320 1510
rect 24340 1485 24360 1560
rect 24515 1555 24535 1650
rect 24560 1605 24600 1615
rect 24560 1585 24570 1605
rect 24590 1595 24600 1605
rect 24725 1595 24745 1720
rect 24855 1700 24875 1720
rect 24765 1690 24875 1700
rect 24765 1670 24775 1690
rect 24795 1680 24875 1690
rect 24795 1670 24825 1680
rect 24765 1660 24825 1670
rect 24590 1585 24780 1595
rect 24560 1575 24780 1585
rect 24650 1555 24670 1575
rect 24760 1555 24780 1575
rect 24805 1555 24825 1660
rect 24850 1605 24890 1615
rect 24850 1585 24860 1605
rect 24880 1595 24890 1605
rect 24925 1595 24945 1720
rect 25035 1595 25055 1720
rect 25165 1670 25185 1730
rect 25220 1720 25250 1730
rect 25275 1750 25345 1760
rect 25275 1730 25280 1750
rect 25300 1730 25320 1750
rect 25340 1730 25345 1750
rect 25275 1720 25345 1730
rect 25375 1750 25420 1760
rect 25375 1730 25395 1750
rect 25415 1730 25420 1750
rect 25375 1720 25420 1730
rect 25445 1750 25475 1760
rect 25445 1730 25450 1750
rect 25470 1730 25475 1750
rect 25445 1720 25475 1730
rect 25500 1750 25530 1760
rect 25500 1730 25505 1750
rect 25525 1730 25530 1750
rect 25500 1720 25530 1730
rect 25570 1750 25600 1760
rect 25570 1730 25575 1750
rect 25595 1730 25600 1750
rect 25570 1720 25600 1730
rect 25625 1750 25655 1760
rect 25625 1730 25630 1750
rect 25650 1730 25655 1750
rect 25625 1720 25655 1730
rect 25680 1750 25710 1760
rect 25870 1750 25900 1760
rect 25680 1730 25685 1750
rect 25705 1730 25710 1750
rect 25680 1720 25710 1730
rect 25815 1730 25875 1750
rect 25895 1730 25900 1750
rect 25085 1660 25185 1670
rect 25085 1640 25095 1660
rect 25115 1650 25185 1660
rect 25115 1640 25125 1650
rect 25085 1630 25125 1640
rect 24880 1585 25055 1595
rect 24850 1575 25055 1585
rect 25035 1555 25055 1575
rect 25165 1555 25185 1650
rect 25210 1605 25250 1615
rect 25210 1585 25220 1605
rect 25240 1595 25250 1605
rect 25375 1595 25395 1720
rect 25505 1700 25525 1720
rect 25415 1690 25525 1700
rect 25415 1670 25425 1690
rect 25445 1680 25525 1690
rect 25445 1670 25475 1680
rect 25415 1660 25475 1670
rect 25240 1585 25430 1595
rect 25210 1575 25430 1585
rect 25300 1555 25320 1575
rect 25410 1555 25430 1575
rect 25455 1555 25475 1660
rect 25500 1605 25540 1615
rect 25500 1585 25510 1605
rect 25530 1595 25540 1605
rect 25575 1595 25595 1720
rect 25685 1595 25705 1720
rect 25815 1670 25835 1730
rect 25870 1720 25900 1730
rect 25925 1750 25995 1760
rect 25925 1730 25930 1750
rect 25950 1730 25970 1750
rect 25990 1730 25995 1750
rect 25925 1720 25995 1730
rect 26025 1750 26070 1760
rect 26025 1730 26045 1750
rect 26065 1730 26070 1750
rect 26025 1720 26070 1730
rect 26095 1750 26125 1760
rect 26095 1730 26100 1750
rect 26120 1730 26125 1750
rect 26095 1720 26125 1730
rect 26150 1750 26180 1760
rect 26150 1730 26155 1750
rect 26175 1730 26180 1750
rect 26150 1720 26180 1730
rect 26220 1750 26250 1760
rect 26220 1730 26225 1750
rect 26245 1730 26250 1750
rect 26220 1720 26250 1730
rect 26275 1750 26305 1760
rect 26275 1730 26280 1750
rect 26300 1730 26305 1750
rect 26275 1720 26305 1730
rect 26330 1750 26360 1760
rect 26330 1730 26335 1750
rect 26355 1730 26360 1750
rect 26330 1720 26360 1730
rect 25735 1660 25835 1670
rect 25735 1640 25745 1660
rect 25765 1650 25835 1660
rect 25765 1640 25775 1650
rect 25735 1630 25775 1640
rect 25530 1585 25705 1595
rect 25500 1575 25705 1585
rect 25685 1555 25705 1575
rect 25815 1555 25835 1650
rect 25860 1605 25900 1615
rect 25860 1585 25870 1605
rect 25890 1595 25900 1605
rect 26025 1595 26045 1720
rect 26155 1700 26175 1720
rect 26065 1690 26175 1700
rect 26065 1670 26075 1690
rect 26095 1680 26175 1690
rect 26095 1670 26125 1680
rect 26065 1660 26125 1670
rect 25890 1585 26080 1595
rect 25860 1575 26080 1585
rect 25950 1555 25970 1575
rect 26060 1555 26080 1575
rect 26105 1555 26125 1660
rect 26150 1605 26190 1615
rect 26150 1585 26160 1605
rect 26180 1595 26190 1605
rect 26225 1595 26245 1720
rect 26335 1595 26355 1720
rect 26376 1661 26405 1670
rect 26376 1644 26382 1661
rect 26399 1644 26405 1661
rect 26376 1630 26405 1644
rect 26180 1585 26355 1595
rect 26150 1575 26355 1585
rect 26335 1555 26355 1575
rect 24465 1545 24495 1555
rect 24465 1525 24470 1545
rect 24490 1525 24495 1545
rect 24515 1545 24565 1555
rect 24515 1525 24540 1545
rect 24560 1525 24565 1545
rect 24465 1515 24495 1525
rect 24535 1515 24565 1525
rect 24590 1545 24620 1555
rect 24590 1525 24595 1545
rect 24615 1525 24620 1545
rect 24590 1515 24620 1525
rect 24645 1545 24675 1555
rect 24645 1525 24650 1545
rect 24670 1525 24675 1545
rect 24645 1515 24675 1525
rect 24700 1545 24730 1555
rect 24700 1525 24705 1545
rect 24725 1525 24730 1545
rect 24700 1515 24730 1525
rect 24755 1545 24785 1555
rect 24755 1525 24760 1545
rect 24780 1525 24785 1545
rect 24805 1545 24895 1555
rect 24805 1535 24870 1545
rect 24755 1515 24785 1525
rect 24865 1525 24870 1535
rect 24890 1525 24895 1545
rect 24865 1515 24895 1525
rect 24920 1545 24950 1555
rect 24920 1525 24925 1545
rect 24945 1525 24950 1545
rect 24920 1515 24950 1525
rect 24975 1545 25005 1555
rect 24975 1525 24980 1545
rect 25000 1525 25005 1545
rect 24975 1515 25005 1525
rect 25030 1545 25060 1555
rect 25030 1525 25035 1545
rect 25055 1525 25060 1545
rect 25030 1515 25060 1525
rect 25115 1545 25145 1555
rect 25115 1525 25120 1545
rect 25140 1525 25145 1545
rect 25165 1545 25215 1555
rect 25165 1525 25190 1545
rect 25210 1525 25215 1545
rect 25115 1515 25145 1525
rect 25185 1515 25215 1525
rect 25240 1545 25270 1555
rect 25240 1525 25245 1545
rect 25265 1525 25270 1545
rect 25240 1515 25270 1525
rect 25295 1545 25325 1555
rect 25295 1525 25300 1545
rect 25320 1525 25325 1545
rect 25295 1515 25325 1525
rect 25350 1545 25380 1555
rect 25350 1525 25355 1545
rect 25375 1525 25380 1545
rect 25350 1515 25380 1525
rect 25405 1545 25435 1555
rect 25405 1525 25410 1545
rect 25430 1525 25435 1545
rect 25455 1545 25545 1555
rect 25455 1535 25520 1545
rect 25405 1515 25435 1525
rect 25515 1525 25520 1535
rect 25540 1525 25545 1545
rect 25515 1515 25545 1525
rect 25570 1545 25600 1555
rect 25570 1525 25575 1545
rect 25595 1525 25600 1545
rect 25570 1515 25600 1525
rect 25625 1545 25655 1555
rect 25625 1525 25630 1545
rect 25650 1525 25655 1545
rect 25625 1515 25655 1525
rect 25680 1545 25710 1555
rect 25680 1525 25685 1545
rect 25705 1525 25710 1545
rect 25680 1515 25710 1525
rect 25765 1545 25795 1555
rect 25765 1525 25770 1545
rect 25790 1525 25795 1545
rect 25815 1545 25865 1555
rect 25815 1525 25840 1545
rect 25860 1525 25865 1545
rect 25765 1515 25795 1525
rect 25835 1515 25865 1525
rect 25890 1545 25920 1555
rect 25890 1525 25895 1545
rect 25915 1525 25920 1545
rect 25890 1515 25920 1525
rect 25945 1545 25975 1555
rect 25945 1525 25950 1545
rect 25970 1525 25975 1545
rect 25945 1515 25975 1525
rect 26000 1545 26030 1555
rect 26000 1525 26005 1545
rect 26025 1525 26030 1545
rect 26000 1515 26030 1525
rect 26055 1545 26085 1555
rect 26055 1525 26060 1545
rect 26080 1525 26085 1545
rect 26105 1545 26195 1555
rect 26105 1535 26170 1545
rect 26055 1515 26085 1525
rect 26165 1525 26170 1535
rect 26190 1525 26195 1545
rect 26165 1515 26195 1525
rect 26220 1545 26250 1555
rect 26220 1525 26225 1545
rect 26245 1525 26250 1545
rect 26220 1515 26250 1525
rect 26275 1545 26305 1555
rect 26275 1525 26280 1545
rect 26300 1525 26305 1545
rect 26275 1515 26305 1525
rect 26330 1545 26360 1555
rect 26330 1525 26335 1545
rect 26355 1525 26360 1545
rect 26330 1515 26360 1525
rect 24470 1485 24490 1515
rect 24595 1485 24615 1515
rect 24705 1485 24725 1515
rect 24980 1485 25000 1515
rect 25120 1485 25140 1515
rect 25245 1485 25265 1515
rect 25355 1485 25375 1515
rect 25630 1485 25650 1515
rect 25770 1485 25790 1515
rect 25895 1485 25915 1515
rect 26005 1485 26025 1515
rect 26280 1485 26300 1515
rect 21250 1475 21290 1485
rect 21250 1455 21260 1475
rect 21280 1455 21290 1475
rect 21250 1445 21290 1455
rect 21360 1475 21400 1485
rect 21360 1455 21370 1475
rect 21390 1455 21400 1475
rect 21360 1445 21400 1455
rect 21595 1475 21635 1485
rect 21595 1455 21605 1475
rect 21625 1455 21635 1475
rect 21595 1445 21635 1455
rect 21765 1475 21805 1485
rect 21765 1455 21775 1475
rect 21795 1455 21805 1475
rect 21765 1445 21805 1455
rect 21875 1475 21915 1485
rect 21875 1455 21885 1475
rect 21905 1455 21915 1475
rect 21875 1445 21915 1455
rect 22095 1475 22135 1485
rect 22095 1455 22105 1475
rect 22125 1455 22135 1475
rect 22095 1445 22135 1455
rect 22330 1475 22370 1485
rect 22330 1455 22340 1475
rect 22360 1455 22370 1475
rect 22330 1445 22370 1455
rect 22455 1475 22495 1485
rect 22455 1455 22465 1475
rect 22485 1455 22495 1475
rect 22455 1445 22495 1455
rect 22565 1475 22605 1485
rect 22565 1455 22575 1475
rect 22595 1455 22605 1475
rect 22565 1445 22605 1455
rect 22800 1475 22840 1485
rect 22800 1455 22810 1475
rect 22830 1455 22840 1475
rect 22800 1445 22840 1455
rect 23030 1475 23070 1485
rect 23030 1455 23040 1475
rect 23060 1455 23070 1475
rect 23030 1445 23070 1455
rect 23205 1475 23245 1485
rect 23205 1455 23215 1475
rect 23235 1455 23245 1475
rect 23205 1445 23245 1455
rect 23330 1475 23370 1485
rect 23330 1455 23340 1475
rect 23360 1455 23370 1475
rect 23330 1445 23370 1455
rect 23440 1475 23480 1485
rect 23440 1455 23450 1475
rect 23470 1455 23480 1475
rect 23440 1445 23480 1455
rect 23605 1475 23645 1485
rect 23605 1455 23615 1475
rect 23635 1455 23645 1475
rect 23605 1445 23645 1455
rect 23935 1475 23975 1485
rect 23935 1455 23945 1475
rect 23965 1455 23975 1475
rect 23935 1445 23975 1455
rect 24045 1475 24085 1485
rect 24045 1455 24055 1475
rect 24075 1455 24085 1475
rect 24045 1445 24085 1455
rect 24330 1475 24370 1485
rect 24330 1455 24340 1475
rect 24360 1455 24370 1475
rect 24330 1445 24370 1455
rect 24460 1475 24500 1485
rect 24460 1455 24470 1475
rect 24490 1455 24500 1475
rect 24460 1445 24500 1455
rect 24585 1475 24625 1485
rect 24585 1455 24595 1475
rect 24615 1455 24625 1475
rect 24585 1445 24625 1455
rect 24695 1475 24735 1485
rect 24695 1455 24705 1475
rect 24725 1455 24735 1475
rect 24695 1445 24735 1455
rect 24970 1475 25010 1485
rect 24970 1455 24980 1475
rect 25000 1455 25010 1475
rect 24970 1445 25010 1455
rect 25110 1475 25150 1485
rect 25110 1455 25120 1475
rect 25140 1455 25150 1475
rect 25110 1445 25150 1455
rect 25235 1475 25275 1485
rect 25235 1455 25245 1475
rect 25265 1455 25275 1475
rect 25235 1445 25275 1455
rect 25345 1475 25385 1485
rect 25345 1455 25355 1475
rect 25375 1455 25385 1475
rect 25345 1445 25385 1455
rect 25620 1475 25660 1485
rect 25620 1455 25630 1475
rect 25650 1455 25660 1475
rect 25620 1445 25660 1455
rect 25760 1475 25800 1485
rect 25760 1455 25770 1475
rect 25790 1455 25800 1475
rect 25760 1445 25800 1455
rect 25885 1475 25925 1485
rect 25885 1455 25895 1475
rect 25915 1455 25925 1475
rect 25885 1445 25925 1455
rect 25995 1475 26035 1485
rect 25995 1455 26005 1475
rect 26025 1455 26035 1475
rect 25995 1445 26035 1455
rect 26270 1475 26310 1485
rect 26270 1455 26280 1475
rect 26300 1455 26310 1475
rect 26270 1445 26310 1455
<< viali >>
rect 21340 1845 21360 1865
rect 21550 1845 21570 1865
rect 21885 1845 21905 1865
rect 22170 1845 22190 1865
rect 22545 1845 22565 1865
rect 22760 1845 22780 1865
rect 22980 1845 23000 1865
rect 23105 1845 23125 1865
rect 23215 1845 23235 1865
rect 23450 1845 23470 1865
rect 23670 1845 23690 1865
rect 23980 1845 24000 1865
rect 24150 1845 24170 1865
rect 24330 1845 24350 1865
rect 24630 1845 24650 1865
rect 24800 1845 24820 1865
rect 24980 1845 25000 1865
rect 25280 1845 25300 1865
rect 25450 1845 25470 1865
rect 25630 1845 25650 1865
rect 25930 1845 25950 1865
rect 26100 1845 26120 1865
rect 26280 1845 26300 1865
rect 21500 1790 21520 1810
rect 21595 1790 21615 1810
rect 21655 1780 21675 1800
rect 22060 1790 22080 1810
rect 22125 1790 22145 1810
rect 22710 1790 22730 1810
rect 22820 1790 22840 1810
rect 23385 1795 23405 1815
rect 23590 1795 23610 1815
rect 24565 1790 24585 1810
rect 24855 1790 24875 1810
rect 25215 1790 25235 1810
rect 25505 1790 25525 1810
rect 25865 1790 25885 1810
rect 26155 1790 26175 1810
rect 21130 1645 21150 1665
rect 22375 1730 22395 1750
rect 21985 1630 22005 1650
rect 22245 1630 22265 1650
rect 23125 1635 23145 1655
rect 21160 1510 21180 1530
rect 21655 1520 21675 1540
rect 21720 1515 21740 1535
rect 22190 1515 22210 1535
rect 22990 1515 23010 1535
rect 24292 1510 24312 1530
rect 26382 1644 26399 1661
rect 21260 1455 21280 1475
rect 21370 1455 21390 1475
rect 21605 1455 21625 1475
rect 21775 1455 21795 1475
rect 21885 1455 21905 1475
rect 22105 1455 22125 1475
rect 22340 1455 22360 1475
rect 22465 1455 22485 1475
rect 22575 1455 22595 1475
rect 22810 1455 22830 1475
rect 23040 1455 23060 1475
rect 23215 1455 23235 1475
rect 23340 1455 23360 1475
rect 23450 1455 23470 1475
rect 23615 1455 23635 1475
rect 23945 1455 23965 1475
rect 24055 1455 24075 1475
rect 24340 1455 24360 1475
rect 24470 1455 24490 1475
rect 24595 1455 24615 1475
rect 24705 1455 24725 1475
rect 24980 1455 25000 1475
rect 25120 1455 25140 1475
rect 25245 1455 25265 1475
rect 25355 1455 25375 1475
rect 25630 1455 25650 1475
rect 25770 1455 25790 1475
rect 25895 1455 25915 1475
rect 26005 1455 26025 1475
rect 26280 1455 26300 1475
<< metal1 >>
rect 21330 1870 21370 1875
rect 21330 1840 21335 1870
rect 21365 1840 21370 1870
rect 21330 1835 21370 1840
rect 21540 1870 21580 1875
rect 21540 1840 21545 1870
rect 21575 1840 21580 1870
rect 21540 1835 21580 1840
rect 21875 1870 21915 1875
rect 21875 1840 21880 1870
rect 21910 1840 21915 1870
rect 21875 1835 21915 1840
rect 22160 1870 22200 1875
rect 22160 1840 22165 1870
rect 22195 1840 22200 1870
rect 22160 1835 22200 1840
rect 22535 1870 22575 1875
rect 22535 1840 22540 1870
rect 22570 1840 22575 1870
rect 22535 1835 22575 1840
rect 22750 1870 22790 1875
rect 22750 1840 22755 1870
rect 22785 1840 22790 1870
rect 22750 1835 22790 1840
rect 22970 1870 23010 1875
rect 22970 1840 22975 1870
rect 23005 1840 23010 1870
rect 22970 1835 23010 1840
rect 23095 1870 23135 1875
rect 23095 1840 23100 1870
rect 23130 1840 23135 1870
rect 23095 1835 23135 1840
rect 23205 1870 23245 1875
rect 23205 1840 23210 1870
rect 23240 1840 23245 1870
rect 23205 1835 23245 1840
rect 23440 1870 23480 1875
rect 23440 1840 23445 1870
rect 23475 1840 23480 1870
rect 23440 1835 23480 1840
rect 23660 1870 23700 1875
rect 23660 1840 23665 1870
rect 23695 1840 23700 1870
rect 23660 1835 23700 1840
rect 23970 1870 24010 1875
rect 23970 1840 23975 1870
rect 24005 1840 24010 1870
rect 23970 1835 24010 1840
rect 24140 1870 24180 1875
rect 24140 1840 24145 1870
rect 24175 1840 24180 1870
rect 24140 1835 24180 1840
rect 24320 1870 24360 1875
rect 24320 1840 24325 1870
rect 24355 1840 24360 1870
rect 24320 1835 24360 1840
rect 24620 1870 24660 1875
rect 24620 1840 24625 1870
rect 24655 1840 24660 1870
rect 24620 1835 24660 1840
rect 24790 1870 24830 1875
rect 24790 1840 24795 1870
rect 24825 1840 24830 1870
rect 24790 1835 24830 1840
rect 24970 1870 25010 1875
rect 24970 1840 24975 1870
rect 25005 1840 25010 1870
rect 24970 1835 25010 1840
rect 25270 1870 25310 1875
rect 25270 1840 25275 1870
rect 25305 1840 25310 1870
rect 25270 1835 25310 1840
rect 25440 1870 25480 1875
rect 25440 1840 25445 1870
rect 25475 1840 25480 1870
rect 25440 1835 25480 1840
rect 25620 1870 25660 1875
rect 25620 1840 25625 1870
rect 25655 1840 25660 1870
rect 25620 1835 25660 1840
rect 25920 1870 25960 1875
rect 25920 1840 25925 1870
rect 25955 1840 25960 1870
rect 25920 1835 25960 1840
rect 26090 1870 26130 1875
rect 26090 1840 26095 1870
rect 26125 1840 26130 1870
rect 26090 1835 26130 1840
rect 26270 1870 26310 1875
rect 26270 1840 26275 1870
rect 26305 1840 26310 1870
rect 26270 1835 26310 1840
rect 21490 1810 21530 1820
rect 21490 1790 21500 1810
rect 21520 1800 21530 1810
rect 21590 1810 21625 1820
rect 22050 1810 22090 1820
rect 21590 1800 21595 1810
rect 21520 1790 21595 1800
rect 21615 1790 21625 1810
rect 21490 1780 21625 1790
rect 21645 1800 21685 1810
rect 22050 1800 22060 1810
rect 21645 1780 21655 1800
rect 21675 1790 22060 1800
rect 22080 1790 22090 1810
rect 21675 1780 22090 1790
rect 22120 1810 22150 1820
rect 22120 1790 22125 1810
rect 22145 1800 22150 1810
rect 22700 1810 22740 1820
rect 22145 1790 22385 1800
rect 22120 1780 22385 1790
rect 22700 1790 22710 1810
rect 22730 1800 22740 1810
rect 22810 1810 22850 1820
rect 22810 1800 22820 1810
rect 22730 1790 22820 1800
rect 22840 1790 22850 1810
rect 22700 1780 22850 1790
rect 23375 1815 23415 1820
rect 23375 1795 23385 1815
rect 23405 1805 23415 1815
rect 23580 1815 23620 1820
rect 23580 1805 23590 1815
rect 23405 1795 23590 1805
rect 23610 1795 23620 1815
rect 23375 1785 23620 1795
rect 24555 1810 24595 1820
rect 24555 1790 24565 1810
rect 24585 1800 24595 1810
rect 24845 1810 24885 1820
rect 24845 1800 24855 1810
rect 24585 1790 24855 1800
rect 24875 1790 24885 1810
rect 24555 1780 24885 1790
rect 25205 1810 25245 1820
rect 25205 1790 25215 1810
rect 25235 1800 25245 1810
rect 25495 1810 25535 1820
rect 25495 1800 25505 1810
rect 25235 1790 25505 1800
rect 25525 1790 25535 1810
rect 25205 1780 25535 1790
rect 25855 1810 25895 1820
rect 25855 1790 25865 1810
rect 25885 1800 25895 1810
rect 26145 1810 26185 1820
rect 26145 1800 26155 1810
rect 25885 1790 26155 1800
rect 26175 1790 26185 1810
rect 25855 1780 26185 1790
rect 21645 1770 21685 1780
rect 22365 1760 22385 1780
rect 24575 1760 24595 1780
rect 25225 1760 25245 1780
rect 25875 1760 25895 1780
rect 22365 1750 22405 1760
rect 22365 1730 22375 1750
rect 22395 1730 22405 1750
rect 22365 1720 22405 1730
rect 21120 1670 21160 1675
rect 21120 1640 21125 1670
rect 21155 1640 21160 1670
rect 26376 1665 26405 1670
rect 23115 1655 23155 1665
rect 21120 1635 21160 1640
rect 21975 1650 22275 1655
rect 21975 1630 21985 1650
rect 22005 1635 22245 1650
rect 22005 1630 22015 1635
rect 21975 1620 22015 1630
rect 22235 1630 22245 1635
rect 22265 1630 22275 1650
rect 22235 1620 22275 1630
rect 23115 1635 23125 1655
rect 23145 1635 23155 1655
rect 23115 1625 23155 1635
rect 26376 1639 26378 1665
rect 26404 1639 26405 1665
rect 26376 1630 26405 1639
rect 21645 1540 21685 1550
rect 23115 1540 23135 1625
rect 21150 1530 21190 1540
rect 21645 1530 21655 1540
rect 21150 1510 21160 1530
rect 21180 1520 21655 1530
rect 21675 1520 21685 1540
rect 21180 1510 21685 1520
rect 21710 1535 21750 1540
rect 21710 1515 21720 1535
rect 21740 1525 21750 1535
rect 22180 1535 22220 1540
rect 22180 1525 22190 1535
rect 21740 1515 22190 1525
rect 22210 1525 22220 1535
rect 22980 1535 23020 1540
rect 22980 1525 22990 1535
rect 22210 1515 22990 1525
rect 23010 1515 23020 1535
rect 23115 1530 24320 1540
rect 23115 1520 24292 1530
rect 21150 1500 21190 1510
rect 21710 1505 23020 1515
rect 24287 1510 24292 1520
rect 24312 1510 24320 1530
rect 24287 1500 24320 1510
rect 21250 1480 21290 1485
rect 21250 1450 21255 1480
rect 21285 1450 21290 1480
rect 21250 1445 21290 1450
rect 21360 1480 21400 1485
rect 21360 1450 21365 1480
rect 21395 1450 21400 1480
rect 21360 1445 21400 1450
rect 21595 1480 21635 1485
rect 21595 1450 21600 1480
rect 21630 1450 21635 1480
rect 21595 1445 21635 1450
rect 21765 1480 21805 1485
rect 21765 1450 21770 1480
rect 21800 1450 21805 1480
rect 21765 1445 21805 1450
rect 21875 1480 21915 1485
rect 21875 1450 21880 1480
rect 21910 1450 21915 1480
rect 21875 1445 21915 1450
rect 22095 1480 22135 1485
rect 22095 1450 22100 1480
rect 22130 1450 22135 1480
rect 22095 1445 22135 1450
rect 22330 1480 22370 1485
rect 22330 1450 22335 1480
rect 22365 1450 22370 1480
rect 22330 1445 22370 1450
rect 22455 1480 22495 1485
rect 22455 1450 22460 1480
rect 22490 1450 22495 1480
rect 22455 1445 22495 1450
rect 22565 1480 22605 1485
rect 22565 1450 22570 1480
rect 22600 1450 22605 1480
rect 22565 1445 22605 1450
rect 22800 1480 22840 1485
rect 22800 1450 22805 1480
rect 22835 1450 22840 1480
rect 22800 1445 22840 1450
rect 23030 1480 23070 1485
rect 23030 1450 23035 1480
rect 23065 1450 23070 1480
rect 23030 1445 23070 1450
rect 23205 1480 23245 1485
rect 23205 1450 23210 1480
rect 23240 1450 23245 1480
rect 23205 1445 23245 1450
rect 23330 1480 23370 1485
rect 23330 1450 23335 1480
rect 23365 1450 23370 1480
rect 23330 1445 23370 1450
rect 23440 1480 23480 1485
rect 23440 1450 23445 1480
rect 23475 1450 23480 1480
rect 23440 1445 23480 1450
rect 23605 1480 23645 1485
rect 23605 1450 23610 1480
rect 23640 1450 23645 1480
rect 23605 1445 23645 1450
rect 23935 1480 23975 1485
rect 23935 1450 23940 1480
rect 23970 1450 23975 1480
rect 23935 1445 23975 1450
rect 24045 1480 24085 1485
rect 24045 1450 24050 1480
rect 24080 1450 24085 1480
rect 24045 1445 24085 1450
rect 24330 1480 24370 1485
rect 24330 1450 24335 1480
rect 24365 1450 24370 1480
rect 24330 1445 24370 1450
rect 24460 1480 24500 1485
rect 24460 1450 24465 1480
rect 24495 1450 24500 1480
rect 24460 1445 24500 1450
rect 24585 1480 24625 1485
rect 24585 1450 24590 1480
rect 24620 1450 24625 1480
rect 24585 1445 24625 1450
rect 24695 1480 24735 1485
rect 24695 1450 24700 1480
rect 24730 1450 24735 1480
rect 24695 1445 24735 1450
rect 24970 1480 25010 1485
rect 24970 1450 24975 1480
rect 25005 1450 25010 1480
rect 24970 1445 25010 1450
rect 25110 1480 25150 1485
rect 25110 1450 25115 1480
rect 25145 1450 25150 1480
rect 25110 1445 25150 1450
rect 25235 1480 25275 1485
rect 25235 1450 25240 1480
rect 25270 1450 25275 1480
rect 25235 1445 25275 1450
rect 25345 1480 25385 1485
rect 25345 1450 25350 1480
rect 25380 1450 25385 1480
rect 25345 1445 25385 1450
rect 25620 1480 25660 1485
rect 25620 1450 25625 1480
rect 25655 1450 25660 1480
rect 25620 1445 25660 1450
rect 25760 1480 25800 1485
rect 25760 1450 25765 1480
rect 25795 1450 25800 1480
rect 25760 1445 25800 1450
rect 25885 1480 25925 1485
rect 25885 1450 25890 1480
rect 25920 1450 25925 1480
rect 25885 1445 25925 1450
rect 25995 1480 26035 1485
rect 25995 1450 26000 1480
rect 26030 1450 26035 1480
rect 25995 1445 26035 1450
rect 26270 1480 26310 1485
rect 26270 1450 26275 1480
rect 26305 1450 26310 1480
rect 26270 1445 26310 1450
<< via1 >>
rect 21335 1865 21365 1870
rect 21335 1845 21340 1865
rect 21340 1845 21360 1865
rect 21360 1845 21365 1865
rect 21335 1840 21365 1845
rect 21545 1865 21575 1870
rect 21545 1845 21550 1865
rect 21550 1845 21570 1865
rect 21570 1845 21575 1865
rect 21545 1840 21575 1845
rect 21880 1865 21910 1870
rect 21880 1845 21885 1865
rect 21885 1845 21905 1865
rect 21905 1845 21910 1865
rect 21880 1840 21910 1845
rect 22165 1865 22195 1870
rect 22165 1845 22170 1865
rect 22170 1845 22190 1865
rect 22190 1845 22195 1865
rect 22165 1840 22195 1845
rect 22540 1865 22570 1870
rect 22540 1845 22545 1865
rect 22545 1845 22565 1865
rect 22565 1845 22570 1865
rect 22540 1840 22570 1845
rect 22755 1865 22785 1870
rect 22755 1845 22760 1865
rect 22760 1845 22780 1865
rect 22780 1845 22785 1865
rect 22755 1840 22785 1845
rect 22975 1865 23005 1870
rect 22975 1845 22980 1865
rect 22980 1845 23000 1865
rect 23000 1845 23005 1865
rect 22975 1840 23005 1845
rect 23100 1865 23130 1870
rect 23100 1845 23105 1865
rect 23105 1845 23125 1865
rect 23125 1845 23130 1865
rect 23100 1840 23130 1845
rect 23210 1865 23240 1870
rect 23210 1845 23215 1865
rect 23215 1845 23235 1865
rect 23235 1845 23240 1865
rect 23210 1840 23240 1845
rect 23445 1865 23475 1870
rect 23445 1845 23450 1865
rect 23450 1845 23470 1865
rect 23470 1845 23475 1865
rect 23445 1840 23475 1845
rect 23665 1865 23695 1870
rect 23665 1845 23670 1865
rect 23670 1845 23690 1865
rect 23690 1845 23695 1865
rect 23665 1840 23695 1845
rect 23975 1865 24005 1870
rect 23975 1845 23980 1865
rect 23980 1845 24000 1865
rect 24000 1845 24005 1865
rect 23975 1840 24005 1845
rect 24145 1865 24175 1870
rect 24145 1845 24150 1865
rect 24150 1845 24170 1865
rect 24170 1845 24175 1865
rect 24145 1840 24175 1845
rect 24325 1865 24355 1870
rect 24325 1845 24330 1865
rect 24330 1845 24350 1865
rect 24350 1845 24355 1865
rect 24325 1840 24355 1845
rect 24625 1865 24655 1870
rect 24625 1845 24630 1865
rect 24630 1845 24650 1865
rect 24650 1845 24655 1865
rect 24625 1840 24655 1845
rect 24795 1865 24825 1870
rect 24795 1845 24800 1865
rect 24800 1845 24820 1865
rect 24820 1845 24825 1865
rect 24795 1840 24825 1845
rect 24975 1865 25005 1870
rect 24975 1845 24980 1865
rect 24980 1845 25000 1865
rect 25000 1845 25005 1865
rect 24975 1840 25005 1845
rect 25275 1865 25305 1870
rect 25275 1845 25280 1865
rect 25280 1845 25300 1865
rect 25300 1845 25305 1865
rect 25275 1840 25305 1845
rect 25445 1865 25475 1870
rect 25445 1845 25450 1865
rect 25450 1845 25470 1865
rect 25470 1845 25475 1865
rect 25445 1840 25475 1845
rect 25625 1865 25655 1870
rect 25625 1845 25630 1865
rect 25630 1845 25650 1865
rect 25650 1845 25655 1865
rect 25625 1840 25655 1845
rect 25925 1865 25955 1870
rect 25925 1845 25930 1865
rect 25930 1845 25950 1865
rect 25950 1845 25955 1865
rect 25925 1840 25955 1845
rect 26095 1865 26125 1870
rect 26095 1845 26100 1865
rect 26100 1845 26120 1865
rect 26120 1845 26125 1865
rect 26095 1840 26125 1845
rect 26275 1865 26305 1870
rect 26275 1845 26280 1865
rect 26280 1845 26300 1865
rect 26300 1845 26305 1865
rect 26275 1840 26305 1845
rect 21125 1665 21155 1670
rect 21125 1645 21130 1665
rect 21130 1645 21150 1665
rect 21150 1645 21155 1665
rect 21125 1640 21155 1645
rect 26378 1661 26404 1665
rect 26378 1644 26382 1661
rect 26382 1644 26399 1661
rect 26399 1644 26404 1661
rect 26378 1639 26404 1644
rect 21255 1475 21285 1480
rect 21255 1455 21260 1475
rect 21260 1455 21280 1475
rect 21280 1455 21285 1475
rect 21255 1450 21285 1455
rect 21365 1475 21395 1480
rect 21365 1455 21370 1475
rect 21370 1455 21390 1475
rect 21390 1455 21395 1475
rect 21365 1450 21395 1455
rect 21600 1475 21630 1480
rect 21600 1455 21605 1475
rect 21605 1455 21625 1475
rect 21625 1455 21630 1475
rect 21600 1450 21630 1455
rect 21770 1475 21800 1480
rect 21770 1455 21775 1475
rect 21775 1455 21795 1475
rect 21795 1455 21800 1475
rect 21770 1450 21800 1455
rect 21880 1475 21910 1480
rect 21880 1455 21885 1475
rect 21885 1455 21905 1475
rect 21905 1455 21910 1475
rect 21880 1450 21910 1455
rect 22100 1475 22130 1480
rect 22100 1455 22105 1475
rect 22105 1455 22125 1475
rect 22125 1455 22130 1475
rect 22100 1450 22130 1455
rect 22335 1475 22365 1480
rect 22335 1455 22340 1475
rect 22340 1455 22360 1475
rect 22360 1455 22365 1475
rect 22335 1450 22365 1455
rect 22460 1475 22490 1480
rect 22460 1455 22465 1475
rect 22465 1455 22485 1475
rect 22485 1455 22490 1475
rect 22460 1450 22490 1455
rect 22570 1475 22600 1480
rect 22570 1455 22575 1475
rect 22575 1455 22595 1475
rect 22595 1455 22600 1475
rect 22570 1450 22600 1455
rect 22805 1475 22835 1480
rect 22805 1455 22810 1475
rect 22810 1455 22830 1475
rect 22830 1455 22835 1475
rect 22805 1450 22835 1455
rect 23035 1475 23065 1480
rect 23035 1455 23040 1475
rect 23040 1455 23060 1475
rect 23060 1455 23065 1475
rect 23035 1450 23065 1455
rect 23210 1475 23240 1480
rect 23210 1455 23215 1475
rect 23215 1455 23235 1475
rect 23235 1455 23240 1475
rect 23210 1450 23240 1455
rect 23335 1475 23365 1480
rect 23335 1455 23340 1475
rect 23340 1455 23360 1475
rect 23360 1455 23365 1475
rect 23335 1450 23365 1455
rect 23445 1475 23475 1480
rect 23445 1455 23450 1475
rect 23450 1455 23470 1475
rect 23470 1455 23475 1475
rect 23445 1450 23475 1455
rect 23610 1475 23640 1480
rect 23610 1455 23615 1475
rect 23615 1455 23635 1475
rect 23635 1455 23640 1475
rect 23610 1450 23640 1455
rect 23940 1475 23970 1480
rect 23940 1455 23945 1475
rect 23945 1455 23965 1475
rect 23965 1455 23970 1475
rect 23940 1450 23970 1455
rect 24050 1475 24080 1480
rect 24050 1455 24055 1475
rect 24055 1455 24075 1475
rect 24075 1455 24080 1475
rect 24050 1450 24080 1455
rect 24335 1475 24365 1480
rect 24335 1455 24340 1475
rect 24340 1455 24360 1475
rect 24360 1455 24365 1475
rect 24335 1450 24365 1455
rect 24465 1475 24495 1480
rect 24465 1455 24470 1475
rect 24470 1455 24490 1475
rect 24490 1455 24495 1475
rect 24465 1450 24495 1455
rect 24590 1475 24620 1480
rect 24590 1455 24595 1475
rect 24595 1455 24615 1475
rect 24615 1455 24620 1475
rect 24590 1450 24620 1455
rect 24700 1475 24730 1480
rect 24700 1455 24705 1475
rect 24705 1455 24725 1475
rect 24725 1455 24730 1475
rect 24700 1450 24730 1455
rect 24975 1475 25005 1480
rect 24975 1455 24980 1475
rect 24980 1455 25000 1475
rect 25000 1455 25005 1475
rect 24975 1450 25005 1455
rect 25115 1475 25145 1480
rect 25115 1455 25120 1475
rect 25120 1455 25140 1475
rect 25140 1455 25145 1475
rect 25115 1450 25145 1455
rect 25240 1475 25270 1480
rect 25240 1455 25245 1475
rect 25245 1455 25265 1475
rect 25265 1455 25270 1475
rect 25240 1450 25270 1455
rect 25350 1475 25380 1480
rect 25350 1455 25355 1475
rect 25355 1455 25375 1475
rect 25375 1455 25380 1475
rect 25350 1450 25380 1455
rect 25625 1475 25655 1480
rect 25625 1455 25630 1475
rect 25630 1455 25650 1475
rect 25650 1455 25655 1475
rect 25625 1450 25655 1455
rect 25765 1475 25795 1480
rect 25765 1455 25770 1475
rect 25770 1455 25790 1475
rect 25790 1455 25795 1475
rect 25765 1450 25795 1455
rect 25890 1475 25920 1480
rect 25890 1455 25895 1475
rect 25895 1455 25915 1475
rect 25915 1455 25920 1475
rect 25890 1450 25920 1455
rect 26000 1475 26030 1480
rect 26000 1455 26005 1475
rect 26005 1455 26025 1475
rect 26025 1455 26030 1475
rect 26000 1450 26030 1455
rect 26275 1475 26305 1480
rect 26275 1455 26280 1475
rect 26280 1455 26300 1475
rect 26300 1455 26305 1475
rect 26275 1450 26305 1455
<< metal2 >>
rect 21130 1870 26310 1875
rect 21130 1840 21335 1870
rect 21365 1840 21545 1870
rect 21575 1840 21880 1870
rect 21910 1840 22165 1870
rect 22195 1840 22540 1870
rect 22570 1840 22755 1870
rect 22785 1840 22975 1870
rect 23005 1840 23100 1870
rect 23130 1840 23210 1870
rect 23240 1840 23445 1870
rect 23475 1840 23665 1870
rect 23695 1840 23975 1870
rect 24005 1840 24145 1870
rect 24175 1840 24325 1870
rect 24355 1840 24625 1870
rect 24655 1840 24795 1870
rect 24825 1840 24975 1870
rect 25005 1840 25275 1870
rect 25305 1840 25445 1870
rect 25475 1840 25625 1870
rect 25655 1840 25925 1870
rect 25955 1840 26095 1870
rect 26125 1840 26275 1870
rect 26305 1840 26310 1870
rect 21130 1835 26310 1840
rect 21065 1670 21160 1675
rect 21065 1640 21125 1670
rect 21155 1640 21160 1670
rect 21065 1635 21160 1640
rect 26376 1665 26405 1670
rect 26376 1639 26378 1665
rect 26404 1639 26405 1665
rect 26376 1630 26405 1639
rect 21130 1480 26310 1485
rect 21130 1450 21255 1480
rect 21285 1450 21365 1480
rect 21395 1450 21600 1480
rect 21630 1450 21770 1480
rect 21800 1450 21880 1480
rect 21910 1450 22100 1480
rect 22130 1450 22335 1480
rect 22365 1450 22460 1480
rect 22490 1450 22570 1480
rect 22600 1450 22805 1480
rect 22835 1450 23035 1480
rect 23065 1450 23210 1480
rect 23240 1450 23335 1480
rect 23365 1450 23445 1480
rect 23475 1450 23610 1480
rect 23640 1450 23940 1480
rect 23970 1450 24050 1480
rect 24080 1450 24335 1480
rect 24365 1450 24465 1480
rect 24495 1450 24590 1480
rect 24620 1450 24700 1480
rect 24730 1450 24975 1480
rect 25005 1450 25115 1480
rect 25145 1450 25240 1480
rect 25270 1450 25350 1480
rect 25380 1450 25625 1480
rect 25655 1450 25765 1480
rect 25795 1450 25890 1480
rect 25920 1450 26000 1480
rect 26030 1450 26275 1480
rect 26305 1450 26310 1480
rect 21130 1445 26310 1450
<< end >>
