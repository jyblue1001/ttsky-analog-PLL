magic
tech sky130A
timestamp 1757089157
<< nwell >>
rect 6130 1695 11385 1800
<< nmos >>
rect 6235 1555 6250 1605
rect 6290 1555 6305 1605
rect 6345 1555 6360 1605
rect 6400 1555 6415 1605
rect 6525 1555 6540 1605
rect 6580 1555 6595 1605
rect 6750 1555 6765 1605
rect 6805 1555 6820 1605
rect 6860 1555 6875 1605
rect 6915 1555 6930 1605
rect 7080 1555 7095 1605
rect 7135 1555 7150 1605
rect 7190 1555 7205 1605
rect 7245 1555 7260 1605
rect 7440 1555 7455 1605
rect 7495 1555 7510 1605
rect 7550 1555 7565 1605
rect 7605 1555 7620 1605
rect 7730 1555 7745 1605
rect 7785 1555 7800 1605
rect 8010 1555 8025 1605
rect 8190 1555 8205 1605
rect 8315 1555 8330 1605
rect 8370 1555 8385 1605
rect 8425 1555 8440 1605
rect 8480 1555 8495 1605
rect 8645 1555 8660 1605
rect 8700 1555 8715 1605
rect 8755 1555 8770 1605
rect 8920 1555 8935 1605
rect 8975 1555 8990 1605
rect 9030 1555 9045 1605
rect 9085 1555 9100 1605
rect 9250 1555 9265 1605
rect 9305 1555 9320 1605
rect 9360 1555 9375 1605
rect 9570 1510 9585 1560
rect 9625 1510 9640 1560
rect 9680 1510 9695 1560
rect 9735 1510 9750 1560
rect 9900 1510 9915 1560
rect 9955 1510 9970 1560
rect 10010 1510 10025 1560
rect 10220 1510 10235 1560
rect 10275 1510 10290 1560
rect 10330 1510 10345 1560
rect 10385 1510 10400 1560
rect 10550 1510 10565 1560
rect 10605 1510 10620 1560
rect 10660 1510 10675 1560
rect 10870 1510 10885 1560
rect 10925 1510 10940 1560
rect 10980 1510 10995 1560
rect 11035 1510 11050 1560
rect 11200 1510 11215 1560
rect 11255 1510 11270 1560
rect 11310 1510 11325 1560
<< pmos >>
rect 6315 1715 6330 1765
rect 6525 1715 6540 1765
rect 6580 1715 6595 1765
rect 6860 1715 6875 1765
rect 6915 1715 6930 1765
rect 7080 1715 7095 1765
rect 7135 1715 7150 1765
rect 7190 1715 7205 1765
rect 7520 1715 7535 1765
rect 7730 1715 7745 1765
rect 7785 1715 7800 1765
rect 7955 1715 7970 1765
rect 8010 1715 8025 1765
rect 8135 1715 8150 1765
rect 8190 1715 8205 1765
rect 8425 1715 8440 1765
rect 8480 1715 8495 1765
rect 8645 1715 8660 1765
rect 8700 1715 8715 1765
rect 8955 1715 8970 1765
rect 9125 1715 9140 1765
rect 9180 1715 9195 1765
rect 9305 1715 9320 1765
rect 9360 1715 9375 1765
rect 9605 1715 9620 1765
rect 9775 1715 9790 1765
rect 9830 1715 9845 1765
rect 9955 1715 9970 1765
rect 10010 1715 10025 1765
rect 10255 1715 10270 1765
rect 10425 1715 10440 1765
rect 10480 1715 10495 1765
rect 10605 1715 10620 1765
rect 10660 1715 10675 1765
rect 10905 1715 10920 1765
rect 11075 1715 11090 1765
rect 11130 1715 11145 1765
rect 11255 1715 11270 1765
rect 11310 1715 11325 1765
<< ndiff >>
rect 6195 1590 6235 1605
rect 6195 1570 6205 1590
rect 6225 1570 6235 1590
rect 6195 1555 6235 1570
rect 6250 1590 6290 1605
rect 6250 1570 6260 1590
rect 6280 1570 6290 1590
rect 6250 1555 6290 1570
rect 6305 1590 6345 1605
rect 6305 1570 6315 1590
rect 6335 1570 6345 1590
rect 6305 1555 6345 1570
rect 6360 1590 6400 1605
rect 6360 1570 6370 1590
rect 6390 1570 6400 1590
rect 6360 1555 6400 1570
rect 6415 1590 6455 1605
rect 6415 1570 6425 1590
rect 6445 1570 6455 1590
rect 6415 1555 6455 1570
rect 6485 1590 6525 1605
rect 6485 1570 6495 1590
rect 6515 1570 6525 1590
rect 6485 1555 6525 1570
rect 6540 1590 6580 1605
rect 6540 1570 6550 1590
rect 6570 1570 6580 1590
rect 6540 1555 6580 1570
rect 6595 1590 6635 1605
rect 6595 1570 6605 1590
rect 6625 1570 6635 1590
rect 6595 1555 6635 1570
rect 6710 1590 6750 1605
rect 6710 1570 6720 1590
rect 6740 1570 6750 1590
rect 6710 1555 6750 1570
rect 6765 1590 6805 1605
rect 6765 1570 6775 1590
rect 6795 1570 6805 1590
rect 6765 1555 6805 1570
rect 6820 1590 6860 1605
rect 6820 1570 6830 1590
rect 6850 1570 6860 1590
rect 6820 1555 6860 1570
rect 6875 1590 6915 1605
rect 6875 1570 6885 1590
rect 6905 1570 6915 1590
rect 6875 1555 6915 1570
rect 6930 1590 6970 1605
rect 6930 1570 6940 1590
rect 6960 1570 6970 1590
rect 6930 1555 6970 1570
rect 7040 1590 7080 1605
rect 7040 1570 7050 1590
rect 7070 1570 7080 1590
rect 7040 1555 7080 1570
rect 7095 1590 7135 1605
rect 7095 1570 7105 1590
rect 7125 1570 7135 1590
rect 7095 1555 7135 1570
rect 7150 1590 7190 1605
rect 7150 1570 7160 1590
rect 7180 1570 7190 1590
rect 7150 1555 7190 1570
rect 7205 1590 7245 1605
rect 7205 1570 7215 1590
rect 7235 1570 7245 1590
rect 7205 1555 7245 1570
rect 7260 1590 7300 1605
rect 7260 1570 7270 1590
rect 7290 1570 7300 1590
rect 7260 1555 7300 1570
rect 7400 1590 7440 1605
rect 7400 1570 7410 1590
rect 7430 1570 7440 1590
rect 7400 1555 7440 1570
rect 7455 1590 7495 1605
rect 7455 1570 7465 1590
rect 7485 1570 7495 1590
rect 7455 1555 7495 1570
rect 7510 1590 7550 1605
rect 7510 1570 7520 1590
rect 7540 1570 7550 1590
rect 7510 1555 7550 1570
rect 7565 1590 7605 1605
rect 7565 1570 7575 1590
rect 7595 1570 7605 1590
rect 7565 1555 7605 1570
rect 7620 1590 7660 1605
rect 7620 1570 7630 1590
rect 7650 1570 7660 1590
rect 7620 1555 7660 1570
rect 7690 1590 7730 1605
rect 7690 1570 7700 1590
rect 7720 1570 7730 1590
rect 7690 1555 7730 1570
rect 7745 1590 7785 1605
rect 7745 1570 7755 1590
rect 7775 1570 7785 1590
rect 7745 1555 7785 1570
rect 7800 1590 7840 1605
rect 7800 1570 7810 1590
rect 7830 1570 7840 1590
rect 7800 1555 7840 1570
rect 7970 1590 8010 1605
rect 7970 1570 7980 1590
rect 8000 1570 8010 1590
rect 7970 1555 8010 1570
rect 8025 1590 8065 1605
rect 8025 1570 8035 1590
rect 8055 1570 8065 1590
rect 8025 1555 8065 1570
rect 8150 1590 8190 1605
rect 8150 1570 8160 1590
rect 8180 1570 8190 1590
rect 8150 1555 8190 1570
rect 8205 1590 8245 1605
rect 8205 1570 8215 1590
rect 8235 1570 8245 1590
rect 8205 1555 8245 1570
rect 8275 1590 8315 1605
rect 8275 1570 8285 1590
rect 8305 1570 8315 1590
rect 8275 1555 8315 1570
rect 8330 1590 8370 1605
rect 8330 1570 8340 1590
rect 8360 1570 8370 1590
rect 8330 1555 8370 1570
rect 8385 1590 8425 1605
rect 8385 1570 8395 1590
rect 8415 1570 8425 1590
rect 8385 1555 8425 1570
rect 8440 1590 8480 1605
rect 8440 1570 8450 1590
rect 8470 1570 8480 1590
rect 8440 1555 8480 1570
rect 8495 1590 8535 1605
rect 8495 1570 8505 1590
rect 8525 1570 8535 1590
rect 8495 1555 8535 1570
rect 8605 1590 8645 1605
rect 8605 1570 8615 1590
rect 8635 1570 8645 1590
rect 8605 1555 8645 1570
rect 8660 1590 8700 1605
rect 8660 1570 8670 1590
rect 8690 1570 8700 1590
rect 8660 1555 8700 1570
rect 8715 1590 8755 1605
rect 8715 1570 8725 1590
rect 8745 1570 8755 1590
rect 8715 1555 8755 1570
rect 8770 1590 8810 1605
rect 8770 1570 8780 1590
rect 8800 1570 8810 1590
rect 8770 1555 8810 1570
rect 8880 1590 8920 1605
rect 8880 1570 8890 1590
rect 8910 1570 8920 1590
rect 8880 1555 8920 1570
rect 8935 1590 8975 1605
rect 8935 1570 8945 1590
rect 8965 1570 8975 1590
rect 8935 1555 8975 1570
rect 8990 1590 9030 1605
rect 8990 1570 9000 1590
rect 9020 1570 9030 1590
rect 8990 1555 9030 1570
rect 9045 1590 9085 1605
rect 9045 1570 9055 1590
rect 9075 1570 9085 1590
rect 9045 1555 9085 1570
rect 9100 1590 9140 1605
rect 9100 1570 9110 1590
rect 9130 1570 9140 1590
rect 9100 1555 9140 1570
rect 9210 1590 9250 1605
rect 9210 1570 9220 1590
rect 9240 1570 9250 1590
rect 9210 1555 9250 1570
rect 9265 1590 9305 1605
rect 9265 1570 9275 1590
rect 9295 1570 9305 1590
rect 9265 1555 9305 1570
rect 9320 1590 9360 1605
rect 9320 1570 9330 1590
rect 9350 1570 9360 1590
rect 9320 1555 9360 1570
rect 9375 1590 9415 1605
rect 9375 1570 9385 1590
rect 9405 1570 9415 1590
rect 9375 1555 9415 1570
rect 9530 1545 9570 1560
rect 9530 1525 9540 1545
rect 9560 1525 9570 1545
rect 9530 1510 9570 1525
rect 9585 1545 9625 1560
rect 9585 1525 9595 1545
rect 9615 1525 9625 1545
rect 9585 1510 9625 1525
rect 9640 1545 9680 1560
rect 9640 1525 9650 1545
rect 9670 1525 9680 1545
rect 9640 1510 9680 1525
rect 9695 1545 9735 1560
rect 9695 1525 9705 1545
rect 9725 1525 9735 1545
rect 9695 1510 9735 1525
rect 9750 1545 9790 1560
rect 9750 1525 9760 1545
rect 9780 1525 9790 1545
rect 9750 1510 9790 1525
rect 9860 1545 9900 1560
rect 9860 1525 9870 1545
rect 9890 1525 9900 1545
rect 9860 1510 9900 1525
rect 9915 1545 9955 1560
rect 9915 1525 9925 1545
rect 9945 1525 9955 1545
rect 9915 1510 9955 1525
rect 9970 1545 10010 1560
rect 9970 1525 9980 1545
rect 10000 1525 10010 1545
rect 9970 1510 10010 1525
rect 10025 1545 10065 1560
rect 10025 1525 10035 1545
rect 10055 1525 10065 1545
rect 10025 1510 10065 1525
rect 10180 1545 10220 1560
rect 10180 1525 10190 1545
rect 10210 1525 10220 1545
rect 10180 1510 10220 1525
rect 10235 1545 10275 1560
rect 10235 1525 10245 1545
rect 10265 1525 10275 1545
rect 10235 1510 10275 1525
rect 10290 1545 10330 1560
rect 10290 1525 10300 1545
rect 10320 1525 10330 1545
rect 10290 1510 10330 1525
rect 10345 1545 10385 1560
rect 10345 1525 10355 1545
rect 10375 1525 10385 1545
rect 10345 1510 10385 1525
rect 10400 1545 10440 1560
rect 10400 1525 10410 1545
rect 10430 1525 10440 1545
rect 10400 1510 10440 1525
rect 10510 1545 10550 1560
rect 10510 1525 10520 1545
rect 10540 1525 10550 1545
rect 10510 1510 10550 1525
rect 10565 1545 10605 1560
rect 10565 1525 10575 1545
rect 10595 1525 10605 1545
rect 10565 1510 10605 1525
rect 10620 1545 10660 1560
rect 10620 1525 10630 1545
rect 10650 1525 10660 1545
rect 10620 1510 10660 1525
rect 10675 1545 10715 1560
rect 10675 1525 10685 1545
rect 10705 1525 10715 1545
rect 10675 1510 10715 1525
rect 10830 1545 10870 1560
rect 10830 1525 10840 1545
rect 10860 1525 10870 1545
rect 10830 1510 10870 1525
rect 10885 1545 10925 1560
rect 10885 1525 10895 1545
rect 10915 1525 10925 1545
rect 10885 1510 10925 1525
rect 10940 1545 10980 1560
rect 10940 1525 10950 1545
rect 10970 1525 10980 1545
rect 10940 1510 10980 1525
rect 10995 1545 11035 1560
rect 10995 1525 11005 1545
rect 11025 1525 11035 1545
rect 10995 1510 11035 1525
rect 11050 1545 11090 1560
rect 11050 1525 11060 1545
rect 11080 1525 11090 1545
rect 11050 1510 11090 1525
rect 11160 1545 11200 1560
rect 11160 1525 11170 1545
rect 11190 1525 11200 1545
rect 11160 1510 11200 1525
rect 11215 1545 11255 1560
rect 11215 1525 11225 1545
rect 11245 1525 11255 1545
rect 11215 1510 11255 1525
rect 11270 1545 11310 1560
rect 11270 1525 11280 1545
rect 11300 1525 11310 1545
rect 11270 1510 11310 1525
rect 11325 1545 11365 1560
rect 11325 1525 11335 1545
rect 11355 1525 11365 1545
rect 11325 1510 11365 1525
<< pdiff >>
rect 6275 1750 6315 1765
rect 6275 1730 6285 1750
rect 6305 1730 6315 1750
rect 6275 1715 6315 1730
rect 6330 1750 6370 1765
rect 6330 1730 6340 1750
rect 6360 1730 6370 1750
rect 6330 1715 6370 1730
rect 6485 1750 6525 1765
rect 6485 1730 6495 1750
rect 6515 1730 6525 1750
rect 6485 1715 6525 1730
rect 6540 1750 6580 1765
rect 6540 1730 6550 1750
rect 6570 1730 6580 1750
rect 6540 1715 6580 1730
rect 6595 1750 6635 1765
rect 6595 1730 6605 1750
rect 6625 1730 6635 1750
rect 6595 1715 6635 1730
rect 6820 1750 6860 1765
rect 6820 1730 6830 1750
rect 6850 1730 6860 1750
rect 6820 1715 6860 1730
rect 6875 1750 6915 1765
rect 6875 1730 6885 1750
rect 6905 1730 6915 1750
rect 6875 1715 6915 1730
rect 6930 1750 6970 1765
rect 6930 1730 6940 1750
rect 6960 1730 6970 1750
rect 6930 1715 6970 1730
rect 7040 1750 7080 1765
rect 7040 1730 7050 1750
rect 7070 1730 7080 1750
rect 7040 1715 7080 1730
rect 7095 1750 7135 1765
rect 7095 1730 7105 1750
rect 7125 1730 7135 1750
rect 7095 1715 7135 1730
rect 7150 1750 7190 1765
rect 7150 1730 7160 1750
rect 7180 1730 7190 1750
rect 7150 1715 7190 1730
rect 7205 1750 7245 1765
rect 7205 1730 7215 1750
rect 7235 1730 7245 1750
rect 7205 1715 7245 1730
rect 7480 1750 7520 1765
rect 7480 1730 7490 1750
rect 7510 1730 7520 1750
rect 7480 1715 7520 1730
rect 7535 1750 7575 1765
rect 7535 1730 7545 1750
rect 7565 1730 7575 1750
rect 7535 1715 7575 1730
rect 7690 1750 7730 1765
rect 7690 1730 7700 1750
rect 7720 1730 7730 1750
rect 7690 1715 7730 1730
rect 7745 1750 7785 1765
rect 7745 1730 7755 1750
rect 7775 1730 7785 1750
rect 7745 1715 7785 1730
rect 7800 1750 7840 1765
rect 7800 1730 7810 1750
rect 7830 1730 7840 1750
rect 7800 1715 7840 1730
rect 7915 1750 7955 1765
rect 7915 1730 7925 1750
rect 7945 1730 7955 1750
rect 7915 1715 7955 1730
rect 7970 1750 8010 1765
rect 7970 1730 7980 1750
rect 8000 1730 8010 1750
rect 7970 1715 8010 1730
rect 8025 1750 8065 1765
rect 8025 1730 8035 1750
rect 8055 1730 8065 1750
rect 8025 1715 8065 1730
rect 8095 1750 8135 1765
rect 8095 1730 8105 1750
rect 8125 1730 8135 1750
rect 8095 1715 8135 1730
rect 8150 1750 8190 1765
rect 8150 1730 8160 1750
rect 8180 1730 8190 1750
rect 8150 1715 8190 1730
rect 8205 1750 8245 1765
rect 8205 1730 8215 1750
rect 8235 1730 8245 1750
rect 8205 1715 8245 1730
rect 8385 1750 8425 1765
rect 8385 1730 8395 1750
rect 8415 1730 8425 1750
rect 8385 1715 8425 1730
rect 8440 1750 8480 1765
rect 8440 1730 8450 1750
rect 8470 1730 8480 1750
rect 8440 1715 8480 1730
rect 8495 1750 8535 1765
rect 8495 1730 8505 1750
rect 8525 1730 8535 1750
rect 8495 1715 8535 1730
rect 8605 1750 8645 1765
rect 8605 1730 8615 1750
rect 8635 1730 8645 1750
rect 8605 1715 8645 1730
rect 8660 1750 8700 1765
rect 8660 1730 8670 1750
rect 8690 1730 8700 1750
rect 8660 1715 8700 1730
rect 8715 1750 8755 1765
rect 8715 1730 8725 1750
rect 8745 1730 8755 1750
rect 8715 1715 8755 1730
rect 8915 1750 8955 1765
rect 8915 1730 8925 1750
rect 8945 1730 8955 1750
rect 8915 1715 8955 1730
rect 8970 1750 9010 1765
rect 8970 1730 8980 1750
rect 9000 1730 9010 1750
rect 8970 1715 9010 1730
rect 9085 1750 9125 1765
rect 9085 1730 9095 1750
rect 9115 1730 9125 1750
rect 9085 1715 9125 1730
rect 9140 1750 9180 1765
rect 9140 1730 9150 1750
rect 9170 1730 9180 1750
rect 9140 1715 9180 1730
rect 9195 1750 9235 1765
rect 9195 1730 9205 1750
rect 9225 1730 9235 1750
rect 9195 1715 9235 1730
rect 9265 1750 9305 1765
rect 9265 1730 9275 1750
rect 9295 1730 9305 1750
rect 9265 1715 9305 1730
rect 9320 1750 9360 1765
rect 9320 1730 9330 1750
rect 9350 1730 9360 1750
rect 9320 1715 9360 1730
rect 9375 1750 9415 1765
rect 9375 1730 9385 1750
rect 9405 1730 9415 1750
rect 9375 1715 9415 1730
rect 9565 1750 9605 1765
rect 9565 1730 9575 1750
rect 9595 1730 9605 1750
rect 9565 1715 9605 1730
rect 9620 1750 9660 1765
rect 9620 1730 9630 1750
rect 9650 1730 9660 1750
rect 9620 1715 9660 1730
rect 9735 1750 9775 1765
rect 9735 1730 9745 1750
rect 9765 1730 9775 1750
rect 9735 1715 9775 1730
rect 9790 1750 9830 1765
rect 9790 1730 9800 1750
rect 9820 1730 9830 1750
rect 9790 1715 9830 1730
rect 9845 1750 9885 1765
rect 9845 1730 9855 1750
rect 9875 1730 9885 1750
rect 9845 1715 9885 1730
rect 9915 1750 9955 1765
rect 9915 1730 9925 1750
rect 9945 1730 9955 1750
rect 9915 1715 9955 1730
rect 9970 1750 10010 1765
rect 9970 1730 9980 1750
rect 10000 1730 10010 1750
rect 9970 1715 10010 1730
rect 10025 1750 10065 1765
rect 10025 1730 10035 1750
rect 10055 1730 10065 1750
rect 10025 1715 10065 1730
rect 10215 1750 10255 1765
rect 10215 1730 10225 1750
rect 10245 1730 10255 1750
rect 10215 1715 10255 1730
rect 10270 1750 10310 1765
rect 10270 1730 10280 1750
rect 10300 1730 10310 1750
rect 10270 1715 10310 1730
rect 10385 1750 10425 1765
rect 10385 1730 10395 1750
rect 10415 1730 10425 1750
rect 10385 1715 10425 1730
rect 10440 1750 10480 1765
rect 10440 1730 10450 1750
rect 10470 1730 10480 1750
rect 10440 1715 10480 1730
rect 10495 1750 10535 1765
rect 10495 1730 10505 1750
rect 10525 1730 10535 1750
rect 10495 1715 10535 1730
rect 10565 1750 10605 1765
rect 10565 1730 10575 1750
rect 10595 1730 10605 1750
rect 10565 1715 10605 1730
rect 10620 1750 10660 1765
rect 10620 1730 10630 1750
rect 10650 1730 10660 1750
rect 10620 1715 10660 1730
rect 10675 1750 10715 1765
rect 10675 1730 10685 1750
rect 10705 1730 10715 1750
rect 10675 1715 10715 1730
rect 10865 1750 10905 1765
rect 10865 1730 10875 1750
rect 10895 1730 10905 1750
rect 10865 1715 10905 1730
rect 10920 1750 10960 1765
rect 10920 1730 10930 1750
rect 10950 1730 10960 1750
rect 10920 1715 10960 1730
rect 11035 1750 11075 1765
rect 11035 1730 11045 1750
rect 11065 1730 11075 1750
rect 11035 1715 11075 1730
rect 11090 1750 11130 1765
rect 11090 1730 11100 1750
rect 11120 1730 11130 1750
rect 11090 1715 11130 1730
rect 11145 1750 11185 1765
rect 11145 1730 11155 1750
rect 11175 1730 11185 1750
rect 11145 1715 11185 1730
rect 11215 1750 11255 1765
rect 11215 1730 11225 1750
rect 11245 1730 11255 1750
rect 11215 1715 11255 1730
rect 11270 1750 11310 1765
rect 11270 1730 11280 1750
rect 11300 1730 11310 1750
rect 11270 1715 11310 1730
rect 11325 1750 11365 1765
rect 11325 1730 11335 1750
rect 11355 1730 11365 1750
rect 11325 1715 11365 1730
<< ndiffc >>
rect 6205 1570 6225 1590
rect 6260 1570 6280 1590
rect 6315 1570 6335 1590
rect 6370 1570 6390 1590
rect 6425 1570 6445 1590
rect 6495 1570 6515 1590
rect 6550 1570 6570 1590
rect 6605 1570 6625 1590
rect 6720 1570 6740 1590
rect 6775 1570 6795 1590
rect 6830 1570 6850 1590
rect 6885 1570 6905 1590
rect 6940 1570 6960 1590
rect 7050 1570 7070 1590
rect 7105 1570 7125 1590
rect 7160 1570 7180 1590
rect 7215 1570 7235 1590
rect 7270 1570 7290 1590
rect 7410 1570 7430 1590
rect 7465 1570 7485 1590
rect 7520 1570 7540 1590
rect 7575 1570 7595 1590
rect 7630 1570 7650 1590
rect 7700 1570 7720 1590
rect 7755 1570 7775 1590
rect 7810 1570 7830 1590
rect 7980 1570 8000 1590
rect 8035 1570 8055 1590
rect 8160 1570 8180 1590
rect 8215 1570 8235 1590
rect 8285 1570 8305 1590
rect 8340 1570 8360 1590
rect 8395 1570 8415 1590
rect 8450 1570 8470 1590
rect 8505 1570 8525 1590
rect 8615 1570 8635 1590
rect 8670 1570 8690 1590
rect 8725 1570 8745 1590
rect 8780 1570 8800 1590
rect 8890 1570 8910 1590
rect 8945 1570 8965 1590
rect 9000 1570 9020 1590
rect 9055 1570 9075 1590
rect 9110 1570 9130 1590
rect 9220 1570 9240 1590
rect 9275 1570 9295 1590
rect 9330 1570 9350 1590
rect 9385 1570 9405 1590
rect 9540 1525 9560 1545
rect 9595 1525 9615 1545
rect 9650 1525 9670 1545
rect 9705 1525 9725 1545
rect 9760 1525 9780 1545
rect 9870 1525 9890 1545
rect 9925 1525 9945 1545
rect 9980 1525 10000 1545
rect 10035 1525 10055 1545
rect 10190 1525 10210 1545
rect 10245 1525 10265 1545
rect 10300 1525 10320 1545
rect 10355 1525 10375 1545
rect 10410 1525 10430 1545
rect 10520 1525 10540 1545
rect 10575 1525 10595 1545
rect 10630 1525 10650 1545
rect 10685 1525 10705 1545
rect 10840 1525 10860 1545
rect 10895 1525 10915 1545
rect 10950 1525 10970 1545
rect 11005 1525 11025 1545
rect 11060 1525 11080 1545
rect 11170 1525 11190 1545
rect 11225 1525 11245 1545
rect 11280 1525 11300 1545
rect 11335 1525 11355 1545
<< pdiffc >>
rect 6285 1730 6305 1750
rect 6340 1730 6360 1750
rect 6495 1730 6515 1750
rect 6550 1730 6570 1750
rect 6605 1730 6625 1750
rect 6830 1730 6850 1750
rect 6885 1730 6905 1750
rect 6940 1730 6960 1750
rect 7050 1730 7070 1750
rect 7105 1730 7125 1750
rect 7160 1730 7180 1750
rect 7215 1730 7235 1750
rect 7490 1730 7510 1750
rect 7545 1730 7565 1750
rect 7700 1730 7720 1750
rect 7755 1730 7775 1750
rect 7810 1730 7830 1750
rect 7925 1730 7945 1750
rect 7980 1730 8000 1750
rect 8035 1730 8055 1750
rect 8105 1730 8125 1750
rect 8160 1730 8180 1750
rect 8215 1730 8235 1750
rect 8395 1730 8415 1750
rect 8450 1730 8470 1750
rect 8505 1730 8525 1750
rect 8615 1730 8635 1750
rect 8670 1730 8690 1750
rect 8725 1730 8745 1750
rect 8925 1730 8945 1750
rect 8980 1730 9000 1750
rect 9095 1730 9115 1750
rect 9150 1730 9170 1750
rect 9205 1730 9225 1750
rect 9275 1730 9295 1750
rect 9330 1730 9350 1750
rect 9385 1730 9405 1750
rect 9575 1730 9595 1750
rect 9630 1730 9650 1750
rect 9745 1730 9765 1750
rect 9800 1730 9820 1750
rect 9855 1730 9875 1750
rect 9925 1730 9945 1750
rect 9980 1730 10000 1750
rect 10035 1730 10055 1750
rect 10225 1730 10245 1750
rect 10280 1730 10300 1750
rect 10395 1730 10415 1750
rect 10450 1730 10470 1750
rect 10505 1730 10525 1750
rect 10575 1730 10595 1750
rect 10630 1730 10650 1750
rect 10685 1730 10705 1750
rect 10875 1730 10895 1750
rect 10930 1730 10950 1750
rect 11045 1730 11065 1750
rect 11100 1730 11120 1750
rect 11155 1730 11175 1750
rect 11225 1730 11245 1750
rect 11280 1730 11300 1750
rect 11335 1730 11355 1750
<< psubdiff >>
rect 7330 1545 7370 1560
rect 7840 1590 7880 1605
rect 7840 1570 7850 1590
rect 7870 1570 7880 1590
rect 7840 1555 7880 1570
rect 8565 1590 8605 1605
rect 8565 1570 8575 1590
rect 8595 1570 8605 1590
rect 8565 1555 8605 1570
rect 7330 1525 7340 1545
rect 7360 1525 7370 1545
rect 9460 1545 9500 1560
rect 7330 1510 7370 1525
rect 9460 1525 9470 1545
rect 9490 1525 9500 1545
rect 9460 1510 9500 1525
rect 10110 1545 10150 1560
rect 10110 1525 10120 1545
rect 10140 1525 10150 1545
rect 10110 1510 10150 1525
rect 10760 1545 10800 1560
rect 10760 1525 10770 1545
rect 10790 1525 10800 1545
rect 10760 1510 10800 1525
<< nsubdiff >>
rect 6370 1750 6410 1765
rect 6370 1730 6380 1750
rect 6400 1730 6410 1750
rect 6370 1715 6410 1730
rect 7575 1750 7615 1765
rect 7575 1730 7585 1750
rect 7605 1730 7615 1750
rect 7575 1715 7615 1730
rect 9010 1750 9050 1765
rect 9010 1730 9020 1750
rect 9040 1730 9050 1750
rect 9010 1715 9050 1730
rect 9660 1750 9700 1765
rect 9660 1730 9670 1750
rect 9690 1730 9700 1750
rect 9660 1715 9700 1730
rect 10310 1750 10350 1765
rect 10310 1730 10320 1750
rect 10340 1730 10350 1750
rect 10310 1715 10350 1730
rect 10960 1750 11000 1765
rect 10960 1730 10970 1750
rect 10990 1730 11000 1750
rect 10960 1715 11000 1730
<< psubdiffcont >>
rect 7850 1570 7870 1590
rect 8575 1570 8595 1590
rect 7340 1525 7360 1545
rect 9470 1525 9490 1545
rect 10120 1525 10140 1545
rect 10770 1525 10790 1545
<< nsubdiffcont >>
rect 6380 1730 6400 1750
rect 7585 1730 7605 1750
rect 9020 1730 9040 1750
rect 9670 1730 9690 1750
rect 10320 1730 10340 1750
rect 10970 1730 10990 1750
<< poly >>
rect 6490 1810 6540 1820
rect 7050 1810 7095 1820
rect 6490 1790 6500 1810
rect 6520 1790 6540 1810
rect 6490 1780 6540 1790
rect 6645 1800 6685 1810
rect 6645 1780 6655 1800
rect 6675 1780 6685 1800
rect 7050 1790 7060 1810
rect 7080 1790 7095 1810
rect 7050 1780 7095 1790
rect 7120 1810 7150 1820
rect 7120 1790 7125 1810
rect 7145 1790 7150 1810
rect 7120 1780 7150 1790
rect 7700 1810 7745 1820
rect 7700 1790 7710 1810
rect 7730 1790 7745 1810
rect 7700 1780 7745 1790
rect 8580 1815 8620 1820
rect 8580 1795 8590 1815
rect 8610 1800 8620 1815
rect 9830 1810 9885 1820
rect 8610 1795 8660 1800
rect 8580 1785 8660 1795
rect 9830 1790 9855 1810
rect 9875 1790 9885 1810
rect 10480 1810 10535 1820
rect 10480 1790 10505 1810
rect 10525 1790 10535 1810
rect 11130 1810 11185 1820
rect 11130 1790 11155 1810
rect 11175 1790 11185 1810
rect 6315 1765 6330 1780
rect 6525 1765 6540 1780
rect 6580 1765 6595 1780
rect 6645 1770 6685 1780
rect 6150 1750 6190 1760
rect 6150 1730 6160 1750
rect 6180 1730 6190 1750
rect 6150 1720 6190 1730
rect 6225 1650 6265 1660
rect 6225 1630 6235 1650
rect 6255 1630 6265 1650
rect 6315 1630 6330 1715
rect 6525 1700 6540 1715
rect 6580 1685 6595 1715
rect 6645 1685 6660 1770
rect 6860 1765 6875 1780
rect 6915 1765 6930 1780
rect 7080 1765 7095 1780
rect 7135 1765 7150 1780
rect 7190 1765 7205 1780
rect 7520 1765 7535 1780
rect 7730 1765 7745 1780
rect 7785 1765 7800 1780
rect 7955 1765 7970 1780
rect 8010 1765 8025 1780
rect 8135 1765 8150 1780
rect 8190 1765 8205 1780
rect 8425 1765 8440 1780
rect 8480 1765 8495 1780
rect 8645 1765 8660 1785
rect 8700 1765 8715 1780
rect 8955 1765 8970 1780
rect 9125 1765 9140 1780
rect 9180 1765 9195 1780
rect 9305 1775 9375 1790
rect 9830 1780 9885 1790
rect 9305 1765 9320 1775
rect 9360 1765 9375 1775
rect 9605 1765 9620 1780
rect 9775 1765 9790 1780
rect 9830 1765 9845 1780
rect 9955 1775 10025 1790
rect 10480 1780 10535 1790
rect 9955 1765 9970 1775
rect 10010 1765 10025 1775
rect 10255 1765 10270 1780
rect 10425 1765 10440 1780
rect 10480 1765 10495 1780
rect 10605 1775 10675 1790
rect 11130 1780 11185 1790
rect 10605 1765 10620 1775
rect 10660 1765 10675 1775
rect 10905 1765 10920 1780
rect 11075 1765 11090 1780
rect 11130 1765 11145 1780
rect 11255 1775 11325 1790
rect 11255 1765 11270 1775
rect 11310 1765 11325 1775
rect 6580 1670 6660 1685
rect 6785 1690 6825 1700
rect 6785 1675 6795 1690
rect 6515 1650 6555 1660
rect 6515 1630 6525 1650
rect 6545 1630 6555 1650
rect 6225 1620 6265 1630
rect 6290 1620 6555 1630
rect 6235 1605 6250 1620
rect 6290 1615 6540 1620
rect 6290 1605 6305 1615
rect 6345 1605 6360 1615
rect 6400 1605 6415 1615
rect 6525 1605 6540 1615
rect 6580 1605 6595 1670
rect 6235 1540 6250 1555
rect 6290 1540 6305 1555
rect 6345 1540 6360 1555
rect 6400 1540 6415 1555
rect 6525 1540 6540 1555
rect 6580 1540 6595 1555
rect 6645 1550 6660 1670
rect 6750 1670 6795 1675
rect 6815 1670 6825 1690
rect 6750 1660 6825 1670
rect 6685 1650 6725 1660
rect 6685 1630 6695 1650
rect 6715 1630 6725 1650
rect 6685 1620 6725 1630
rect 6750 1605 6765 1660
rect 6860 1635 6875 1715
rect 6915 1700 6930 1715
rect 6985 1710 7025 1720
rect 6985 1700 6995 1710
rect 6915 1690 6995 1700
rect 7015 1690 7025 1710
rect 6915 1685 7025 1690
rect 6985 1680 7025 1685
rect 6975 1650 7015 1655
rect 6975 1635 6985 1650
rect 6805 1630 6985 1635
rect 7005 1630 7015 1650
rect 6805 1620 7015 1630
rect 6805 1605 6820 1620
rect 6860 1605 6875 1620
rect 6915 1605 6930 1620
rect 7080 1605 7095 1715
rect 7135 1605 7150 1715
rect 7190 1605 7205 1715
rect 7520 1695 7535 1715
rect 7730 1700 7745 1715
rect 7355 1680 7535 1695
rect 7235 1650 7275 1655
rect 7235 1630 7245 1650
rect 7265 1635 7275 1650
rect 7355 1635 7370 1680
rect 7265 1630 7370 1635
rect 7235 1620 7370 1630
rect 7430 1650 7470 1655
rect 7430 1630 7440 1650
rect 7460 1630 7470 1650
rect 7520 1630 7535 1680
rect 7785 1695 7800 1715
rect 7855 1710 7895 1720
rect 7855 1695 7865 1710
rect 7785 1690 7865 1695
rect 7885 1690 7895 1710
rect 7955 1705 7970 1715
rect 8010 1705 8025 1715
rect 7955 1690 8025 1705
rect 8135 1705 8150 1715
rect 8190 1705 8205 1715
rect 8135 1690 8205 1705
rect 7785 1680 7895 1690
rect 7720 1650 7760 1660
rect 7720 1630 7730 1650
rect 7750 1630 7760 1650
rect 7430 1620 7470 1630
rect 7495 1620 7760 1630
rect 7245 1605 7260 1620
rect 7440 1605 7455 1620
rect 7495 1615 7745 1620
rect 7495 1605 7510 1615
rect 7550 1605 7565 1615
rect 7605 1605 7620 1615
rect 7730 1605 7745 1615
rect 7785 1605 7800 1680
rect 7825 1650 7865 1655
rect 7945 1650 7985 1660
rect 7825 1630 7835 1650
rect 7855 1635 7955 1650
rect 7855 1630 7865 1635
rect 7825 1620 7865 1630
rect 7945 1630 7955 1635
rect 7975 1630 7985 1650
rect 7945 1620 7985 1630
rect 8010 1605 8025 1690
rect 8190 1670 8205 1690
rect 8350 1690 8390 1700
rect 8250 1675 8290 1685
rect 8350 1675 8360 1690
rect 8250 1670 8260 1675
rect 8115 1655 8155 1665
rect 8115 1635 8125 1655
rect 8145 1635 8155 1655
rect 8115 1625 8155 1635
rect 8190 1655 8260 1670
rect 8280 1655 8290 1675
rect 8190 1605 8205 1655
rect 8250 1645 8290 1655
rect 8315 1670 8360 1675
rect 8380 1670 8390 1690
rect 8315 1660 8390 1670
rect 8315 1605 8330 1660
rect 8425 1635 8440 1715
rect 8480 1700 8495 1715
rect 8550 1710 8590 1720
rect 8845 1750 8885 1760
rect 8845 1735 8855 1750
rect 8765 1730 8855 1735
rect 8875 1730 8885 1750
rect 8765 1720 8885 1730
rect 8550 1700 8560 1710
rect 8480 1690 8560 1700
rect 8580 1690 8590 1710
rect 8480 1685 8590 1690
rect 8550 1680 8590 1685
rect 8565 1650 8605 1655
rect 8565 1635 8575 1650
rect 8370 1630 8575 1635
rect 8595 1630 8605 1650
rect 8370 1620 8605 1630
rect 8370 1605 8385 1620
rect 8425 1605 8440 1620
rect 8480 1605 8495 1620
rect 8645 1605 8660 1715
rect 8700 1695 8715 1715
rect 8765 1695 8780 1720
rect 8955 1695 8970 1715
rect 9125 1700 9140 1715
rect 9180 1705 9195 1715
rect 8700 1680 8780 1695
rect 8835 1680 8990 1695
rect 8700 1605 8715 1680
rect 8745 1650 8785 1655
rect 8745 1630 8755 1650
rect 8775 1635 8785 1650
rect 8835 1635 8850 1680
rect 8775 1630 8850 1635
rect 8745 1620 8850 1630
rect 8910 1650 8950 1655
rect 8910 1630 8920 1650
rect 8940 1630 8950 1650
rect 8910 1620 8950 1630
rect 8975 1630 8990 1680
rect 9115 1690 9155 1700
rect 9180 1690 9280 1705
rect 9305 1700 9320 1715
rect 9115 1670 9125 1690
rect 9145 1670 9155 1690
rect 9115 1660 9155 1670
rect 9265 1675 9280 1690
rect 9265 1660 9320 1675
rect 9200 1650 9240 1660
rect 9200 1630 9210 1650
rect 9230 1630 9240 1650
rect 8755 1605 8770 1620
rect 8920 1605 8935 1620
rect 8975 1615 9265 1630
rect 8975 1605 8990 1615
rect 9030 1605 9045 1615
rect 9085 1605 9100 1615
rect 9250 1605 9265 1615
rect 9305 1605 9320 1660
rect 9360 1660 9375 1715
rect 9605 1700 9620 1715
rect 9775 1700 9790 1715
rect 9605 1685 9640 1700
rect 9435 1660 9475 1670
rect 9360 1645 9445 1660
rect 9360 1605 9375 1645
rect 9435 1640 9445 1645
rect 9465 1640 9475 1660
rect 9435 1630 9475 1640
rect 9560 1605 9600 1615
rect 6645 1540 6685 1550
rect 6750 1540 6765 1555
rect 6805 1540 6820 1555
rect 6860 1540 6875 1555
rect 6915 1540 6930 1555
rect 7080 1540 7095 1555
rect 7135 1540 7150 1555
rect 7190 1540 7205 1555
rect 7245 1540 7260 1555
rect 9560 1585 9570 1605
rect 9590 1585 9600 1605
rect 9560 1575 9600 1585
rect 9625 1585 9640 1685
rect 9765 1690 9805 1700
rect 9765 1670 9775 1690
rect 9795 1670 9805 1690
rect 9765 1660 9805 1670
rect 9830 1660 9845 1715
rect 9955 1700 9970 1715
rect 10010 1660 10025 1715
rect 10255 1700 10270 1715
rect 10425 1700 10440 1715
rect 10255 1685 10290 1700
rect 10085 1660 10125 1670
rect 9830 1645 9970 1660
rect 9850 1605 9890 1615
rect 9850 1585 9860 1605
rect 9880 1585 9890 1605
rect 9570 1560 9585 1575
rect 9625 1570 9915 1585
rect 9625 1560 9640 1570
rect 9680 1560 9695 1570
rect 9735 1560 9750 1570
rect 9900 1560 9915 1570
rect 9955 1560 9970 1645
rect 10010 1645 10095 1660
rect 10010 1560 10025 1645
rect 10085 1640 10095 1645
rect 10115 1640 10125 1660
rect 10085 1630 10125 1640
rect 10210 1605 10250 1615
rect 10210 1585 10220 1605
rect 10240 1585 10250 1605
rect 10210 1575 10250 1585
rect 10275 1585 10290 1685
rect 10415 1690 10455 1700
rect 10415 1670 10425 1690
rect 10445 1670 10455 1690
rect 10415 1660 10455 1670
rect 10480 1660 10495 1715
rect 10605 1700 10620 1715
rect 10660 1660 10675 1715
rect 10905 1700 10920 1715
rect 11075 1700 11090 1715
rect 10905 1685 10940 1700
rect 10735 1660 10775 1670
rect 10480 1645 10620 1660
rect 10500 1605 10540 1615
rect 10500 1585 10510 1605
rect 10530 1585 10540 1605
rect 10220 1560 10235 1575
rect 10275 1570 10565 1585
rect 10275 1560 10290 1570
rect 10330 1560 10345 1570
rect 10385 1560 10400 1570
rect 10550 1560 10565 1570
rect 10605 1560 10620 1645
rect 10660 1645 10745 1660
rect 10660 1560 10675 1645
rect 10735 1640 10745 1645
rect 10765 1640 10775 1660
rect 10735 1630 10775 1640
rect 10860 1605 10900 1615
rect 10860 1585 10870 1605
rect 10890 1585 10900 1605
rect 10860 1575 10900 1585
rect 10925 1585 10940 1685
rect 11065 1690 11105 1700
rect 11065 1670 11075 1690
rect 11095 1670 11105 1690
rect 11065 1660 11105 1670
rect 11130 1660 11145 1715
rect 11255 1700 11270 1715
rect 11310 1660 11325 1715
rect 11376 1661 11405 1670
rect 11376 1660 11382 1661
rect 11130 1645 11270 1660
rect 11150 1605 11190 1615
rect 11150 1585 11160 1605
rect 11180 1585 11190 1605
rect 10870 1560 10885 1575
rect 10925 1570 11215 1585
rect 10925 1560 10940 1570
rect 10980 1560 10995 1570
rect 11035 1560 11050 1570
rect 11200 1560 11215 1570
rect 11255 1560 11270 1645
rect 11310 1645 11382 1660
rect 11310 1560 11325 1645
rect 11376 1644 11382 1645
rect 11399 1644 11405 1661
rect 11376 1630 11405 1644
rect 6150 1530 6190 1540
rect 6150 1510 6160 1530
rect 6180 1510 6190 1530
rect 6645 1520 6655 1540
rect 6675 1520 6685 1540
rect 6645 1510 6685 1520
rect 7180 1535 7220 1540
rect 7180 1515 7190 1535
rect 7210 1515 7220 1535
rect 6150 1500 6190 1510
rect 7180 1505 7220 1515
rect 7440 1540 7455 1555
rect 7495 1540 7510 1555
rect 7550 1540 7565 1555
rect 7605 1540 7620 1555
rect 7730 1540 7745 1555
rect 7785 1540 7800 1555
rect 8010 1540 8025 1555
rect 8190 1540 8205 1555
rect 8315 1540 8330 1555
rect 8370 1540 8385 1555
rect 8425 1540 8440 1555
rect 8480 1540 8495 1555
rect 8645 1540 8660 1555
rect 8700 1540 8715 1555
rect 8755 1540 8770 1555
rect 8920 1540 8935 1555
rect 8975 1540 8990 1555
rect 9030 1540 9045 1555
rect 9085 1540 9100 1555
rect 9250 1540 9265 1555
rect 9305 1540 9320 1555
rect 9360 1540 9375 1555
rect 7980 1535 8025 1540
rect 7980 1515 7990 1535
rect 8010 1515 8025 1535
rect 7980 1505 8025 1515
rect 9287 1530 9320 1540
rect 9287 1510 9292 1530
rect 9312 1510 9320 1530
rect 9287 1500 9320 1510
rect 9570 1495 9585 1510
rect 9625 1495 9640 1510
rect 9680 1495 9695 1510
rect 9735 1495 9750 1510
rect 9900 1495 9915 1510
rect 9955 1495 9970 1510
rect 10010 1495 10025 1510
rect 10220 1495 10235 1510
rect 10275 1495 10290 1510
rect 10330 1495 10345 1510
rect 10385 1495 10400 1510
rect 10550 1495 10565 1510
rect 10605 1495 10620 1510
rect 10660 1495 10675 1510
rect 10870 1495 10885 1510
rect 10925 1495 10940 1510
rect 10980 1495 10995 1510
rect 11035 1495 11050 1510
rect 11200 1495 11215 1510
rect 11255 1495 11270 1510
rect 11310 1495 11325 1510
<< polycont >>
rect 6500 1790 6520 1810
rect 6655 1780 6675 1800
rect 7060 1790 7080 1810
rect 7125 1790 7145 1810
rect 7710 1790 7730 1810
rect 8590 1795 8610 1815
rect 9855 1790 9875 1810
rect 10505 1790 10525 1810
rect 11155 1790 11175 1810
rect 6160 1730 6180 1750
rect 6235 1630 6255 1650
rect 6525 1630 6545 1650
rect 6795 1670 6815 1690
rect 6695 1630 6715 1650
rect 6995 1690 7015 1710
rect 6985 1630 7005 1650
rect 7245 1630 7265 1650
rect 7440 1630 7460 1650
rect 7865 1690 7885 1710
rect 7730 1630 7750 1650
rect 7835 1630 7855 1650
rect 7955 1630 7975 1650
rect 8125 1635 8145 1655
rect 8260 1655 8280 1675
rect 8360 1670 8380 1690
rect 8855 1730 8875 1750
rect 8560 1690 8580 1710
rect 8575 1630 8595 1650
rect 8755 1630 8775 1650
rect 8920 1630 8940 1650
rect 9125 1670 9145 1690
rect 9210 1630 9230 1650
rect 9445 1640 9465 1660
rect 9570 1585 9590 1605
rect 9775 1670 9795 1690
rect 9860 1585 9880 1605
rect 10095 1640 10115 1660
rect 10220 1585 10240 1605
rect 10425 1670 10445 1690
rect 10510 1585 10530 1605
rect 10745 1640 10765 1660
rect 10870 1585 10890 1605
rect 11075 1670 11095 1690
rect 11160 1585 11180 1605
rect 11382 1644 11399 1661
rect 6160 1510 6180 1530
rect 6655 1520 6675 1540
rect 7190 1515 7210 1535
rect 7990 1515 8010 1535
rect 9292 1510 9312 1530
<< locali >>
rect 6330 1865 6370 1875
rect 6330 1845 6340 1865
rect 6360 1845 6370 1865
rect 6330 1835 6370 1845
rect 6540 1865 6580 1875
rect 6540 1845 6550 1865
rect 6570 1845 6580 1865
rect 6540 1835 6580 1845
rect 6875 1865 6915 1875
rect 6875 1845 6885 1865
rect 6905 1845 6915 1865
rect 6875 1835 6915 1845
rect 7160 1865 7200 1875
rect 7160 1845 7170 1865
rect 7190 1845 7200 1865
rect 7160 1835 7200 1845
rect 7535 1865 7575 1875
rect 7535 1845 7545 1865
rect 7565 1845 7575 1865
rect 7535 1835 7575 1845
rect 7750 1865 7790 1875
rect 7750 1845 7760 1865
rect 7780 1845 7790 1865
rect 7750 1835 7790 1845
rect 7970 1865 8010 1875
rect 7970 1845 7980 1865
rect 8000 1845 8010 1865
rect 7970 1835 8010 1845
rect 8095 1865 8135 1875
rect 8095 1845 8105 1865
rect 8125 1845 8135 1865
rect 8095 1835 8135 1845
rect 8205 1865 8245 1875
rect 8205 1845 8215 1865
rect 8235 1845 8245 1865
rect 8205 1835 8245 1845
rect 8440 1865 8480 1875
rect 8440 1845 8450 1865
rect 8470 1845 8480 1865
rect 8440 1835 8480 1845
rect 8660 1865 8700 1875
rect 8660 1845 8670 1865
rect 8690 1845 8700 1865
rect 8660 1835 8700 1845
rect 8970 1865 9010 1875
rect 8970 1845 8980 1865
rect 9000 1845 9010 1865
rect 8970 1835 9010 1845
rect 9140 1865 9180 1875
rect 9140 1845 9150 1865
rect 9170 1845 9180 1865
rect 9140 1835 9180 1845
rect 9320 1865 9360 1875
rect 9320 1845 9330 1865
rect 9350 1845 9360 1865
rect 9320 1835 9360 1845
rect 9620 1865 9660 1875
rect 9620 1845 9630 1865
rect 9650 1845 9660 1865
rect 9620 1835 9660 1845
rect 9790 1865 9830 1875
rect 9790 1845 9800 1865
rect 9820 1845 9830 1865
rect 9790 1835 9830 1845
rect 9970 1865 10010 1875
rect 9970 1845 9980 1865
rect 10000 1845 10010 1865
rect 9970 1835 10010 1845
rect 10270 1865 10310 1875
rect 10270 1845 10280 1865
rect 10300 1845 10310 1865
rect 10270 1835 10310 1845
rect 10440 1865 10480 1875
rect 10440 1845 10450 1865
rect 10470 1845 10480 1865
rect 10440 1835 10480 1845
rect 10620 1865 10660 1875
rect 10620 1845 10630 1865
rect 10650 1845 10660 1865
rect 10620 1835 10660 1845
rect 10920 1865 10960 1875
rect 10920 1845 10930 1865
rect 10950 1845 10960 1865
rect 10920 1835 10960 1845
rect 11090 1865 11130 1875
rect 11090 1845 11100 1865
rect 11120 1845 11130 1865
rect 11090 1835 11130 1845
rect 11270 1865 11310 1875
rect 11270 1845 11280 1865
rect 11300 1845 11310 1865
rect 11270 1835 11310 1845
rect 6340 1760 6360 1835
rect 6490 1810 6530 1820
rect 6490 1790 6500 1810
rect 6520 1790 6530 1810
rect 6490 1780 6530 1790
rect 6550 1760 6570 1835
rect 6590 1810 6625 1820
rect 6590 1790 6595 1810
rect 6615 1790 6625 1810
rect 6590 1780 6625 1790
rect 6605 1760 6625 1780
rect 6645 1800 6685 1810
rect 6645 1780 6655 1800
rect 6675 1780 6685 1800
rect 6645 1770 6685 1780
rect 6885 1760 6905 1835
rect 7050 1810 7090 1820
rect 7050 1790 7060 1810
rect 7080 1790 7090 1810
rect 7050 1780 7090 1790
rect 7120 1810 7150 1820
rect 7120 1790 7125 1810
rect 7145 1790 7150 1810
rect 7120 1780 7150 1790
rect 7170 1760 7190 1835
rect 7545 1760 7565 1835
rect 7700 1810 7740 1820
rect 7700 1790 7710 1810
rect 7730 1790 7740 1810
rect 7700 1780 7740 1790
rect 7760 1760 7780 1835
rect 7810 1810 7850 1820
rect 7810 1790 7820 1810
rect 7840 1790 7850 1810
rect 7810 1780 7850 1790
rect 7810 1760 7830 1780
rect 7980 1760 8000 1835
rect 8105 1760 8125 1835
rect 8215 1760 8235 1835
rect 8375 1815 8415 1820
rect 8375 1795 8385 1815
rect 8405 1795 8415 1815
rect 8375 1785 8415 1795
rect 8395 1760 8415 1785
rect 8450 1760 8470 1835
rect 8580 1815 8620 1820
rect 8580 1795 8590 1815
rect 8610 1795 8620 1815
rect 8580 1785 8620 1795
rect 8670 1760 8690 1835
rect 8980 1760 9000 1835
rect 9150 1760 9170 1835
rect 9330 1760 9350 1835
rect 9555 1810 9595 1820
rect 9555 1790 9565 1810
rect 9585 1790 9595 1810
rect 9555 1780 9595 1790
rect 9575 1760 9595 1780
rect 9630 1760 9650 1835
rect 9800 1760 9820 1835
rect 9845 1810 9885 1820
rect 9845 1790 9855 1810
rect 9875 1790 9885 1810
rect 9845 1780 9885 1790
rect 9980 1760 10000 1835
rect 10205 1810 10245 1820
rect 10205 1790 10215 1810
rect 10235 1790 10245 1810
rect 10205 1780 10245 1790
rect 10225 1760 10245 1780
rect 10280 1760 10300 1835
rect 10450 1760 10470 1835
rect 10495 1810 10535 1820
rect 10495 1790 10505 1810
rect 10525 1790 10535 1810
rect 10495 1780 10535 1790
rect 10630 1760 10650 1835
rect 10855 1810 10895 1820
rect 10855 1790 10865 1810
rect 10885 1790 10895 1810
rect 10855 1780 10895 1790
rect 10875 1760 10895 1780
rect 10930 1760 10950 1835
rect 11100 1760 11120 1835
rect 11145 1810 11185 1820
rect 11145 1790 11155 1810
rect 11175 1790 11185 1810
rect 11145 1780 11185 1790
rect 11280 1760 11300 1835
rect 6150 1750 6190 1760
rect 6280 1750 6310 1760
rect 6150 1730 6160 1750
rect 6180 1730 6285 1750
rect 6305 1730 6310 1750
rect 6150 1720 6190 1730
rect 6280 1720 6310 1730
rect 6335 1750 6405 1760
rect 6490 1750 6520 1760
rect 6335 1730 6340 1750
rect 6360 1730 6380 1750
rect 6400 1730 6405 1750
rect 6335 1720 6405 1730
rect 6425 1730 6495 1750
rect 6515 1730 6520 1750
rect 6160 1675 6180 1720
rect 6120 1665 6180 1675
rect 6120 1645 6130 1665
rect 6150 1645 6180 1665
rect 6120 1635 6180 1645
rect 6160 1540 6180 1635
rect 6225 1650 6265 1660
rect 6225 1630 6235 1650
rect 6255 1640 6265 1650
rect 6425 1640 6445 1730
rect 6490 1720 6520 1730
rect 6545 1750 6575 1760
rect 6545 1730 6550 1750
rect 6570 1730 6575 1750
rect 6545 1720 6575 1730
rect 6600 1750 6630 1760
rect 6825 1750 6855 1760
rect 6600 1730 6605 1750
rect 6625 1730 6630 1750
rect 6600 1720 6630 1730
rect 6715 1730 6830 1750
rect 6850 1730 6855 1750
rect 6605 1700 6625 1720
rect 6255 1630 6445 1640
rect 6225 1620 6445 1630
rect 6315 1600 6335 1620
rect 6425 1600 6445 1620
rect 6470 1680 6625 1700
rect 6470 1600 6490 1680
rect 6715 1660 6735 1730
rect 6825 1720 6855 1730
rect 6880 1750 6910 1760
rect 6880 1730 6885 1750
rect 6905 1730 6910 1750
rect 6880 1720 6910 1730
rect 6935 1750 6965 1760
rect 6935 1730 6940 1750
rect 6960 1730 6965 1750
rect 6935 1720 6965 1730
rect 7045 1750 7075 1760
rect 7045 1730 7050 1750
rect 7070 1730 7075 1750
rect 7045 1720 7075 1730
rect 7100 1750 7130 1760
rect 7100 1730 7105 1750
rect 7125 1730 7130 1750
rect 7100 1720 7130 1730
rect 7155 1750 7190 1760
rect 7155 1730 7160 1750
rect 7180 1730 7190 1750
rect 7155 1720 7190 1730
rect 7210 1750 7240 1760
rect 7210 1730 7215 1750
rect 7235 1730 7240 1750
rect 7210 1720 7240 1730
rect 7365 1750 7405 1760
rect 7485 1750 7515 1760
rect 7365 1730 7375 1750
rect 7395 1730 7490 1750
rect 7510 1730 7515 1750
rect 7365 1720 7405 1730
rect 7485 1720 7515 1730
rect 7540 1750 7610 1760
rect 7695 1750 7725 1760
rect 7540 1730 7545 1750
rect 7565 1730 7585 1750
rect 7605 1730 7610 1750
rect 7540 1720 7610 1730
rect 7630 1730 7700 1750
rect 7720 1730 7725 1750
rect 6785 1690 6825 1700
rect 6785 1670 6795 1690
rect 6815 1670 6825 1690
rect 6785 1660 6825 1670
rect 6515 1650 6555 1660
rect 6685 1650 6735 1660
rect 6515 1630 6525 1650
rect 6545 1630 6695 1650
rect 6715 1630 6735 1650
rect 6515 1620 6555 1630
rect 6685 1620 6735 1630
rect 6805 1640 6825 1660
rect 6935 1640 6955 1720
rect 6985 1710 7025 1720
rect 6985 1690 6995 1710
rect 7015 1700 7025 1710
rect 7050 1700 7070 1720
rect 7215 1700 7235 1720
rect 7015 1690 7315 1700
rect 6985 1680 7315 1690
rect 6805 1620 6955 1640
rect 6975 1650 7015 1655
rect 6975 1630 6985 1650
rect 7005 1630 7015 1650
rect 7235 1650 7275 1655
rect 6975 1620 7015 1630
rect 7050 1620 7180 1640
rect 7235 1630 7245 1650
rect 7265 1630 7275 1650
rect 7235 1620 7275 1630
rect 6715 1600 6735 1620
rect 6825 1600 6845 1620
rect 6935 1600 6955 1620
rect 7050 1600 7070 1620
rect 7160 1600 7180 1620
rect 7295 1600 7315 1680
rect 6200 1590 6230 1600
rect 6200 1570 6205 1590
rect 6225 1570 6230 1590
rect 6200 1560 6230 1570
rect 6255 1590 6285 1600
rect 6255 1570 6260 1590
rect 6280 1570 6285 1590
rect 6255 1560 6285 1570
rect 6310 1590 6340 1600
rect 6310 1570 6315 1590
rect 6335 1570 6340 1590
rect 6310 1560 6340 1570
rect 6365 1590 6395 1600
rect 6365 1570 6370 1590
rect 6390 1570 6395 1590
rect 6365 1560 6395 1570
rect 6420 1590 6450 1600
rect 6420 1570 6425 1590
rect 6445 1570 6450 1590
rect 6470 1590 6520 1600
rect 6470 1570 6495 1590
rect 6515 1570 6520 1590
rect 6420 1560 6450 1570
rect 6490 1560 6520 1570
rect 6545 1590 6575 1600
rect 6545 1570 6550 1590
rect 6570 1570 6575 1590
rect 6545 1560 6575 1570
rect 6600 1590 6630 1600
rect 6600 1570 6605 1590
rect 6625 1570 6630 1590
rect 6600 1560 6630 1570
rect 6715 1590 6745 1600
rect 6715 1570 6720 1590
rect 6740 1570 6745 1590
rect 6715 1560 6745 1570
rect 6770 1590 6800 1600
rect 6770 1570 6775 1590
rect 6795 1570 6800 1590
rect 6770 1560 6800 1570
rect 6825 1590 6855 1600
rect 6825 1570 6830 1590
rect 6850 1570 6855 1590
rect 6825 1560 6855 1570
rect 6880 1590 6910 1600
rect 6880 1570 6885 1590
rect 6905 1570 6910 1590
rect 6880 1560 6910 1570
rect 6935 1590 6965 1600
rect 6935 1570 6940 1590
rect 6960 1570 6965 1590
rect 6935 1560 6965 1570
rect 7045 1590 7075 1600
rect 7045 1570 7050 1590
rect 7070 1570 7075 1590
rect 7045 1560 7075 1570
rect 7100 1590 7130 1600
rect 7100 1570 7105 1590
rect 7125 1570 7130 1590
rect 7100 1560 7130 1570
rect 7155 1590 7185 1600
rect 7155 1570 7160 1590
rect 7180 1570 7185 1590
rect 7155 1560 7185 1570
rect 7210 1590 7240 1600
rect 7210 1570 7215 1590
rect 7235 1570 7240 1590
rect 7210 1560 7240 1570
rect 7265 1590 7315 1600
rect 7265 1570 7270 1590
rect 7290 1570 7315 1590
rect 7385 1600 7405 1720
rect 7430 1650 7470 1655
rect 7430 1630 7440 1650
rect 7460 1640 7470 1650
rect 7630 1640 7650 1730
rect 7695 1720 7725 1730
rect 7750 1750 7780 1760
rect 7750 1730 7755 1750
rect 7775 1730 7780 1750
rect 7750 1720 7780 1730
rect 7805 1750 7835 1760
rect 7805 1730 7810 1750
rect 7830 1730 7835 1750
rect 7805 1720 7835 1730
rect 7920 1750 7950 1760
rect 7920 1730 7925 1750
rect 7945 1730 7950 1750
rect 7920 1720 7950 1730
rect 7975 1750 8005 1760
rect 7975 1730 7980 1750
rect 8000 1730 8005 1750
rect 7975 1720 8005 1730
rect 8030 1750 8060 1760
rect 8030 1730 8035 1750
rect 8055 1730 8060 1750
rect 8030 1720 8060 1730
rect 8100 1750 8130 1760
rect 8100 1730 8105 1750
rect 8125 1730 8130 1750
rect 8100 1720 8130 1730
rect 8155 1750 8185 1760
rect 8155 1730 8160 1750
rect 8180 1730 8185 1750
rect 8155 1720 8185 1730
rect 8210 1750 8240 1760
rect 8390 1750 8420 1760
rect 8210 1730 8215 1750
rect 8235 1730 8240 1750
rect 8210 1720 8240 1730
rect 8280 1730 8395 1750
rect 8415 1730 8420 1750
rect 7810 1700 7830 1720
rect 7460 1630 7650 1640
rect 7430 1620 7650 1630
rect 7520 1600 7540 1620
rect 7630 1600 7650 1620
rect 7675 1680 7830 1700
rect 7855 1710 7895 1720
rect 7855 1690 7865 1710
rect 7885 1700 7895 1710
rect 7925 1700 7945 1720
rect 8035 1700 8055 1720
rect 7885 1690 8055 1700
rect 7855 1680 8055 1690
rect 7675 1600 7695 1680
rect 7720 1650 7760 1660
rect 7825 1650 7865 1655
rect 7720 1630 7730 1650
rect 7750 1630 7835 1650
rect 7855 1630 7865 1650
rect 7720 1620 7760 1630
rect 7825 1620 7865 1630
rect 7385 1590 7435 1600
rect 7385 1570 7410 1590
rect 7430 1570 7435 1590
rect 7265 1560 7295 1570
rect 7405 1560 7435 1570
rect 7460 1590 7490 1600
rect 7460 1570 7465 1590
rect 7485 1570 7490 1590
rect 7460 1560 7490 1570
rect 7515 1590 7545 1600
rect 7515 1570 7520 1590
rect 7540 1570 7545 1590
rect 7515 1560 7545 1570
rect 7570 1590 7600 1600
rect 7570 1570 7575 1590
rect 7595 1570 7600 1590
rect 7570 1560 7600 1570
rect 7625 1590 7655 1600
rect 7625 1570 7630 1590
rect 7650 1570 7655 1590
rect 7675 1590 7725 1600
rect 7675 1570 7700 1590
rect 7720 1570 7725 1590
rect 7625 1560 7655 1570
rect 7695 1560 7725 1570
rect 7750 1590 7780 1600
rect 7750 1570 7755 1590
rect 7775 1570 7780 1590
rect 7750 1560 7780 1570
rect 7805 1590 7875 1600
rect 7805 1570 7810 1590
rect 7830 1570 7850 1590
rect 7870 1570 7875 1590
rect 7895 1590 7915 1680
rect 8160 1665 8180 1720
rect 8280 1685 8300 1730
rect 8390 1720 8420 1730
rect 8445 1750 8475 1760
rect 8445 1730 8450 1750
rect 8470 1730 8475 1750
rect 8445 1720 8475 1730
rect 8500 1750 8530 1760
rect 8500 1730 8505 1750
rect 8525 1730 8530 1750
rect 8500 1720 8530 1730
rect 8610 1750 8640 1760
rect 8610 1730 8615 1750
rect 8635 1730 8640 1750
rect 8610 1720 8640 1730
rect 8665 1750 8695 1760
rect 8665 1730 8670 1750
rect 8690 1730 8695 1750
rect 8665 1720 8695 1730
rect 8720 1750 8750 1760
rect 8845 1750 8885 1760
rect 8920 1750 8950 1760
rect 8720 1730 8725 1750
rect 8745 1730 8825 1750
rect 8720 1720 8750 1730
rect 8115 1660 8180 1665
rect 7945 1655 8180 1660
rect 7945 1650 8125 1655
rect 7945 1630 7955 1650
rect 7975 1640 8125 1650
rect 7975 1630 7985 1640
rect 7945 1620 7985 1630
rect 8115 1635 8125 1640
rect 8145 1635 8180 1655
rect 8250 1675 8300 1685
rect 8250 1655 8260 1675
rect 8280 1655 8300 1675
rect 8350 1690 8390 1700
rect 8350 1670 8360 1690
rect 8380 1670 8390 1690
rect 8350 1660 8390 1670
rect 8250 1645 8300 1655
rect 8115 1625 8180 1635
rect 8160 1600 8180 1625
rect 8280 1600 8300 1645
rect 8370 1640 8390 1660
rect 8500 1640 8520 1720
rect 8550 1710 8590 1720
rect 8550 1690 8560 1710
rect 8580 1700 8590 1710
rect 8615 1700 8635 1720
rect 8725 1700 8745 1720
rect 8580 1690 8745 1700
rect 8550 1680 8745 1690
rect 8370 1620 8520 1640
rect 8565 1650 8605 1655
rect 8745 1650 8785 1655
rect 8565 1630 8575 1650
rect 8595 1630 8755 1650
rect 8775 1630 8785 1650
rect 8565 1620 8605 1630
rect 8745 1620 8785 1630
rect 8390 1600 8410 1620
rect 8500 1600 8520 1620
rect 8805 1600 8825 1730
rect 8845 1730 8855 1750
rect 8875 1730 8925 1750
rect 8945 1730 8950 1750
rect 8845 1720 8885 1730
rect 8920 1720 8950 1730
rect 8975 1750 9045 1760
rect 8975 1730 8980 1750
rect 9000 1730 9020 1750
rect 9040 1730 9045 1750
rect 8975 1720 9045 1730
rect 9075 1750 9120 1760
rect 9075 1730 9095 1750
rect 9115 1730 9120 1750
rect 9075 1720 9120 1730
rect 9145 1750 9175 1760
rect 9145 1730 9150 1750
rect 9170 1730 9175 1750
rect 9145 1720 9175 1730
rect 9200 1750 9230 1760
rect 9200 1730 9205 1750
rect 9225 1730 9230 1750
rect 9200 1720 9230 1730
rect 9270 1750 9300 1760
rect 9270 1730 9275 1750
rect 9295 1730 9300 1750
rect 9270 1720 9300 1730
rect 9325 1750 9355 1760
rect 9325 1730 9330 1750
rect 9350 1730 9355 1750
rect 9325 1720 9355 1730
rect 9380 1750 9410 1760
rect 9570 1750 9600 1760
rect 9380 1730 9385 1750
rect 9405 1730 9410 1750
rect 9380 1720 9410 1730
rect 9515 1730 9575 1750
rect 9595 1730 9600 1750
rect 7975 1590 8005 1600
rect 7895 1570 7980 1590
rect 8000 1570 8005 1590
rect 7805 1560 7875 1570
rect 7975 1560 8005 1570
rect 8030 1590 8060 1600
rect 8030 1570 8035 1590
rect 8055 1570 8060 1590
rect 8030 1560 8060 1570
rect 8155 1590 8185 1600
rect 8155 1570 8160 1590
rect 8180 1570 8185 1590
rect 8155 1560 8185 1570
rect 8210 1590 8240 1600
rect 8210 1570 8215 1590
rect 8235 1570 8240 1590
rect 8210 1560 8240 1570
rect 8280 1590 8310 1600
rect 8280 1570 8285 1590
rect 8305 1570 8310 1590
rect 8280 1560 8310 1570
rect 8335 1590 8365 1600
rect 8335 1570 8340 1590
rect 8360 1570 8365 1590
rect 8335 1560 8365 1570
rect 8390 1590 8420 1600
rect 8390 1570 8395 1590
rect 8415 1570 8420 1590
rect 8390 1560 8420 1570
rect 8445 1590 8475 1600
rect 8445 1570 8450 1590
rect 8470 1570 8475 1590
rect 8445 1560 8475 1570
rect 8500 1590 8530 1600
rect 8500 1570 8505 1590
rect 8525 1570 8530 1590
rect 8500 1560 8530 1570
rect 8570 1590 8640 1600
rect 8570 1570 8575 1590
rect 8595 1570 8615 1590
rect 8635 1570 8640 1590
rect 8570 1560 8640 1570
rect 8665 1590 8695 1600
rect 8665 1570 8670 1590
rect 8690 1570 8695 1590
rect 8665 1560 8695 1570
rect 8720 1590 8750 1600
rect 8720 1570 8725 1590
rect 8745 1570 8750 1590
rect 8720 1560 8750 1570
rect 8775 1590 8825 1600
rect 8775 1570 8780 1590
rect 8800 1570 8825 1590
rect 8865 1600 8885 1720
rect 8910 1650 8950 1655
rect 8910 1630 8920 1650
rect 8940 1640 8950 1650
rect 9075 1640 9095 1720
rect 9205 1700 9225 1720
rect 9115 1690 9225 1700
rect 9115 1670 9125 1690
rect 9145 1680 9225 1690
rect 9145 1670 9175 1680
rect 9115 1660 9175 1670
rect 8940 1630 9130 1640
rect 8910 1620 9130 1630
rect 9000 1600 9020 1620
rect 9110 1600 9130 1620
rect 9155 1600 9175 1660
rect 9200 1650 9240 1660
rect 9200 1630 9210 1650
rect 9230 1640 9240 1650
rect 9275 1640 9295 1720
rect 9385 1640 9405 1720
rect 9515 1670 9535 1730
rect 9570 1720 9600 1730
rect 9625 1750 9695 1760
rect 9625 1730 9630 1750
rect 9650 1730 9670 1750
rect 9690 1730 9695 1750
rect 9625 1720 9695 1730
rect 9725 1750 9770 1760
rect 9725 1730 9745 1750
rect 9765 1730 9770 1750
rect 9725 1720 9770 1730
rect 9795 1750 9825 1760
rect 9795 1730 9800 1750
rect 9820 1730 9825 1750
rect 9795 1720 9825 1730
rect 9850 1750 9880 1760
rect 9850 1730 9855 1750
rect 9875 1730 9880 1750
rect 9850 1720 9880 1730
rect 9920 1750 9950 1760
rect 9920 1730 9925 1750
rect 9945 1730 9950 1750
rect 9920 1720 9950 1730
rect 9975 1750 10005 1760
rect 9975 1730 9980 1750
rect 10000 1730 10005 1750
rect 9975 1720 10005 1730
rect 10030 1750 10060 1760
rect 10220 1750 10250 1760
rect 10030 1730 10035 1750
rect 10055 1730 10060 1750
rect 10030 1720 10060 1730
rect 10165 1730 10225 1750
rect 10245 1730 10250 1750
rect 9230 1630 9405 1640
rect 9435 1660 9535 1670
rect 9435 1640 9445 1660
rect 9465 1650 9535 1660
rect 9465 1640 9475 1650
rect 9435 1630 9475 1640
rect 9200 1620 9405 1630
rect 9385 1600 9405 1620
rect 8865 1590 8915 1600
rect 8865 1570 8890 1590
rect 8910 1570 8915 1590
rect 8775 1560 8805 1570
rect 8885 1560 8915 1570
rect 8940 1590 8970 1600
rect 8940 1570 8945 1590
rect 8965 1570 8970 1590
rect 8940 1560 8970 1570
rect 8995 1590 9025 1600
rect 8995 1570 9000 1590
rect 9020 1570 9025 1590
rect 8995 1560 9025 1570
rect 9050 1590 9080 1600
rect 9050 1570 9055 1590
rect 9075 1570 9080 1590
rect 9050 1560 9080 1570
rect 9105 1590 9135 1600
rect 9105 1570 9110 1590
rect 9130 1570 9135 1590
rect 9155 1590 9245 1600
rect 9155 1580 9220 1590
rect 9105 1560 9135 1570
rect 9215 1570 9220 1580
rect 9240 1570 9245 1590
rect 9215 1560 9245 1570
rect 9270 1590 9300 1600
rect 9270 1570 9275 1590
rect 9295 1570 9300 1590
rect 9270 1560 9300 1570
rect 9325 1590 9360 1600
rect 9325 1570 9330 1590
rect 9350 1570 9360 1590
rect 9325 1560 9360 1570
rect 9380 1590 9410 1600
rect 9380 1570 9385 1590
rect 9405 1570 9410 1590
rect 9380 1560 9410 1570
rect 6150 1530 6190 1540
rect 6150 1510 6160 1530
rect 6180 1510 6190 1530
rect 6150 1500 6190 1510
rect 6260 1485 6280 1560
rect 6370 1485 6390 1560
rect 6605 1485 6625 1560
rect 6645 1540 6685 1550
rect 6720 1540 6740 1560
rect 6645 1520 6655 1540
rect 6675 1520 6685 1540
rect 6645 1510 6685 1520
rect 6710 1535 6750 1540
rect 6710 1515 6720 1535
rect 6740 1515 6750 1535
rect 6710 1505 6750 1515
rect 6775 1485 6795 1560
rect 6885 1485 6905 1560
rect 7105 1485 7125 1560
rect 7335 1545 7365 1555
rect 7180 1535 7220 1540
rect 7180 1515 7190 1535
rect 7210 1515 7220 1535
rect 7335 1525 7340 1545
rect 7360 1525 7365 1545
rect 7335 1515 7365 1525
rect 7180 1505 7220 1515
rect 7340 1485 7360 1515
rect 7465 1485 7485 1560
rect 7575 1485 7595 1560
rect 7810 1485 7830 1560
rect 7980 1535 8020 1540
rect 7980 1515 7990 1535
rect 8010 1515 8020 1535
rect 7980 1505 8020 1515
rect 8040 1485 8060 1560
rect 8215 1485 8235 1560
rect 8340 1485 8360 1560
rect 8450 1485 8470 1560
rect 8615 1485 8635 1560
rect 8945 1485 8965 1560
rect 9055 1485 9075 1560
rect 9287 1530 9320 1540
rect 9287 1510 9292 1530
rect 9312 1510 9320 1530
rect 9287 1500 9320 1510
rect 9340 1485 9360 1560
rect 9515 1555 9535 1650
rect 9560 1605 9600 1615
rect 9560 1585 9570 1605
rect 9590 1595 9600 1605
rect 9725 1595 9745 1720
rect 9855 1700 9875 1720
rect 9765 1690 9875 1700
rect 9765 1670 9775 1690
rect 9795 1680 9875 1690
rect 9795 1670 9825 1680
rect 9765 1660 9825 1670
rect 9590 1585 9780 1595
rect 9560 1575 9780 1585
rect 9650 1555 9670 1575
rect 9760 1555 9780 1575
rect 9805 1555 9825 1660
rect 9850 1605 9890 1615
rect 9850 1585 9860 1605
rect 9880 1595 9890 1605
rect 9925 1595 9945 1720
rect 10035 1595 10055 1720
rect 10165 1670 10185 1730
rect 10220 1720 10250 1730
rect 10275 1750 10345 1760
rect 10275 1730 10280 1750
rect 10300 1730 10320 1750
rect 10340 1730 10345 1750
rect 10275 1720 10345 1730
rect 10375 1750 10420 1760
rect 10375 1730 10395 1750
rect 10415 1730 10420 1750
rect 10375 1720 10420 1730
rect 10445 1750 10475 1760
rect 10445 1730 10450 1750
rect 10470 1730 10475 1750
rect 10445 1720 10475 1730
rect 10500 1750 10530 1760
rect 10500 1730 10505 1750
rect 10525 1730 10530 1750
rect 10500 1720 10530 1730
rect 10570 1750 10600 1760
rect 10570 1730 10575 1750
rect 10595 1730 10600 1750
rect 10570 1720 10600 1730
rect 10625 1750 10655 1760
rect 10625 1730 10630 1750
rect 10650 1730 10655 1750
rect 10625 1720 10655 1730
rect 10680 1750 10710 1760
rect 10870 1750 10900 1760
rect 10680 1730 10685 1750
rect 10705 1730 10710 1750
rect 10680 1720 10710 1730
rect 10815 1730 10875 1750
rect 10895 1730 10900 1750
rect 10085 1660 10185 1670
rect 10085 1640 10095 1660
rect 10115 1650 10185 1660
rect 10115 1640 10125 1650
rect 10085 1630 10125 1640
rect 9880 1585 10055 1595
rect 9850 1575 10055 1585
rect 10035 1555 10055 1575
rect 10165 1555 10185 1650
rect 10210 1605 10250 1615
rect 10210 1585 10220 1605
rect 10240 1595 10250 1605
rect 10375 1595 10395 1720
rect 10505 1700 10525 1720
rect 10415 1690 10525 1700
rect 10415 1670 10425 1690
rect 10445 1680 10525 1690
rect 10445 1670 10475 1680
rect 10415 1660 10475 1670
rect 10240 1585 10430 1595
rect 10210 1575 10430 1585
rect 10300 1555 10320 1575
rect 10410 1555 10430 1575
rect 10455 1555 10475 1660
rect 10500 1605 10540 1615
rect 10500 1585 10510 1605
rect 10530 1595 10540 1605
rect 10575 1595 10595 1720
rect 10685 1595 10705 1720
rect 10815 1670 10835 1730
rect 10870 1720 10900 1730
rect 10925 1750 10995 1760
rect 10925 1730 10930 1750
rect 10950 1730 10970 1750
rect 10990 1730 10995 1750
rect 10925 1720 10995 1730
rect 11025 1750 11070 1760
rect 11025 1730 11045 1750
rect 11065 1730 11070 1750
rect 11025 1720 11070 1730
rect 11095 1750 11125 1760
rect 11095 1730 11100 1750
rect 11120 1730 11125 1750
rect 11095 1720 11125 1730
rect 11150 1750 11180 1760
rect 11150 1730 11155 1750
rect 11175 1730 11180 1750
rect 11150 1720 11180 1730
rect 11220 1750 11250 1760
rect 11220 1730 11225 1750
rect 11245 1730 11250 1750
rect 11220 1720 11250 1730
rect 11275 1750 11305 1760
rect 11275 1730 11280 1750
rect 11300 1730 11305 1750
rect 11275 1720 11305 1730
rect 11330 1750 11360 1760
rect 11330 1730 11335 1750
rect 11355 1730 11360 1750
rect 11330 1720 11360 1730
rect 10735 1660 10835 1670
rect 10735 1640 10745 1660
rect 10765 1650 10835 1660
rect 10765 1640 10775 1650
rect 10735 1630 10775 1640
rect 10530 1585 10705 1595
rect 10500 1575 10705 1585
rect 10685 1555 10705 1575
rect 10815 1555 10835 1650
rect 10860 1605 10900 1615
rect 10860 1585 10870 1605
rect 10890 1595 10900 1605
rect 11025 1595 11045 1720
rect 11155 1700 11175 1720
rect 11065 1690 11175 1700
rect 11065 1670 11075 1690
rect 11095 1680 11175 1690
rect 11095 1670 11125 1680
rect 11065 1660 11125 1670
rect 10890 1585 11080 1595
rect 10860 1575 11080 1585
rect 10950 1555 10970 1575
rect 11060 1555 11080 1575
rect 11105 1555 11125 1660
rect 11150 1605 11190 1615
rect 11150 1585 11160 1605
rect 11180 1595 11190 1605
rect 11225 1595 11245 1720
rect 11335 1595 11355 1720
rect 11376 1661 11405 1670
rect 11376 1644 11382 1661
rect 11399 1644 11405 1661
rect 11376 1630 11405 1644
rect 11180 1585 11355 1595
rect 11150 1575 11355 1585
rect 11335 1555 11355 1575
rect 9465 1545 9495 1555
rect 9465 1525 9470 1545
rect 9490 1525 9495 1545
rect 9515 1545 9565 1555
rect 9515 1525 9540 1545
rect 9560 1525 9565 1545
rect 9465 1515 9495 1525
rect 9535 1515 9565 1525
rect 9590 1545 9620 1555
rect 9590 1525 9595 1545
rect 9615 1525 9620 1545
rect 9590 1515 9620 1525
rect 9645 1545 9675 1555
rect 9645 1525 9650 1545
rect 9670 1525 9675 1545
rect 9645 1515 9675 1525
rect 9700 1545 9730 1555
rect 9700 1525 9705 1545
rect 9725 1525 9730 1545
rect 9700 1515 9730 1525
rect 9755 1545 9785 1555
rect 9755 1525 9760 1545
rect 9780 1525 9785 1545
rect 9805 1545 9895 1555
rect 9805 1535 9870 1545
rect 9755 1515 9785 1525
rect 9865 1525 9870 1535
rect 9890 1525 9895 1545
rect 9865 1515 9895 1525
rect 9920 1545 9950 1555
rect 9920 1525 9925 1545
rect 9945 1525 9950 1545
rect 9920 1515 9950 1525
rect 9975 1545 10005 1555
rect 9975 1525 9980 1545
rect 10000 1525 10005 1545
rect 9975 1515 10005 1525
rect 10030 1545 10060 1555
rect 10030 1525 10035 1545
rect 10055 1525 10060 1545
rect 10030 1515 10060 1525
rect 10115 1545 10145 1555
rect 10115 1525 10120 1545
rect 10140 1525 10145 1545
rect 10165 1545 10215 1555
rect 10165 1525 10190 1545
rect 10210 1525 10215 1545
rect 10115 1515 10145 1525
rect 10185 1515 10215 1525
rect 10240 1545 10270 1555
rect 10240 1525 10245 1545
rect 10265 1525 10270 1545
rect 10240 1515 10270 1525
rect 10295 1545 10325 1555
rect 10295 1525 10300 1545
rect 10320 1525 10325 1545
rect 10295 1515 10325 1525
rect 10350 1545 10380 1555
rect 10350 1525 10355 1545
rect 10375 1525 10380 1545
rect 10350 1515 10380 1525
rect 10405 1545 10435 1555
rect 10405 1525 10410 1545
rect 10430 1525 10435 1545
rect 10455 1545 10545 1555
rect 10455 1535 10520 1545
rect 10405 1515 10435 1525
rect 10515 1525 10520 1535
rect 10540 1525 10545 1545
rect 10515 1515 10545 1525
rect 10570 1545 10600 1555
rect 10570 1525 10575 1545
rect 10595 1525 10600 1545
rect 10570 1515 10600 1525
rect 10625 1545 10655 1555
rect 10625 1525 10630 1545
rect 10650 1525 10655 1545
rect 10625 1515 10655 1525
rect 10680 1545 10710 1555
rect 10680 1525 10685 1545
rect 10705 1525 10710 1545
rect 10680 1515 10710 1525
rect 10765 1545 10795 1555
rect 10765 1525 10770 1545
rect 10790 1525 10795 1545
rect 10815 1545 10865 1555
rect 10815 1525 10840 1545
rect 10860 1525 10865 1545
rect 10765 1515 10795 1525
rect 10835 1515 10865 1525
rect 10890 1545 10920 1555
rect 10890 1525 10895 1545
rect 10915 1525 10920 1545
rect 10890 1515 10920 1525
rect 10945 1545 10975 1555
rect 10945 1525 10950 1545
rect 10970 1525 10975 1545
rect 10945 1515 10975 1525
rect 11000 1545 11030 1555
rect 11000 1525 11005 1545
rect 11025 1525 11030 1545
rect 11000 1515 11030 1525
rect 11055 1545 11085 1555
rect 11055 1525 11060 1545
rect 11080 1525 11085 1545
rect 11105 1545 11195 1555
rect 11105 1535 11170 1545
rect 11055 1515 11085 1525
rect 11165 1525 11170 1535
rect 11190 1525 11195 1545
rect 11165 1515 11195 1525
rect 11220 1545 11250 1555
rect 11220 1525 11225 1545
rect 11245 1525 11250 1545
rect 11220 1515 11250 1525
rect 11275 1545 11305 1555
rect 11275 1525 11280 1545
rect 11300 1525 11305 1545
rect 11275 1515 11305 1525
rect 11330 1545 11360 1555
rect 11330 1525 11335 1545
rect 11355 1525 11360 1545
rect 11330 1515 11360 1525
rect 9470 1485 9490 1515
rect 9595 1485 9615 1515
rect 9705 1485 9725 1515
rect 9980 1485 10000 1515
rect 10120 1485 10140 1515
rect 10245 1485 10265 1515
rect 10355 1485 10375 1515
rect 10630 1485 10650 1515
rect 10770 1485 10790 1515
rect 10895 1485 10915 1515
rect 11005 1485 11025 1515
rect 11280 1485 11300 1515
rect 6250 1475 6290 1485
rect 6250 1455 6260 1475
rect 6280 1455 6290 1475
rect 6250 1445 6290 1455
rect 6360 1475 6400 1485
rect 6360 1455 6370 1475
rect 6390 1455 6400 1475
rect 6360 1445 6400 1455
rect 6595 1475 6635 1485
rect 6595 1455 6605 1475
rect 6625 1455 6635 1475
rect 6595 1445 6635 1455
rect 6765 1475 6805 1485
rect 6765 1455 6775 1475
rect 6795 1455 6805 1475
rect 6765 1445 6805 1455
rect 6875 1475 6915 1485
rect 6875 1455 6885 1475
rect 6905 1455 6915 1475
rect 6875 1445 6915 1455
rect 7095 1475 7135 1485
rect 7095 1455 7105 1475
rect 7125 1455 7135 1475
rect 7095 1445 7135 1455
rect 7330 1475 7370 1485
rect 7330 1455 7340 1475
rect 7360 1455 7370 1475
rect 7330 1445 7370 1455
rect 7455 1475 7495 1485
rect 7455 1455 7465 1475
rect 7485 1455 7495 1475
rect 7455 1445 7495 1455
rect 7565 1475 7605 1485
rect 7565 1455 7575 1475
rect 7595 1455 7605 1475
rect 7565 1445 7605 1455
rect 7800 1475 7840 1485
rect 7800 1455 7810 1475
rect 7830 1455 7840 1475
rect 7800 1445 7840 1455
rect 8030 1475 8070 1485
rect 8030 1455 8040 1475
rect 8060 1455 8070 1475
rect 8030 1445 8070 1455
rect 8205 1475 8245 1485
rect 8205 1455 8215 1475
rect 8235 1455 8245 1475
rect 8205 1445 8245 1455
rect 8330 1475 8370 1485
rect 8330 1455 8340 1475
rect 8360 1455 8370 1475
rect 8330 1445 8370 1455
rect 8440 1475 8480 1485
rect 8440 1455 8450 1475
rect 8470 1455 8480 1475
rect 8440 1445 8480 1455
rect 8605 1475 8645 1485
rect 8605 1455 8615 1475
rect 8635 1455 8645 1475
rect 8605 1445 8645 1455
rect 8935 1475 8975 1485
rect 8935 1455 8945 1475
rect 8965 1455 8975 1475
rect 8935 1445 8975 1455
rect 9045 1475 9085 1485
rect 9045 1455 9055 1475
rect 9075 1455 9085 1475
rect 9045 1445 9085 1455
rect 9330 1475 9370 1485
rect 9330 1455 9340 1475
rect 9360 1455 9370 1475
rect 9330 1445 9370 1455
rect 9460 1475 9500 1485
rect 9460 1455 9470 1475
rect 9490 1455 9500 1475
rect 9460 1445 9500 1455
rect 9585 1475 9625 1485
rect 9585 1455 9595 1475
rect 9615 1455 9625 1475
rect 9585 1445 9625 1455
rect 9695 1475 9735 1485
rect 9695 1455 9705 1475
rect 9725 1455 9735 1475
rect 9695 1445 9735 1455
rect 9970 1475 10010 1485
rect 9970 1455 9980 1475
rect 10000 1455 10010 1475
rect 9970 1445 10010 1455
rect 10110 1475 10150 1485
rect 10110 1455 10120 1475
rect 10140 1455 10150 1475
rect 10110 1445 10150 1455
rect 10235 1475 10275 1485
rect 10235 1455 10245 1475
rect 10265 1455 10275 1475
rect 10235 1445 10275 1455
rect 10345 1475 10385 1485
rect 10345 1455 10355 1475
rect 10375 1455 10385 1475
rect 10345 1445 10385 1455
rect 10620 1475 10660 1485
rect 10620 1455 10630 1475
rect 10650 1455 10660 1475
rect 10620 1445 10660 1455
rect 10760 1475 10800 1485
rect 10760 1455 10770 1475
rect 10790 1455 10800 1475
rect 10760 1445 10800 1455
rect 10885 1475 10925 1485
rect 10885 1455 10895 1475
rect 10915 1455 10925 1475
rect 10885 1445 10925 1455
rect 10995 1475 11035 1485
rect 10995 1455 11005 1475
rect 11025 1455 11035 1475
rect 10995 1445 11035 1455
rect 11270 1475 11310 1485
rect 11270 1455 11280 1475
rect 11300 1455 11310 1475
rect 11270 1445 11310 1455
<< viali >>
rect 6340 1845 6360 1865
rect 6550 1845 6570 1865
rect 6885 1845 6905 1865
rect 7170 1845 7190 1865
rect 7545 1845 7565 1865
rect 7760 1845 7780 1865
rect 7980 1845 8000 1865
rect 8105 1845 8125 1865
rect 8215 1845 8235 1865
rect 8450 1845 8470 1865
rect 8670 1845 8690 1865
rect 8980 1845 9000 1865
rect 9150 1845 9170 1865
rect 9330 1845 9350 1865
rect 9630 1845 9650 1865
rect 9800 1845 9820 1865
rect 9980 1845 10000 1865
rect 10280 1845 10300 1865
rect 10450 1845 10470 1865
rect 10630 1845 10650 1865
rect 10930 1845 10950 1865
rect 11100 1845 11120 1865
rect 11280 1845 11300 1865
rect 6500 1790 6520 1810
rect 6595 1790 6615 1810
rect 6655 1780 6675 1800
rect 7060 1790 7080 1810
rect 7125 1790 7145 1810
rect 7710 1790 7730 1810
rect 7820 1790 7840 1810
rect 8385 1795 8405 1815
rect 8590 1795 8610 1815
rect 9565 1790 9585 1810
rect 9855 1790 9875 1810
rect 10215 1790 10235 1810
rect 10505 1790 10525 1810
rect 10865 1790 10885 1810
rect 11155 1790 11175 1810
rect 6130 1645 6150 1665
rect 7375 1730 7395 1750
rect 6985 1630 7005 1650
rect 7245 1630 7265 1650
rect 8125 1635 8145 1655
rect 6160 1510 6180 1530
rect 6655 1520 6675 1540
rect 6720 1515 6740 1535
rect 7190 1515 7210 1535
rect 7990 1515 8010 1535
rect 9292 1510 9312 1530
rect 11382 1644 11399 1661
rect 6260 1455 6280 1475
rect 6370 1455 6390 1475
rect 6605 1455 6625 1475
rect 6775 1455 6795 1475
rect 6885 1455 6905 1475
rect 7105 1455 7125 1475
rect 7340 1455 7360 1475
rect 7465 1455 7485 1475
rect 7575 1455 7595 1475
rect 7810 1455 7830 1475
rect 8040 1455 8060 1475
rect 8215 1455 8235 1475
rect 8340 1455 8360 1475
rect 8450 1455 8470 1475
rect 8615 1455 8635 1475
rect 8945 1455 8965 1475
rect 9055 1455 9075 1475
rect 9340 1455 9360 1475
rect 9470 1455 9490 1475
rect 9595 1455 9615 1475
rect 9705 1455 9725 1475
rect 9980 1455 10000 1475
rect 10120 1455 10140 1475
rect 10245 1455 10265 1475
rect 10355 1455 10375 1475
rect 10630 1455 10650 1475
rect 10770 1455 10790 1475
rect 10895 1455 10915 1475
rect 11005 1455 11025 1475
rect 11280 1455 11300 1475
<< metal1 >>
rect 6330 1870 6370 1875
rect 6330 1840 6335 1870
rect 6365 1840 6370 1870
rect 6330 1835 6370 1840
rect 6540 1870 6580 1875
rect 6540 1840 6545 1870
rect 6575 1840 6580 1870
rect 6540 1835 6580 1840
rect 6875 1870 6915 1875
rect 6875 1840 6880 1870
rect 6910 1840 6915 1870
rect 6875 1835 6915 1840
rect 7160 1870 7200 1875
rect 7160 1840 7165 1870
rect 7195 1840 7200 1870
rect 7160 1835 7200 1840
rect 7535 1870 7575 1875
rect 7535 1840 7540 1870
rect 7570 1840 7575 1870
rect 7535 1835 7575 1840
rect 7750 1870 7790 1875
rect 7750 1840 7755 1870
rect 7785 1840 7790 1870
rect 7750 1835 7790 1840
rect 7970 1870 8010 1875
rect 7970 1840 7975 1870
rect 8005 1840 8010 1870
rect 7970 1835 8010 1840
rect 8095 1870 8135 1875
rect 8095 1840 8100 1870
rect 8130 1840 8135 1870
rect 8095 1835 8135 1840
rect 8205 1870 8245 1875
rect 8205 1840 8210 1870
rect 8240 1840 8245 1870
rect 8205 1835 8245 1840
rect 8440 1870 8480 1875
rect 8440 1840 8445 1870
rect 8475 1840 8480 1870
rect 8440 1835 8480 1840
rect 8660 1870 8700 1875
rect 8660 1840 8665 1870
rect 8695 1840 8700 1870
rect 8660 1835 8700 1840
rect 8970 1870 9010 1875
rect 8970 1840 8975 1870
rect 9005 1840 9010 1870
rect 8970 1835 9010 1840
rect 9140 1870 9180 1875
rect 9140 1840 9145 1870
rect 9175 1840 9180 1870
rect 9140 1835 9180 1840
rect 9320 1870 9360 1875
rect 9320 1840 9325 1870
rect 9355 1840 9360 1870
rect 9320 1835 9360 1840
rect 9620 1870 9660 1875
rect 9620 1840 9625 1870
rect 9655 1840 9660 1870
rect 9620 1835 9660 1840
rect 9790 1870 9830 1875
rect 9790 1840 9795 1870
rect 9825 1840 9830 1870
rect 9790 1835 9830 1840
rect 9970 1870 10010 1875
rect 9970 1840 9975 1870
rect 10005 1840 10010 1870
rect 9970 1835 10010 1840
rect 10270 1870 10310 1875
rect 10270 1840 10275 1870
rect 10305 1840 10310 1870
rect 10270 1835 10310 1840
rect 10440 1870 10480 1875
rect 10440 1840 10445 1870
rect 10475 1840 10480 1870
rect 10440 1835 10480 1840
rect 10620 1870 10660 1875
rect 10620 1840 10625 1870
rect 10655 1840 10660 1870
rect 10620 1835 10660 1840
rect 10920 1870 10960 1875
rect 10920 1840 10925 1870
rect 10955 1840 10960 1870
rect 10920 1835 10960 1840
rect 11090 1870 11130 1875
rect 11090 1840 11095 1870
rect 11125 1840 11130 1870
rect 11090 1835 11130 1840
rect 11270 1870 11310 1875
rect 11270 1840 11275 1870
rect 11305 1840 11310 1870
rect 11270 1835 11310 1840
rect 6490 1810 6530 1820
rect 6490 1790 6500 1810
rect 6520 1800 6530 1810
rect 6590 1810 6625 1820
rect 7050 1810 7090 1820
rect 6590 1800 6595 1810
rect 6520 1790 6595 1800
rect 6615 1790 6625 1810
rect 6490 1780 6625 1790
rect 6645 1800 6685 1810
rect 7050 1800 7060 1810
rect 6645 1780 6655 1800
rect 6675 1790 7060 1800
rect 7080 1790 7090 1810
rect 6675 1780 7090 1790
rect 7120 1810 7150 1820
rect 7120 1790 7125 1810
rect 7145 1800 7150 1810
rect 7700 1810 7740 1820
rect 7145 1790 7385 1800
rect 7120 1780 7385 1790
rect 7700 1790 7710 1810
rect 7730 1800 7740 1810
rect 7810 1810 7850 1820
rect 7810 1800 7820 1810
rect 7730 1790 7820 1800
rect 7840 1790 7850 1810
rect 7700 1780 7850 1790
rect 8375 1815 8415 1820
rect 8375 1795 8385 1815
rect 8405 1805 8415 1815
rect 8580 1815 8620 1820
rect 8580 1805 8590 1815
rect 8405 1795 8590 1805
rect 8610 1795 8620 1815
rect 8375 1785 8620 1795
rect 9555 1810 9595 1820
rect 9555 1790 9565 1810
rect 9585 1800 9595 1810
rect 9845 1810 9885 1820
rect 9845 1800 9855 1810
rect 9585 1790 9855 1800
rect 9875 1790 9885 1810
rect 9555 1780 9885 1790
rect 10205 1810 10245 1820
rect 10205 1790 10215 1810
rect 10235 1800 10245 1810
rect 10495 1810 10535 1820
rect 10495 1800 10505 1810
rect 10235 1790 10505 1800
rect 10525 1790 10535 1810
rect 10205 1780 10535 1790
rect 10855 1810 10895 1820
rect 10855 1790 10865 1810
rect 10885 1800 10895 1810
rect 11145 1810 11185 1820
rect 11145 1800 11155 1810
rect 10885 1790 11155 1800
rect 11175 1790 11185 1810
rect 10855 1780 11185 1790
rect 6645 1770 6685 1780
rect 7365 1760 7385 1780
rect 9575 1760 9595 1780
rect 10225 1760 10245 1780
rect 10875 1760 10895 1780
rect 7365 1750 7405 1760
rect 7365 1730 7375 1750
rect 7395 1730 7405 1750
rect 7365 1720 7405 1730
rect 6120 1670 6160 1675
rect 6120 1640 6125 1670
rect 6155 1640 6160 1670
rect 11376 1665 11405 1670
rect 8115 1655 8155 1665
rect 6120 1635 6160 1640
rect 6975 1650 7275 1655
rect 6975 1630 6985 1650
rect 7005 1635 7245 1650
rect 7005 1630 7015 1635
rect 6975 1620 7015 1630
rect 7235 1630 7245 1635
rect 7265 1630 7275 1650
rect 7235 1620 7275 1630
rect 8115 1635 8125 1655
rect 8145 1635 8155 1655
rect 8115 1625 8155 1635
rect 11376 1639 11378 1665
rect 11404 1639 11405 1665
rect 11376 1630 11405 1639
rect 6645 1540 6685 1550
rect 8115 1540 8135 1625
rect 6150 1530 6190 1540
rect 6645 1530 6655 1540
rect 6150 1510 6160 1530
rect 6180 1520 6655 1530
rect 6675 1520 6685 1540
rect 6180 1510 6685 1520
rect 6710 1535 6750 1540
rect 6710 1515 6720 1535
rect 6740 1525 6750 1535
rect 7180 1535 7220 1540
rect 7180 1525 7190 1535
rect 6740 1515 7190 1525
rect 7210 1525 7220 1535
rect 7980 1535 8020 1540
rect 7980 1525 7990 1535
rect 7210 1515 7990 1525
rect 8010 1515 8020 1535
rect 8115 1530 9320 1540
rect 8115 1520 9292 1530
rect 6150 1500 6190 1510
rect 6710 1505 8020 1515
rect 9287 1510 9292 1520
rect 9312 1510 9320 1530
rect 9287 1500 9320 1510
rect 6250 1480 6290 1485
rect 6250 1450 6255 1480
rect 6285 1450 6290 1480
rect 6250 1445 6290 1450
rect 6360 1480 6400 1485
rect 6360 1450 6365 1480
rect 6395 1450 6400 1480
rect 6360 1445 6400 1450
rect 6595 1480 6635 1485
rect 6595 1450 6600 1480
rect 6630 1450 6635 1480
rect 6595 1445 6635 1450
rect 6765 1480 6805 1485
rect 6765 1450 6770 1480
rect 6800 1450 6805 1480
rect 6765 1445 6805 1450
rect 6875 1480 6915 1485
rect 6875 1450 6880 1480
rect 6910 1450 6915 1480
rect 6875 1445 6915 1450
rect 7095 1480 7135 1485
rect 7095 1450 7100 1480
rect 7130 1450 7135 1480
rect 7095 1445 7135 1450
rect 7330 1480 7370 1485
rect 7330 1450 7335 1480
rect 7365 1450 7370 1480
rect 7330 1445 7370 1450
rect 7455 1480 7495 1485
rect 7455 1450 7460 1480
rect 7490 1450 7495 1480
rect 7455 1445 7495 1450
rect 7565 1480 7605 1485
rect 7565 1450 7570 1480
rect 7600 1450 7605 1480
rect 7565 1445 7605 1450
rect 7800 1480 7840 1485
rect 7800 1450 7805 1480
rect 7835 1450 7840 1480
rect 7800 1445 7840 1450
rect 8030 1480 8070 1485
rect 8030 1450 8035 1480
rect 8065 1450 8070 1480
rect 8030 1445 8070 1450
rect 8205 1480 8245 1485
rect 8205 1450 8210 1480
rect 8240 1450 8245 1480
rect 8205 1445 8245 1450
rect 8330 1480 8370 1485
rect 8330 1450 8335 1480
rect 8365 1450 8370 1480
rect 8330 1445 8370 1450
rect 8440 1480 8480 1485
rect 8440 1450 8445 1480
rect 8475 1450 8480 1480
rect 8440 1445 8480 1450
rect 8605 1480 8645 1485
rect 8605 1450 8610 1480
rect 8640 1450 8645 1480
rect 8605 1445 8645 1450
rect 8935 1480 8975 1485
rect 8935 1450 8940 1480
rect 8970 1450 8975 1480
rect 8935 1445 8975 1450
rect 9045 1480 9085 1485
rect 9045 1450 9050 1480
rect 9080 1450 9085 1480
rect 9045 1445 9085 1450
rect 9330 1480 9370 1485
rect 9330 1450 9335 1480
rect 9365 1450 9370 1480
rect 9330 1445 9370 1450
rect 9460 1480 9500 1485
rect 9460 1450 9465 1480
rect 9495 1450 9500 1480
rect 9460 1445 9500 1450
rect 9585 1480 9625 1485
rect 9585 1450 9590 1480
rect 9620 1450 9625 1480
rect 9585 1445 9625 1450
rect 9695 1480 9735 1485
rect 9695 1450 9700 1480
rect 9730 1450 9735 1480
rect 9695 1445 9735 1450
rect 9970 1480 10010 1485
rect 9970 1450 9975 1480
rect 10005 1450 10010 1480
rect 9970 1445 10010 1450
rect 10110 1480 10150 1485
rect 10110 1450 10115 1480
rect 10145 1450 10150 1480
rect 10110 1445 10150 1450
rect 10235 1480 10275 1485
rect 10235 1450 10240 1480
rect 10270 1450 10275 1480
rect 10235 1445 10275 1450
rect 10345 1480 10385 1485
rect 10345 1450 10350 1480
rect 10380 1450 10385 1480
rect 10345 1445 10385 1450
rect 10620 1480 10660 1485
rect 10620 1450 10625 1480
rect 10655 1450 10660 1480
rect 10620 1445 10660 1450
rect 10760 1480 10800 1485
rect 10760 1450 10765 1480
rect 10795 1450 10800 1480
rect 10760 1445 10800 1450
rect 10885 1480 10925 1485
rect 10885 1450 10890 1480
rect 10920 1450 10925 1480
rect 10885 1445 10925 1450
rect 10995 1480 11035 1485
rect 10995 1450 11000 1480
rect 11030 1450 11035 1480
rect 10995 1445 11035 1450
rect 11270 1480 11310 1485
rect 11270 1450 11275 1480
rect 11305 1450 11310 1480
rect 11270 1445 11310 1450
<< via1 >>
rect 6335 1865 6365 1870
rect 6335 1845 6340 1865
rect 6340 1845 6360 1865
rect 6360 1845 6365 1865
rect 6335 1840 6365 1845
rect 6545 1865 6575 1870
rect 6545 1845 6550 1865
rect 6550 1845 6570 1865
rect 6570 1845 6575 1865
rect 6545 1840 6575 1845
rect 6880 1865 6910 1870
rect 6880 1845 6885 1865
rect 6885 1845 6905 1865
rect 6905 1845 6910 1865
rect 6880 1840 6910 1845
rect 7165 1865 7195 1870
rect 7165 1845 7170 1865
rect 7170 1845 7190 1865
rect 7190 1845 7195 1865
rect 7165 1840 7195 1845
rect 7540 1865 7570 1870
rect 7540 1845 7545 1865
rect 7545 1845 7565 1865
rect 7565 1845 7570 1865
rect 7540 1840 7570 1845
rect 7755 1865 7785 1870
rect 7755 1845 7760 1865
rect 7760 1845 7780 1865
rect 7780 1845 7785 1865
rect 7755 1840 7785 1845
rect 7975 1865 8005 1870
rect 7975 1845 7980 1865
rect 7980 1845 8000 1865
rect 8000 1845 8005 1865
rect 7975 1840 8005 1845
rect 8100 1865 8130 1870
rect 8100 1845 8105 1865
rect 8105 1845 8125 1865
rect 8125 1845 8130 1865
rect 8100 1840 8130 1845
rect 8210 1865 8240 1870
rect 8210 1845 8215 1865
rect 8215 1845 8235 1865
rect 8235 1845 8240 1865
rect 8210 1840 8240 1845
rect 8445 1865 8475 1870
rect 8445 1845 8450 1865
rect 8450 1845 8470 1865
rect 8470 1845 8475 1865
rect 8445 1840 8475 1845
rect 8665 1865 8695 1870
rect 8665 1845 8670 1865
rect 8670 1845 8690 1865
rect 8690 1845 8695 1865
rect 8665 1840 8695 1845
rect 8975 1865 9005 1870
rect 8975 1845 8980 1865
rect 8980 1845 9000 1865
rect 9000 1845 9005 1865
rect 8975 1840 9005 1845
rect 9145 1865 9175 1870
rect 9145 1845 9150 1865
rect 9150 1845 9170 1865
rect 9170 1845 9175 1865
rect 9145 1840 9175 1845
rect 9325 1865 9355 1870
rect 9325 1845 9330 1865
rect 9330 1845 9350 1865
rect 9350 1845 9355 1865
rect 9325 1840 9355 1845
rect 9625 1865 9655 1870
rect 9625 1845 9630 1865
rect 9630 1845 9650 1865
rect 9650 1845 9655 1865
rect 9625 1840 9655 1845
rect 9795 1865 9825 1870
rect 9795 1845 9800 1865
rect 9800 1845 9820 1865
rect 9820 1845 9825 1865
rect 9795 1840 9825 1845
rect 9975 1865 10005 1870
rect 9975 1845 9980 1865
rect 9980 1845 10000 1865
rect 10000 1845 10005 1865
rect 9975 1840 10005 1845
rect 10275 1865 10305 1870
rect 10275 1845 10280 1865
rect 10280 1845 10300 1865
rect 10300 1845 10305 1865
rect 10275 1840 10305 1845
rect 10445 1865 10475 1870
rect 10445 1845 10450 1865
rect 10450 1845 10470 1865
rect 10470 1845 10475 1865
rect 10445 1840 10475 1845
rect 10625 1865 10655 1870
rect 10625 1845 10630 1865
rect 10630 1845 10650 1865
rect 10650 1845 10655 1865
rect 10625 1840 10655 1845
rect 10925 1865 10955 1870
rect 10925 1845 10930 1865
rect 10930 1845 10950 1865
rect 10950 1845 10955 1865
rect 10925 1840 10955 1845
rect 11095 1865 11125 1870
rect 11095 1845 11100 1865
rect 11100 1845 11120 1865
rect 11120 1845 11125 1865
rect 11095 1840 11125 1845
rect 11275 1865 11305 1870
rect 11275 1845 11280 1865
rect 11280 1845 11300 1865
rect 11300 1845 11305 1865
rect 11275 1840 11305 1845
rect 6125 1665 6155 1670
rect 6125 1645 6130 1665
rect 6130 1645 6150 1665
rect 6150 1645 6155 1665
rect 6125 1640 6155 1645
rect 11378 1661 11404 1665
rect 11378 1644 11382 1661
rect 11382 1644 11399 1661
rect 11399 1644 11404 1661
rect 11378 1639 11404 1644
rect 6255 1475 6285 1480
rect 6255 1455 6260 1475
rect 6260 1455 6280 1475
rect 6280 1455 6285 1475
rect 6255 1450 6285 1455
rect 6365 1475 6395 1480
rect 6365 1455 6370 1475
rect 6370 1455 6390 1475
rect 6390 1455 6395 1475
rect 6365 1450 6395 1455
rect 6600 1475 6630 1480
rect 6600 1455 6605 1475
rect 6605 1455 6625 1475
rect 6625 1455 6630 1475
rect 6600 1450 6630 1455
rect 6770 1475 6800 1480
rect 6770 1455 6775 1475
rect 6775 1455 6795 1475
rect 6795 1455 6800 1475
rect 6770 1450 6800 1455
rect 6880 1475 6910 1480
rect 6880 1455 6885 1475
rect 6885 1455 6905 1475
rect 6905 1455 6910 1475
rect 6880 1450 6910 1455
rect 7100 1475 7130 1480
rect 7100 1455 7105 1475
rect 7105 1455 7125 1475
rect 7125 1455 7130 1475
rect 7100 1450 7130 1455
rect 7335 1475 7365 1480
rect 7335 1455 7340 1475
rect 7340 1455 7360 1475
rect 7360 1455 7365 1475
rect 7335 1450 7365 1455
rect 7460 1475 7490 1480
rect 7460 1455 7465 1475
rect 7465 1455 7485 1475
rect 7485 1455 7490 1475
rect 7460 1450 7490 1455
rect 7570 1475 7600 1480
rect 7570 1455 7575 1475
rect 7575 1455 7595 1475
rect 7595 1455 7600 1475
rect 7570 1450 7600 1455
rect 7805 1475 7835 1480
rect 7805 1455 7810 1475
rect 7810 1455 7830 1475
rect 7830 1455 7835 1475
rect 7805 1450 7835 1455
rect 8035 1475 8065 1480
rect 8035 1455 8040 1475
rect 8040 1455 8060 1475
rect 8060 1455 8065 1475
rect 8035 1450 8065 1455
rect 8210 1475 8240 1480
rect 8210 1455 8215 1475
rect 8215 1455 8235 1475
rect 8235 1455 8240 1475
rect 8210 1450 8240 1455
rect 8335 1475 8365 1480
rect 8335 1455 8340 1475
rect 8340 1455 8360 1475
rect 8360 1455 8365 1475
rect 8335 1450 8365 1455
rect 8445 1475 8475 1480
rect 8445 1455 8450 1475
rect 8450 1455 8470 1475
rect 8470 1455 8475 1475
rect 8445 1450 8475 1455
rect 8610 1475 8640 1480
rect 8610 1455 8615 1475
rect 8615 1455 8635 1475
rect 8635 1455 8640 1475
rect 8610 1450 8640 1455
rect 8940 1475 8970 1480
rect 8940 1455 8945 1475
rect 8945 1455 8965 1475
rect 8965 1455 8970 1475
rect 8940 1450 8970 1455
rect 9050 1475 9080 1480
rect 9050 1455 9055 1475
rect 9055 1455 9075 1475
rect 9075 1455 9080 1475
rect 9050 1450 9080 1455
rect 9335 1475 9365 1480
rect 9335 1455 9340 1475
rect 9340 1455 9360 1475
rect 9360 1455 9365 1475
rect 9335 1450 9365 1455
rect 9465 1475 9495 1480
rect 9465 1455 9470 1475
rect 9470 1455 9490 1475
rect 9490 1455 9495 1475
rect 9465 1450 9495 1455
rect 9590 1475 9620 1480
rect 9590 1455 9595 1475
rect 9595 1455 9615 1475
rect 9615 1455 9620 1475
rect 9590 1450 9620 1455
rect 9700 1475 9730 1480
rect 9700 1455 9705 1475
rect 9705 1455 9725 1475
rect 9725 1455 9730 1475
rect 9700 1450 9730 1455
rect 9975 1475 10005 1480
rect 9975 1455 9980 1475
rect 9980 1455 10000 1475
rect 10000 1455 10005 1475
rect 9975 1450 10005 1455
rect 10115 1475 10145 1480
rect 10115 1455 10120 1475
rect 10120 1455 10140 1475
rect 10140 1455 10145 1475
rect 10115 1450 10145 1455
rect 10240 1475 10270 1480
rect 10240 1455 10245 1475
rect 10245 1455 10265 1475
rect 10265 1455 10270 1475
rect 10240 1450 10270 1455
rect 10350 1475 10380 1480
rect 10350 1455 10355 1475
rect 10355 1455 10375 1475
rect 10375 1455 10380 1475
rect 10350 1450 10380 1455
rect 10625 1475 10655 1480
rect 10625 1455 10630 1475
rect 10630 1455 10650 1475
rect 10650 1455 10655 1475
rect 10625 1450 10655 1455
rect 10765 1475 10795 1480
rect 10765 1455 10770 1475
rect 10770 1455 10790 1475
rect 10790 1455 10795 1475
rect 10765 1450 10795 1455
rect 10890 1475 10920 1480
rect 10890 1455 10895 1475
rect 10895 1455 10915 1475
rect 10915 1455 10920 1475
rect 10890 1450 10920 1455
rect 11000 1475 11030 1480
rect 11000 1455 11005 1475
rect 11005 1455 11025 1475
rect 11025 1455 11030 1475
rect 11000 1450 11030 1455
rect 11275 1475 11305 1480
rect 11275 1455 11280 1475
rect 11280 1455 11300 1475
rect 11300 1455 11305 1475
rect 11275 1450 11305 1455
<< metal2 >>
rect 6130 1870 11310 1875
rect 6130 1840 6335 1870
rect 6365 1840 6545 1870
rect 6575 1840 6880 1870
rect 6910 1840 7165 1870
rect 7195 1840 7540 1870
rect 7570 1840 7755 1870
rect 7785 1840 7975 1870
rect 8005 1840 8100 1870
rect 8130 1840 8210 1870
rect 8240 1840 8445 1870
rect 8475 1840 8665 1870
rect 8695 1840 8975 1870
rect 9005 1840 9145 1870
rect 9175 1840 9325 1870
rect 9355 1840 9625 1870
rect 9655 1840 9795 1870
rect 9825 1840 9975 1870
rect 10005 1840 10275 1870
rect 10305 1840 10445 1870
rect 10475 1840 10625 1870
rect 10655 1840 10925 1870
rect 10955 1840 11095 1870
rect 11125 1840 11275 1870
rect 11305 1840 11310 1870
rect 6130 1835 11310 1840
rect 6065 1670 6160 1675
rect 6065 1640 6125 1670
rect 6155 1640 6160 1670
rect 6065 1635 6160 1640
rect 11376 1665 11405 1670
rect 11376 1639 11378 1665
rect 11404 1639 11405 1665
rect 11376 1630 11405 1639
rect 6130 1480 11310 1485
rect 6130 1450 6255 1480
rect 6285 1450 6365 1480
rect 6395 1450 6600 1480
rect 6630 1450 6770 1480
rect 6800 1450 6880 1480
rect 6910 1450 7100 1480
rect 7130 1450 7335 1480
rect 7365 1450 7460 1480
rect 7490 1450 7570 1480
rect 7600 1450 7805 1480
rect 7835 1450 8035 1480
rect 8065 1450 8210 1480
rect 8240 1450 8335 1480
rect 8365 1450 8445 1480
rect 8475 1450 8610 1480
rect 8640 1450 8940 1480
rect 8970 1450 9050 1480
rect 9080 1450 9335 1480
rect 9365 1450 9465 1480
rect 9495 1450 9590 1480
rect 9620 1450 9700 1480
rect 9730 1450 9975 1480
rect 10005 1450 10115 1480
rect 10145 1450 10240 1480
rect 10270 1450 10350 1480
rect 10380 1450 10625 1480
rect 10655 1450 10765 1480
rect 10795 1450 10890 1480
rect 10920 1450 11000 1480
rect 11030 1450 11275 1480
rect 11305 1450 11310 1480
rect 6130 1445 11310 1450
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
