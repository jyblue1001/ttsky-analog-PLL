magic
tech sky130A
magscale 1 2
timestamp 1757393692
<< nwell >>
rect 49300 11490 52740 12800
rect 52997 11427 53521 13791
rect 52997 9157 53521 11171
<< nmos >>
rect 49540 10960 49570 11060
rect 49670 10960 49700 11060
rect 49800 10960 49830 11060
rect 49930 10960 49960 11060
rect 50060 10960 50090 11060
rect 50190 10960 50220 11060
rect 50680 10960 50710 11060
rect 50810 10960 50840 11060
rect 50940 10960 50970 11060
rect 51070 10960 51100 11060
rect 51200 10960 51230 11060
rect 51330 10960 51360 11060
rect 51820 10960 51850 11060
rect 51950 10960 51980 11060
rect 52080 10960 52110 11060
rect 52210 10960 52240 11060
rect 52340 10960 52370 11060
rect 52470 10960 52500 11060
rect 49490 10270 49590 10520
rect 49690 10270 49790 10520
rect 49890 10270 49990 10520
rect 50090 10270 50190 10520
rect 50290 10270 50390 10520
rect 50490 10270 50590 10520
rect 50690 10270 50790 10520
rect 50890 10270 50990 10520
rect 51090 10270 51190 10520
rect 51290 10270 51390 10520
<< pmos >>
rect 49610 12190 49710 12690
rect 49810 12190 49910 12690
rect 50010 12190 50110 12690
rect 50210 12190 50310 12690
rect 50410 12190 50510 12690
rect 50610 12190 50710 12690
rect 50810 12190 50910 12690
rect 51010 12190 51110 12690
rect 51210 12190 51310 12690
rect 51410 12190 51510 12690
rect 49540 11540 49570 11740
rect 49670 11540 49700 11740
rect 49800 11540 49830 11740
rect 49930 11540 49960 11740
rect 50060 11540 50090 11740
rect 50190 11540 50220 11740
rect 50680 11540 50710 11740
rect 50810 11540 50840 11740
rect 50940 11540 50970 11740
rect 51070 11540 51100 11740
rect 51200 11540 51230 11740
rect 51330 11540 51360 11740
rect 51820 11540 51850 11740
rect 51950 11540 51980 11740
rect 52080 11540 52110 11740
rect 52210 11540 52240 11740
rect 52340 11540 52370 11740
rect 52470 11540 52500 11740
<< ndiff >>
rect 49440 11030 49540 11060
rect 49440 10990 49470 11030
rect 49510 10990 49540 11030
rect 49440 10960 49540 10990
rect 49570 11030 49670 11060
rect 49570 10990 49600 11030
rect 49640 10990 49670 11030
rect 49570 10960 49670 10990
rect 49700 11030 49800 11060
rect 49700 10990 49730 11030
rect 49770 10990 49800 11030
rect 49700 10960 49800 10990
rect 49830 11030 49930 11060
rect 49830 10990 49860 11030
rect 49900 10990 49930 11030
rect 49830 10960 49930 10990
rect 49960 11030 50060 11060
rect 49960 10990 49990 11030
rect 50030 10990 50060 11030
rect 49960 10960 50060 10990
rect 50090 11030 50190 11060
rect 50090 10990 50120 11030
rect 50160 10990 50190 11030
rect 50090 10960 50190 10990
rect 50220 11030 50320 11060
rect 50220 10990 50250 11030
rect 50290 10990 50320 11030
rect 50220 10960 50320 10990
rect 50580 11030 50680 11060
rect 50580 10990 50610 11030
rect 50650 10990 50680 11030
rect 50580 10960 50680 10990
rect 50710 11030 50810 11060
rect 50710 10990 50740 11030
rect 50780 10990 50810 11030
rect 50710 10960 50810 10990
rect 50840 11030 50940 11060
rect 50840 10990 50870 11030
rect 50910 10990 50940 11030
rect 50840 10960 50940 10990
rect 50970 11030 51070 11060
rect 50970 10990 51000 11030
rect 51040 10990 51070 11030
rect 50970 10960 51070 10990
rect 51100 11030 51200 11060
rect 51100 10990 51130 11030
rect 51170 10990 51200 11030
rect 51100 10960 51200 10990
rect 51230 11030 51330 11060
rect 51230 10990 51260 11030
rect 51300 10990 51330 11030
rect 51230 10960 51330 10990
rect 51360 11030 51460 11060
rect 51360 10990 51390 11030
rect 51430 10990 51460 11030
rect 51360 10960 51460 10990
rect 51720 11030 51820 11060
rect 51720 10990 51750 11030
rect 51790 10990 51820 11030
rect 51720 10960 51820 10990
rect 51850 11030 51950 11060
rect 51850 10990 51880 11030
rect 51920 10990 51950 11030
rect 51850 10960 51950 10990
rect 51980 11030 52080 11060
rect 51980 10990 52010 11030
rect 52050 10990 52080 11030
rect 51980 10960 52080 10990
rect 52110 11030 52210 11060
rect 52110 10990 52140 11030
rect 52180 10990 52210 11030
rect 52110 10960 52210 10990
rect 52240 11030 52340 11060
rect 52240 10990 52270 11030
rect 52310 10990 52340 11030
rect 52240 10960 52340 10990
rect 52370 11030 52470 11060
rect 52370 10990 52400 11030
rect 52440 10990 52470 11030
rect 52370 10960 52470 10990
rect 52500 11030 52600 11060
rect 52500 10990 52530 11030
rect 52570 10990 52600 11030
rect 52500 10960 52600 10990
rect 49390 10490 49490 10520
rect 49390 10440 49420 10490
rect 49460 10440 49490 10490
rect 49390 10350 49490 10440
rect 49390 10300 49420 10350
rect 49460 10300 49490 10350
rect 49390 10270 49490 10300
rect 49590 10490 49690 10520
rect 49590 10440 49620 10490
rect 49660 10440 49690 10490
rect 49590 10350 49690 10440
rect 49590 10300 49620 10350
rect 49660 10300 49690 10350
rect 49590 10270 49690 10300
rect 49790 10490 49890 10520
rect 49790 10440 49820 10490
rect 49860 10440 49890 10490
rect 49790 10350 49890 10440
rect 49790 10300 49820 10350
rect 49860 10300 49890 10350
rect 49790 10270 49890 10300
rect 49990 10490 50090 10520
rect 49990 10440 50020 10490
rect 50060 10440 50090 10490
rect 49990 10350 50090 10440
rect 49990 10300 50020 10350
rect 50060 10300 50090 10350
rect 49990 10270 50090 10300
rect 50190 10490 50290 10520
rect 50190 10440 50220 10490
rect 50260 10440 50290 10490
rect 50190 10350 50290 10440
rect 50190 10300 50220 10350
rect 50260 10300 50290 10350
rect 50190 10270 50290 10300
rect 50390 10490 50490 10520
rect 50390 10440 50420 10490
rect 50460 10440 50490 10490
rect 50390 10350 50490 10440
rect 50390 10300 50420 10350
rect 50460 10300 50490 10350
rect 50390 10270 50490 10300
rect 50590 10490 50690 10520
rect 50590 10440 50620 10490
rect 50660 10440 50690 10490
rect 50590 10350 50690 10440
rect 50590 10300 50620 10350
rect 50660 10300 50690 10350
rect 50590 10270 50690 10300
rect 50790 10490 50890 10520
rect 50790 10440 50820 10490
rect 50860 10440 50890 10490
rect 50790 10350 50890 10440
rect 50790 10300 50820 10350
rect 50860 10300 50890 10350
rect 50790 10270 50890 10300
rect 50990 10490 51090 10520
rect 50990 10440 51020 10490
rect 51060 10440 51090 10490
rect 50990 10350 51090 10440
rect 50990 10300 51020 10350
rect 51060 10300 51090 10350
rect 50990 10270 51090 10300
rect 51190 10490 51290 10520
rect 51190 10440 51220 10490
rect 51260 10440 51290 10490
rect 51190 10350 51290 10440
rect 51190 10300 51220 10350
rect 51260 10300 51290 10350
rect 51190 10270 51290 10300
rect 51390 10490 51490 10520
rect 51390 10440 51420 10490
rect 51460 10440 51490 10490
rect 51390 10350 51490 10440
rect 51390 10300 51420 10350
rect 51460 10300 51490 10350
rect 51390 10270 51490 10300
<< pdiff >>
rect 49510 12660 49610 12690
rect 49510 12620 49540 12660
rect 49580 12620 49610 12660
rect 49510 12560 49610 12620
rect 49510 12520 49540 12560
rect 49580 12520 49610 12560
rect 49510 12460 49610 12520
rect 49510 12420 49540 12460
rect 49580 12420 49610 12460
rect 49510 12360 49610 12420
rect 49510 12320 49540 12360
rect 49580 12320 49610 12360
rect 49510 12260 49610 12320
rect 49510 12220 49540 12260
rect 49580 12220 49610 12260
rect 49510 12190 49610 12220
rect 49710 12660 49810 12690
rect 49710 12620 49740 12660
rect 49780 12620 49810 12660
rect 49710 12560 49810 12620
rect 49710 12520 49740 12560
rect 49780 12520 49810 12560
rect 49710 12460 49810 12520
rect 49710 12420 49740 12460
rect 49780 12420 49810 12460
rect 49710 12360 49810 12420
rect 49710 12320 49740 12360
rect 49780 12320 49810 12360
rect 49710 12260 49810 12320
rect 49710 12220 49740 12260
rect 49780 12220 49810 12260
rect 49710 12190 49810 12220
rect 49910 12660 50010 12690
rect 49910 12620 49940 12660
rect 49980 12620 50010 12660
rect 49910 12560 50010 12620
rect 49910 12520 49940 12560
rect 49980 12520 50010 12560
rect 49910 12460 50010 12520
rect 49910 12420 49940 12460
rect 49980 12420 50010 12460
rect 49910 12360 50010 12420
rect 49910 12320 49940 12360
rect 49980 12320 50010 12360
rect 49910 12260 50010 12320
rect 49910 12220 49940 12260
rect 49980 12220 50010 12260
rect 49910 12190 50010 12220
rect 50110 12660 50210 12690
rect 50110 12620 50140 12660
rect 50180 12620 50210 12660
rect 50110 12560 50210 12620
rect 50110 12520 50140 12560
rect 50180 12520 50210 12560
rect 50110 12460 50210 12520
rect 50110 12420 50140 12460
rect 50180 12420 50210 12460
rect 50110 12360 50210 12420
rect 50110 12320 50140 12360
rect 50180 12320 50210 12360
rect 50110 12260 50210 12320
rect 50110 12220 50140 12260
rect 50180 12220 50210 12260
rect 50110 12190 50210 12220
rect 50310 12660 50410 12690
rect 50310 12620 50340 12660
rect 50380 12620 50410 12660
rect 50310 12560 50410 12620
rect 50310 12520 50340 12560
rect 50380 12520 50410 12560
rect 50310 12460 50410 12520
rect 50310 12420 50340 12460
rect 50380 12420 50410 12460
rect 50310 12360 50410 12420
rect 50310 12320 50340 12360
rect 50380 12320 50410 12360
rect 50310 12260 50410 12320
rect 50310 12220 50340 12260
rect 50380 12220 50410 12260
rect 50310 12190 50410 12220
rect 50510 12660 50610 12690
rect 50510 12620 50540 12660
rect 50580 12620 50610 12660
rect 50510 12560 50610 12620
rect 50510 12520 50540 12560
rect 50580 12520 50610 12560
rect 50510 12460 50610 12520
rect 50510 12420 50540 12460
rect 50580 12420 50610 12460
rect 50510 12360 50610 12420
rect 50510 12320 50540 12360
rect 50580 12320 50610 12360
rect 50510 12260 50610 12320
rect 50510 12220 50540 12260
rect 50580 12220 50610 12260
rect 50510 12190 50610 12220
rect 50710 12660 50810 12690
rect 50710 12620 50740 12660
rect 50780 12620 50810 12660
rect 50710 12560 50810 12620
rect 50710 12520 50740 12560
rect 50780 12520 50810 12560
rect 50710 12460 50810 12520
rect 50710 12420 50740 12460
rect 50780 12420 50810 12460
rect 50710 12360 50810 12420
rect 50710 12320 50740 12360
rect 50780 12320 50810 12360
rect 50710 12260 50810 12320
rect 50710 12220 50740 12260
rect 50780 12220 50810 12260
rect 50710 12190 50810 12220
rect 50910 12660 51010 12690
rect 50910 12620 50940 12660
rect 50980 12620 51010 12660
rect 50910 12560 51010 12620
rect 50910 12520 50940 12560
rect 50980 12520 51010 12560
rect 50910 12460 51010 12520
rect 50910 12420 50940 12460
rect 50980 12420 51010 12460
rect 50910 12360 51010 12420
rect 50910 12320 50940 12360
rect 50980 12320 51010 12360
rect 50910 12260 51010 12320
rect 50910 12220 50940 12260
rect 50980 12220 51010 12260
rect 50910 12190 51010 12220
rect 51110 12660 51210 12690
rect 51110 12620 51140 12660
rect 51180 12620 51210 12660
rect 51110 12560 51210 12620
rect 51110 12520 51140 12560
rect 51180 12520 51210 12560
rect 51110 12460 51210 12520
rect 51110 12420 51140 12460
rect 51180 12420 51210 12460
rect 51110 12360 51210 12420
rect 51110 12320 51140 12360
rect 51180 12320 51210 12360
rect 51110 12260 51210 12320
rect 51110 12220 51140 12260
rect 51180 12220 51210 12260
rect 51110 12190 51210 12220
rect 51310 12660 51410 12690
rect 51310 12620 51340 12660
rect 51380 12620 51410 12660
rect 51310 12560 51410 12620
rect 51310 12520 51340 12560
rect 51380 12520 51410 12560
rect 51310 12460 51410 12520
rect 51310 12420 51340 12460
rect 51380 12420 51410 12460
rect 51310 12360 51410 12420
rect 51310 12320 51340 12360
rect 51380 12320 51410 12360
rect 51310 12260 51410 12320
rect 51310 12220 51340 12260
rect 51380 12220 51410 12260
rect 51310 12190 51410 12220
rect 51510 12660 51610 12690
rect 51510 12620 51540 12660
rect 51580 12620 51610 12660
rect 51510 12560 51610 12620
rect 51510 12520 51540 12560
rect 51580 12520 51610 12560
rect 51510 12460 51610 12520
rect 51510 12420 51540 12460
rect 51580 12420 51610 12460
rect 51510 12360 51610 12420
rect 51510 12320 51540 12360
rect 51580 12320 51610 12360
rect 51510 12260 51610 12320
rect 51510 12220 51540 12260
rect 51580 12220 51610 12260
rect 51510 12190 51610 12220
rect 49440 11710 49540 11740
rect 49440 11670 49470 11710
rect 49510 11670 49540 11710
rect 49440 11610 49540 11670
rect 49440 11570 49470 11610
rect 49510 11570 49540 11610
rect 49440 11540 49540 11570
rect 49570 11710 49670 11740
rect 49570 11670 49600 11710
rect 49640 11670 49670 11710
rect 49570 11610 49670 11670
rect 49570 11570 49600 11610
rect 49640 11570 49670 11610
rect 49570 11540 49670 11570
rect 49700 11710 49800 11740
rect 49700 11670 49730 11710
rect 49770 11670 49800 11710
rect 49700 11610 49800 11670
rect 49700 11570 49730 11610
rect 49770 11570 49800 11610
rect 49700 11540 49800 11570
rect 49830 11710 49930 11740
rect 49830 11670 49860 11710
rect 49900 11670 49930 11710
rect 49830 11610 49930 11670
rect 49830 11570 49860 11610
rect 49900 11570 49930 11610
rect 49830 11540 49930 11570
rect 49960 11710 50060 11740
rect 49960 11670 49990 11710
rect 50030 11670 50060 11710
rect 49960 11610 50060 11670
rect 49960 11570 49990 11610
rect 50030 11570 50060 11610
rect 49960 11540 50060 11570
rect 50090 11710 50190 11740
rect 50090 11670 50120 11710
rect 50160 11670 50190 11710
rect 50090 11610 50190 11670
rect 50090 11570 50120 11610
rect 50160 11570 50190 11610
rect 50090 11540 50190 11570
rect 50220 11710 50320 11740
rect 50220 11670 50250 11710
rect 50290 11670 50320 11710
rect 50220 11610 50320 11670
rect 50220 11570 50250 11610
rect 50290 11570 50320 11610
rect 50220 11540 50320 11570
rect 50580 11710 50680 11740
rect 50580 11670 50610 11710
rect 50650 11670 50680 11710
rect 50580 11610 50680 11670
rect 50580 11570 50610 11610
rect 50650 11570 50680 11610
rect 50580 11540 50680 11570
rect 50710 11710 50810 11740
rect 50710 11670 50740 11710
rect 50780 11670 50810 11710
rect 50710 11610 50810 11670
rect 50710 11570 50740 11610
rect 50780 11570 50810 11610
rect 50710 11540 50810 11570
rect 50840 11710 50940 11740
rect 50840 11670 50870 11710
rect 50910 11670 50940 11710
rect 50840 11610 50940 11670
rect 50840 11570 50870 11610
rect 50910 11570 50940 11610
rect 50840 11540 50940 11570
rect 50970 11710 51070 11740
rect 50970 11670 51000 11710
rect 51040 11670 51070 11710
rect 50970 11610 51070 11670
rect 50970 11570 51000 11610
rect 51040 11570 51070 11610
rect 50970 11540 51070 11570
rect 51100 11710 51200 11740
rect 51100 11670 51130 11710
rect 51170 11670 51200 11710
rect 51100 11610 51200 11670
rect 51100 11570 51130 11610
rect 51170 11570 51200 11610
rect 51100 11540 51200 11570
rect 51230 11710 51330 11740
rect 51230 11670 51260 11710
rect 51300 11670 51330 11710
rect 51230 11610 51330 11670
rect 51230 11570 51260 11610
rect 51300 11570 51330 11610
rect 51230 11540 51330 11570
rect 51360 11710 51460 11740
rect 51360 11670 51390 11710
rect 51430 11670 51460 11710
rect 51360 11610 51460 11670
rect 51360 11570 51390 11610
rect 51430 11570 51460 11610
rect 51360 11540 51460 11570
rect 51720 11710 51820 11740
rect 51720 11670 51750 11710
rect 51790 11670 51820 11710
rect 51720 11610 51820 11670
rect 51720 11570 51750 11610
rect 51790 11570 51820 11610
rect 51720 11540 51820 11570
rect 51850 11710 51950 11740
rect 51850 11670 51880 11710
rect 51920 11670 51950 11710
rect 51850 11610 51950 11670
rect 51850 11570 51880 11610
rect 51920 11570 51950 11610
rect 51850 11540 51950 11570
rect 51980 11710 52080 11740
rect 51980 11670 52010 11710
rect 52050 11670 52080 11710
rect 51980 11610 52080 11670
rect 51980 11570 52010 11610
rect 52050 11570 52080 11610
rect 51980 11540 52080 11570
rect 52110 11710 52210 11740
rect 52110 11670 52140 11710
rect 52180 11670 52210 11710
rect 52110 11610 52210 11670
rect 52110 11570 52140 11610
rect 52180 11570 52210 11610
rect 52110 11540 52210 11570
rect 52240 11710 52340 11740
rect 52240 11670 52270 11710
rect 52310 11670 52340 11710
rect 52240 11610 52340 11670
rect 52240 11570 52270 11610
rect 52310 11570 52340 11610
rect 52240 11540 52340 11570
rect 52370 11710 52470 11740
rect 52370 11670 52400 11710
rect 52440 11670 52470 11710
rect 52370 11610 52470 11670
rect 52370 11570 52400 11610
rect 52440 11570 52470 11610
rect 52370 11540 52470 11570
rect 52500 11710 52600 11740
rect 52500 11670 52530 11710
rect 52570 11670 52600 11710
rect 52500 11610 52600 11670
rect 52500 11570 52530 11610
rect 52570 11570 52600 11610
rect 52500 11540 52600 11570
<< ndiffc >>
rect 49470 10990 49510 11030
rect 49600 10990 49640 11030
rect 49730 10990 49770 11030
rect 49860 10990 49900 11030
rect 49990 10990 50030 11030
rect 50120 10990 50160 11030
rect 50250 10990 50290 11030
rect 50610 10990 50650 11030
rect 50740 10990 50780 11030
rect 50870 10990 50910 11030
rect 51000 10990 51040 11030
rect 51130 10990 51170 11030
rect 51260 10990 51300 11030
rect 51390 10990 51430 11030
rect 51750 10990 51790 11030
rect 51880 10990 51920 11030
rect 52010 10990 52050 11030
rect 52140 10990 52180 11030
rect 52270 10990 52310 11030
rect 52400 10990 52440 11030
rect 52530 10990 52570 11030
rect 49420 10440 49460 10490
rect 49420 10300 49460 10350
rect 49620 10440 49660 10490
rect 49620 10300 49660 10350
rect 49820 10440 49860 10490
rect 49820 10300 49860 10350
rect 50020 10440 50060 10490
rect 50020 10300 50060 10350
rect 50220 10440 50260 10490
rect 50220 10300 50260 10350
rect 50420 10440 50460 10490
rect 50420 10300 50460 10350
rect 50620 10440 50660 10490
rect 50620 10300 50660 10350
rect 50820 10440 50860 10490
rect 50820 10300 50860 10350
rect 51020 10440 51060 10490
rect 51020 10300 51060 10350
rect 51220 10440 51260 10490
rect 51220 10300 51260 10350
rect 51420 10440 51460 10490
rect 51420 10300 51460 10350
<< pdiffc >>
rect 49540 12620 49580 12660
rect 49540 12520 49580 12560
rect 49540 12420 49580 12460
rect 49540 12320 49580 12360
rect 49540 12220 49580 12260
rect 49740 12620 49780 12660
rect 49740 12520 49780 12560
rect 49740 12420 49780 12460
rect 49740 12320 49780 12360
rect 49740 12220 49780 12260
rect 49940 12620 49980 12660
rect 49940 12520 49980 12560
rect 49940 12420 49980 12460
rect 49940 12320 49980 12360
rect 49940 12220 49980 12260
rect 50140 12620 50180 12660
rect 50140 12520 50180 12560
rect 50140 12420 50180 12460
rect 50140 12320 50180 12360
rect 50140 12220 50180 12260
rect 50340 12620 50380 12660
rect 50340 12520 50380 12560
rect 50340 12420 50380 12460
rect 50340 12320 50380 12360
rect 50340 12220 50380 12260
rect 50540 12620 50580 12660
rect 50540 12520 50580 12560
rect 50540 12420 50580 12460
rect 50540 12320 50580 12360
rect 50540 12220 50580 12260
rect 50740 12620 50780 12660
rect 50740 12520 50780 12560
rect 50740 12420 50780 12460
rect 50740 12320 50780 12360
rect 50740 12220 50780 12260
rect 50940 12620 50980 12660
rect 50940 12520 50980 12560
rect 50940 12420 50980 12460
rect 50940 12320 50980 12360
rect 50940 12220 50980 12260
rect 51140 12620 51180 12660
rect 51140 12520 51180 12560
rect 51140 12420 51180 12460
rect 51140 12320 51180 12360
rect 51140 12220 51180 12260
rect 51340 12620 51380 12660
rect 51340 12520 51380 12560
rect 51340 12420 51380 12460
rect 51340 12320 51380 12360
rect 51340 12220 51380 12260
rect 51540 12620 51580 12660
rect 51540 12520 51580 12560
rect 51540 12420 51580 12460
rect 51540 12320 51580 12360
rect 51540 12220 51580 12260
rect 49470 11670 49510 11710
rect 49470 11570 49510 11610
rect 49600 11670 49640 11710
rect 49600 11570 49640 11610
rect 49730 11670 49770 11710
rect 49730 11570 49770 11610
rect 49860 11670 49900 11710
rect 49860 11570 49900 11610
rect 49990 11670 50030 11710
rect 49990 11570 50030 11610
rect 50120 11670 50160 11710
rect 50120 11570 50160 11610
rect 50250 11670 50290 11710
rect 50250 11570 50290 11610
rect 50610 11670 50650 11710
rect 50610 11570 50650 11610
rect 50740 11670 50780 11710
rect 50740 11570 50780 11610
rect 50870 11670 50910 11710
rect 50870 11570 50910 11610
rect 51000 11670 51040 11710
rect 51000 11570 51040 11610
rect 51130 11670 51170 11710
rect 51130 11570 51170 11610
rect 51260 11670 51300 11710
rect 51260 11570 51300 11610
rect 51390 11670 51430 11710
rect 51390 11570 51430 11610
rect 51750 11670 51790 11710
rect 51750 11570 51790 11610
rect 51880 11670 51920 11710
rect 51880 11570 51920 11610
rect 52010 11670 52050 11710
rect 52010 11570 52050 11610
rect 52140 11670 52180 11710
rect 52140 11570 52180 11610
rect 52270 11670 52310 11710
rect 52270 11570 52310 11610
rect 52400 11670 52440 11710
rect 52400 11570 52440 11610
rect 52530 11670 52570 11710
rect 52530 11570 52570 11610
<< psubdiff >>
rect 49340 11030 49440 11060
rect 49340 10990 49370 11030
rect 49410 10990 49440 11030
rect 49340 10960 49440 10990
rect 50320 11030 50420 11060
rect 50320 10990 50350 11030
rect 50390 10990 50420 11030
rect 50320 10960 50420 10990
rect 51620 11030 51720 11060
rect 51620 10990 51650 11030
rect 51690 10990 51720 11030
rect 51620 10960 51720 10990
rect 52600 11030 52700 11060
rect 52600 10990 52630 11030
rect 52670 10990 52700 11030
rect 52600 10960 52700 10990
rect 49290 10490 49390 10520
rect 49290 10440 49320 10490
rect 49360 10440 49390 10490
rect 49290 10350 49390 10440
rect 49290 10300 49320 10350
rect 49360 10300 49390 10350
rect 49290 10270 49390 10300
rect 51490 10490 51590 10520
rect 51490 10440 51520 10490
rect 51560 10440 51590 10490
rect 51490 10350 51590 10440
rect 51490 10300 51520 10350
rect 51560 10300 51590 10350
rect 51490 10270 51590 10300
<< nsubdiff >>
rect 53033 13721 53129 13755
rect 53389 13721 53485 13755
rect 53033 13659 53067 13721
rect 49410 12660 49510 12690
rect 49410 12620 49440 12660
rect 49480 12620 49510 12660
rect 49410 12560 49510 12620
rect 49410 12520 49440 12560
rect 49480 12520 49510 12560
rect 49410 12460 49510 12520
rect 49410 12420 49440 12460
rect 49480 12420 49510 12460
rect 49410 12360 49510 12420
rect 49410 12320 49440 12360
rect 49480 12320 49510 12360
rect 49410 12260 49510 12320
rect 49410 12220 49440 12260
rect 49480 12220 49510 12260
rect 49410 12190 49510 12220
rect 51610 12660 51710 12690
rect 51610 12620 51640 12660
rect 51680 12620 51710 12660
rect 51610 12560 51710 12620
rect 51610 12520 51640 12560
rect 51680 12520 51710 12560
rect 51610 12460 51710 12520
rect 51610 12420 51640 12460
rect 51680 12420 51710 12460
rect 51610 12360 51710 12420
rect 51610 12320 51640 12360
rect 51680 12320 51710 12360
rect 51610 12260 51710 12320
rect 51610 12220 51640 12260
rect 51680 12220 51710 12260
rect 51610 12190 51710 12220
rect 50480 11710 50580 11740
rect 50480 11670 50510 11710
rect 50550 11670 50580 11710
rect 50480 11610 50580 11670
rect 50480 11570 50510 11610
rect 50550 11570 50580 11610
rect 50480 11540 50580 11570
rect 51460 11710 51560 11740
rect 51460 11670 51490 11710
rect 51530 11670 51560 11710
rect 51460 11610 51560 11670
rect 51460 11570 51490 11610
rect 51530 11570 51560 11610
rect 51460 11540 51560 11570
rect 51620 11710 51720 11740
rect 51620 11670 51650 11710
rect 51690 11670 51720 11710
rect 51620 11610 51720 11670
rect 51620 11570 51650 11610
rect 51690 11570 51720 11610
rect 51620 11540 51720 11570
rect 52600 11710 52700 11740
rect 52600 11670 52630 11710
rect 52670 11670 52700 11710
rect 52600 11610 52700 11670
rect 52600 11570 52630 11610
rect 52670 11570 52700 11610
rect 52600 11540 52700 11570
rect 53451 13659 53485 13721
rect 53033 11497 53067 11559
rect 53451 11497 53485 11559
rect 53033 11463 53129 11497
rect 53389 11463 53485 11497
rect 53033 11101 53129 11135
rect 53389 11101 53485 11135
rect 53033 11039 53067 11101
rect 53451 11039 53485 11101
rect 53033 9227 53067 9289
rect 53451 9227 53485 9289
rect 53033 9193 53129 9227
rect 53389 9193 53485 9227
<< psubdiffcont >>
rect 49370 10990 49410 11030
rect 50350 10990 50390 11030
rect 51650 10990 51690 11030
rect 52630 10990 52670 11030
rect 49320 10440 49360 10490
rect 49320 10300 49360 10350
rect 51520 10440 51560 10490
rect 51520 10300 51560 10350
<< nsubdiffcont >>
rect 53129 13721 53389 13755
rect 49440 12620 49480 12660
rect 49440 12520 49480 12560
rect 49440 12420 49480 12460
rect 49440 12320 49480 12360
rect 49440 12220 49480 12260
rect 51640 12620 51680 12660
rect 51640 12520 51680 12560
rect 51640 12420 51680 12460
rect 51640 12320 51680 12360
rect 51640 12220 51680 12260
rect 50510 11670 50550 11710
rect 50510 11570 50550 11610
rect 51490 11670 51530 11710
rect 51490 11570 51530 11610
rect 51650 11670 51690 11710
rect 51650 11570 51690 11610
rect 52630 11670 52670 11710
rect 52630 11570 52670 11610
rect 53033 11559 53067 13659
rect 53451 11559 53485 13659
rect 53129 11463 53389 11497
rect 53129 11101 53389 11135
rect 53033 9289 53067 11039
rect 53451 9289 53485 11039
rect 53129 9193 53389 9227
<< poly >>
rect 50320 12780 50400 12800
rect 50320 12740 50340 12780
rect 50380 12740 50400 12780
rect 50720 12780 50800 12800
rect 50720 12740 50740 12780
rect 50780 12740 50800 12780
rect 49610 12690 49710 12720
rect 49810 12710 51310 12740
rect 49810 12690 49910 12710
rect 50010 12690 50110 12710
rect 50210 12690 50310 12710
rect 50410 12690 50510 12710
rect 50610 12690 50710 12710
rect 50810 12690 50910 12710
rect 51010 12690 51110 12710
rect 51210 12690 51310 12710
rect 51410 12690 51510 12720
rect 49610 12160 49710 12190
rect 49810 12160 49910 12190
rect 50010 12160 50110 12190
rect 50210 12160 50310 12190
rect 50410 12160 50510 12190
rect 50610 12160 50710 12190
rect 50810 12160 50910 12190
rect 51010 12160 51110 12190
rect 51210 12160 51310 12190
rect 51410 12160 51510 12190
rect 49520 12140 49710 12160
rect 49520 12100 49540 12140
rect 49580 12130 49710 12140
rect 51410 12140 51600 12160
rect 51410 12130 51540 12140
rect 49580 12100 49600 12130
rect 49520 12080 49600 12100
rect 51520 12100 51540 12130
rect 51580 12100 51600 12140
rect 51520 12080 51600 12100
rect 49510 11830 49590 11850
rect 49510 11790 49530 11830
rect 49570 11790 49590 11830
rect 49510 11770 49590 11790
rect 50170 11830 50250 11850
rect 50170 11790 50190 11830
rect 50230 11790 50250 11830
rect 50170 11770 50250 11790
rect 50650 11830 50730 11850
rect 50650 11790 50670 11830
rect 50710 11790 50730 11830
rect 50650 11770 50730 11790
rect 51310 11830 51390 11850
rect 51310 11790 51330 11830
rect 51370 11790 51390 11830
rect 51310 11770 51390 11790
rect 51790 11830 51870 11850
rect 51790 11790 51810 11830
rect 51850 11790 51870 11830
rect 51790 11770 51870 11790
rect 52450 11830 52530 11850
rect 52450 11790 52470 11830
rect 52510 11790 52530 11830
rect 52450 11770 52530 11790
rect 49540 11740 49570 11770
rect 49670 11740 49700 11770
rect 49800 11740 49830 11770
rect 49930 11740 49960 11770
rect 50060 11740 50090 11770
rect 50190 11740 50220 11770
rect 50680 11740 50710 11770
rect 50810 11740 50840 11770
rect 50940 11740 50970 11770
rect 51070 11740 51100 11770
rect 51200 11740 51230 11770
rect 51330 11740 51360 11770
rect 51820 11740 51850 11770
rect 51950 11740 51980 11770
rect 52080 11740 52110 11770
rect 52210 11740 52240 11770
rect 52340 11740 52370 11770
rect 52470 11740 52500 11770
rect 49540 11510 49570 11540
rect 49670 11520 49700 11540
rect 49800 11520 49830 11540
rect 49670 11510 49830 11520
rect 49620 11490 49830 11510
rect 49930 11520 49960 11540
rect 50060 11520 50090 11540
rect 49930 11510 50090 11520
rect 50190 11510 50220 11540
rect 50680 11510 50710 11540
rect 50810 11520 50840 11540
rect 50940 11520 50970 11540
rect 51070 11520 51100 11540
rect 51200 11520 51230 11540
rect 49930 11490 50140 11510
rect 50810 11490 51230 11520
rect 51330 11510 51360 11540
rect 51820 11510 51850 11540
rect 51950 11510 51980 11540
rect 51900 11490 51980 11510
rect 49620 11450 49640 11490
rect 49680 11450 49700 11490
rect 49620 11430 49700 11450
rect 50060 11450 50080 11490
rect 50120 11450 50140 11490
rect 50060 11430 50140 11450
rect 50850 11480 50930 11490
rect 50850 11440 50870 11480
rect 50910 11440 50930 11480
rect 50850 11420 50930 11440
rect 51900 11450 51920 11490
rect 51960 11460 51980 11490
rect 52080 11460 52110 11540
rect 52210 11460 52240 11540
rect 52340 11460 52370 11540
rect 52470 11510 52500 11540
rect 52740 11490 52820 11510
rect 52740 11460 52760 11490
rect 51960 11450 52760 11460
rect 52800 11450 52820 11490
rect 51900 11430 52820 11450
rect 51900 11270 51980 11290
rect 51900 11230 51920 11270
rect 51960 11230 51980 11270
rect 51900 11210 51980 11230
rect 51950 11170 51980 11210
rect 49710 11150 49790 11170
rect 49710 11110 49730 11150
rect 49770 11110 49790 11150
rect 50760 11150 50840 11170
rect 50760 11110 50780 11150
rect 50820 11110 50840 11150
rect 51200 11150 51280 11170
rect 51200 11110 51220 11150
rect 51260 11110 51280 11150
rect 49540 11060 49570 11090
rect 49670 11080 50090 11110
rect 50760 11090 50970 11110
rect 49670 11060 49700 11080
rect 49800 11060 49830 11080
rect 49930 11060 49960 11080
rect 50060 11060 50090 11080
rect 50190 11060 50220 11090
rect 50680 11060 50710 11090
rect 50810 11080 50970 11090
rect 50810 11060 50840 11080
rect 50940 11060 50970 11080
rect 51070 11090 51280 11110
rect 51950 11150 52820 11170
rect 51950 11140 52760 11150
rect 51070 11080 51230 11090
rect 51070 11060 51100 11080
rect 51200 11060 51230 11080
rect 51330 11060 51360 11090
rect 51820 11060 51850 11090
rect 51950 11060 51980 11140
rect 52080 11060 52110 11140
rect 52210 11060 52240 11140
rect 52340 11060 52370 11140
rect 52740 11110 52760 11140
rect 52800 11110 52820 11150
rect 52740 11090 52820 11110
rect 52470 11060 52500 11090
rect 49540 10930 49570 10960
rect 49670 10930 49700 10960
rect 49800 10930 49830 10960
rect 49930 10930 49960 10960
rect 50060 10930 50090 10960
rect 50190 10930 50220 10960
rect 50680 10930 50710 10960
rect 50810 10930 50840 10960
rect 50940 10930 50970 10960
rect 51070 10930 51100 10960
rect 51200 10930 51230 10960
rect 51330 10930 51360 10960
rect 51820 10930 51850 10960
rect 51950 10930 51980 10960
rect 52080 10930 52110 10960
rect 52210 10930 52240 10960
rect 52340 10930 52370 10960
rect 52470 10930 52500 10960
rect 49510 10910 49600 10930
rect 49510 10860 49530 10910
rect 49580 10860 49600 10910
rect 49510 10840 49600 10860
rect 50160 10910 50250 10930
rect 50160 10860 50180 10910
rect 50230 10860 50250 10910
rect 50160 10840 50250 10860
rect 50650 10910 50730 10930
rect 50650 10870 50670 10910
rect 50710 10870 50730 10910
rect 50650 10850 50730 10870
rect 51310 10910 51390 10930
rect 51310 10870 51330 10910
rect 51370 10870 51390 10910
rect 51310 10850 51390 10870
rect 51790 10910 51870 10930
rect 51790 10870 51810 10910
rect 51850 10870 51870 10910
rect 51790 10850 51870 10870
rect 52450 10910 52530 10930
rect 52450 10870 52470 10910
rect 52510 10870 52530 10910
rect 52450 10850 52530 10870
rect 49400 10610 49480 10630
rect 49400 10570 49420 10610
rect 49460 10580 49480 10610
rect 51400 10610 51480 10630
rect 51400 10580 51420 10610
rect 49460 10570 49590 10580
rect 49400 10550 49590 10570
rect 51290 10570 51420 10580
rect 51460 10570 51480 10610
rect 51290 10550 51480 10570
rect 49490 10520 49590 10550
rect 49690 10520 49790 10550
rect 49890 10520 49990 10550
rect 50090 10520 50190 10550
rect 50290 10520 50390 10550
rect 50490 10520 50590 10550
rect 50690 10520 50790 10550
rect 50890 10520 50990 10550
rect 51090 10520 51190 10550
rect 51290 10520 51390 10550
rect 49490 10240 49590 10270
rect 49690 10250 49790 10270
rect 49890 10250 49990 10270
rect 50090 10250 50190 10270
rect 50290 10250 50390 10270
rect 50490 10250 50590 10270
rect 50690 10250 50790 10270
rect 50890 10250 50990 10270
rect 51090 10250 51190 10270
rect 49690 10220 51190 10250
rect 51290 10240 51390 10270
rect 50200 10180 50220 10220
rect 50260 10180 50280 10220
rect 50200 10160 50280 10180
rect 50600 10180 50620 10220
rect 50660 10180 50680 10220
rect 50600 10160 50680 10180
rect 49244 10024 49674 10040
rect 49244 9990 49260 10024
rect 49294 9990 49674 10024
rect 49244 9974 49674 9990
rect 50154 10024 50584 10040
rect 50154 9990 50534 10024
rect 50568 9990 50584 10024
rect 50154 9974 50584 9990
<< polycont >>
rect 50340 12740 50380 12780
rect 50740 12740 50780 12780
rect 49540 12100 49580 12140
rect 51540 12100 51580 12140
rect 49530 11790 49570 11830
rect 50190 11790 50230 11830
rect 50670 11790 50710 11830
rect 51330 11790 51370 11830
rect 51810 11790 51850 11830
rect 52470 11790 52510 11830
rect 49640 11450 49680 11490
rect 50080 11450 50120 11490
rect 50870 11440 50910 11480
rect 51920 11450 51960 11490
rect 52760 11450 52800 11490
rect 51920 11230 51960 11270
rect 49730 11110 49770 11150
rect 50780 11110 50820 11150
rect 51220 11110 51260 11150
rect 52760 11110 52800 11150
rect 49530 10860 49580 10910
rect 50180 10860 50230 10910
rect 50670 10870 50710 10910
rect 51330 10870 51370 10910
rect 51810 10870 51850 10910
rect 52470 10870 52510 10910
rect 49420 10570 49460 10610
rect 51420 10570 51460 10610
rect 50220 10180 50260 10220
rect 50620 10180 50660 10220
rect 49260 9990 49294 10024
rect 50534 9990 50568 10024
<< xpolycontact >>
rect 53224 13184 53294 13616
rect 53224 11602 53294 12034
rect 53224 10564 53294 10996
rect 53224 9332 53294 9764
<< npolyres >>
rect 49674 9974 50154 10040
<< ppolyres >>
rect 53224 12034 53294 13184
rect 53224 9764 53294 10564
<< locali >>
rect 53033 13721 53129 13755
rect 53389 13721 53485 13755
rect 53033 13659 53067 13721
rect 53010 13170 53033 13190
rect 53451 13659 53485 13721
rect 53067 13170 53090 13190
rect 53010 13130 53030 13170
rect 53070 13130 53090 13170
rect 53010 13110 53033 13130
rect 50320 12780 50400 12800
rect 50320 12740 50340 12780
rect 50380 12740 50400 12780
rect 50320 12720 50400 12740
rect 50720 12780 50800 12800
rect 50720 12740 50740 12780
rect 50780 12740 50800 12780
rect 50720 12720 50800 12740
rect 49420 12660 49600 12680
rect 49420 12620 49440 12660
rect 49480 12620 49540 12660
rect 49580 12620 49600 12660
rect 49420 12560 49600 12620
rect 49420 12520 49440 12560
rect 49480 12520 49540 12560
rect 49580 12520 49600 12560
rect 49420 12460 49600 12520
rect 49420 12420 49440 12460
rect 49480 12420 49540 12460
rect 49580 12420 49600 12460
rect 49420 12360 49600 12420
rect 49420 12320 49440 12360
rect 49480 12320 49540 12360
rect 49580 12320 49600 12360
rect 49420 12260 49600 12320
rect 49420 12220 49440 12260
rect 49480 12220 49540 12260
rect 49580 12220 49600 12260
rect 49420 12200 49600 12220
rect 49720 12660 49800 12680
rect 49720 12620 49740 12660
rect 49780 12620 49800 12660
rect 49720 12560 49800 12620
rect 49720 12520 49740 12560
rect 49780 12520 49800 12560
rect 49720 12460 49800 12520
rect 49720 12420 49740 12460
rect 49780 12420 49800 12460
rect 49720 12360 49800 12420
rect 49720 12320 49740 12360
rect 49780 12320 49800 12360
rect 49720 12260 49800 12320
rect 49720 12220 49740 12260
rect 49780 12220 49800 12260
rect 49720 12200 49800 12220
rect 49920 12660 50000 12680
rect 49920 12620 49940 12660
rect 49980 12620 50000 12660
rect 49920 12560 50000 12620
rect 49920 12520 49940 12560
rect 49980 12520 50000 12560
rect 49920 12460 50000 12520
rect 49920 12420 49940 12460
rect 49980 12420 50000 12460
rect 49920 12360 50000 12420
rect 49920 12320 49940 12360
rect 49980 12320 50000 12360
rect 49920 12260 50000 12320
rect 49920 12220 49940 12260
rect 49980 12220 50000 12260
rect 49920 12200 50000 12220
rect 50120 12660 50200 12680
rect 50120 12620 50140 12660
rect 50180 12620 50200 12660
rect 50120 12560 50200 12620
rect 50120 12520 50140 12560
rect 50180 12520 50200 12560
rect 50120 12460 50200 12520
rect 50120 12420 50140 12460
rect 50180 12420 50200 12460
rect 50120 12360 50200 12420
rect 50120 12320 50140 12360
rect 50180 12320 50200 12360
rect 50120 12260 50200 12320
rect 50120 12220 50140 12260
rect 50180 12220 50200 12260
rect 50120 12200 50200 12220
rect 50320 12660 50400 12680
rect 50320 12620 50340 12660
rect 50380 12620 50400 12660
rect 50320 12560 50400 12620
rect 50320 12520 50340 12560
rect 50380 12520 50400 12560
rect 50320 12460 50400 12520
rect 50320 12420 50340 12460
rect 50380 12420 50400 12460
rect 50320 12360 50400 12420
rect 50320 12320 50340 12360
rect 50380 12320 50400 12360
rect 50320 12260 50400 12320
rect 50320 12220 50340 12260
rect 50380 12220 50400 12260
rect 50320 12200 50400 12220
rect 50520 12660 50600 12680
rect 50520 12620 50540 12660
rect 50580 12620 50600 12660
rect 50520 12560 50600 12620
rect 50520 12520 50540 12560
rect 50580 12520 50600 12560
rect 50520 12460 50600 12520
rect 50520 12420 50540 12460
rect 50580 12420 50600 12460
rect 50520 12360 50600 12420
rect 50520 12320 50540 12360
rect 50580 12320 50600 12360
rect 50520 12260 50600 12320
rect 50520 12220 50540 12260
rect 50580 12220 50600 12260
rect 50520 12200 50600 12220
rect 50720 12660 50800 12680
rect 50720 12620 50740 12660
rect 50780 12620 50800 12660
rect 50720 12560 50800 12620
rect 50720 12520 50740 12560
rect 50780 12520 50800 12560
rect 50720 12460 50800 12520
rect 50720 12420 50740 12460
rect 50780 12420 50800 12460
rect 50720 12360 50800 12420
rect 50720 12320 50740 12360
rect 50780 12320 50800 12360
rect 50720 12260 50800 12320
rect 50720 12220 50740 12260
rect 50780 12220 50800 12260
rect 50720 12200 50800 12220
rect 50920 12660 51000 12680
rect 50920 12620 50940 12660
rect 50980 12620 51000 12660
rect 50920 12560 51000 12620
rect 50920 12520 50940 12560
rect 50980 12520 51000 12560
rect 50920 12460 51000 12520
rect 50920 12420 50940 12460
rect 50980 12420 51000 12460
rect 50920 12360 51000 12420
rect 50920 12320 50940 12360
rect 50980 12320 51000 12360
rect 50920 12260 51000 12320
rect 50920 12220 50940 12260
rect 50980 12220 51000 12260
rect 50920 12200 51000 12220
rect 51120 12660 51200 12680
rect 51120 12620 51140 12660
rect 51180 12620 51200 12660
rect 51120 12560 51200 12620
rect 51120 12520 51140 12560
rect 51180 12520 51200 12560
rect 51120 12460 51200 12520
rect 51120 12420 51140 12460
rect 51180 12420 51200 12460
rect 51120 12360 51200 12420
rect 51120 12320 51140 12360
rect 51180 12320 51200 12360
rect 51120 12260 51200 12320
rect 51120 12220 51140 12260
rect 51180 12220 51200 12260
rect 51120 12200 51200 12220
rect 51320 12660 51400 12680
rect 51320 12620 51340 12660
rect 51380 12620 51400 12660
rect 51320 12560 51400 12620
rect 51320 12520 51340 12560
rect 51380 12520 51400 12560
rect 51320 12460 51400 12520
rect 51320 12420 51340 12460
rect 51380 12420 51400 12460
rect 51320 12360 51400 12420
rect 51320 12320 51340 12360
rect 51380 12320 51400 12360
rect 51320 12260 51400 12320
rect 51320 12220 51340 12260
rect 51380 12220 51400 12260
rect 51320 12200 51400 12220
rect 51520 12660 51700 12680
rect 51520 12620 51540 12660
rect 51580 12620 51640 12660
rect 51680 12620 51700 12660
rect 51520 12560 51700 12620
rect 51520 12520 51540 12560
rect 51580 12520 51640 12560
rect 51680 12520 51700 12560
rect 51520 12460 51700 12520
rect 51520 12420 51540 12460
rect 51580 12420 51640 12460
rect 51680 12420 51700 12460
rect 51520 12360 51700 12420
rect 51520 12320 51540 12360
rect 51580 12320 51640 12360
rect 51680 12320 51700 12360
rect 51520 12260 51700 12320
rect 51520 12220 51540 12260
rect 51580 12220 51640 12260
rect 51680 12220 51700 12260
rect 51520 12200 51700 12220
rect 49520 12140 49600 12200
rect 49520 12100 49540 12140
rect 49580 12100 49600 12140
rect 49520 12080 49600 12100
rect 51520 12140 51600 12160
rect 51520 12100 51540 12140
rect 51580 12100 51600 12140
rect 51520 12080 51600 12100
rect 51000 11980 51080 12000
rect 51000 11940 51020 11980
rect 51060 11940 51080 11980
rect 51000 11920 51080 11940
rect 52120 11980 52200 12000
rect 52120 11940 52140 11980
rect 52180 11940 52200 11980
rect 52120 11920 52200 11940
rect 49920 11870 50000 11890
rect 49510 11830 49590 11850
rect 49510 11810 49530 11830
rect 49470 11790 49530 11810
rect 49570 11810 49590 11830
rect 49920 11830 49940 11870
rect 49980 11830 50000 11870
rect 49920 11810 50000 11830
rect 50170 11830 50250 11850
rect 50170 11810 50190 11830
rect 49570 11790 50190 11810
rect 50230 11810 50250 11830
rect 50650 11830 50730 11850
rect 50650 11810 50670 11830
rect 50230 11790 50290 11810
rect 49470 11770 50290 11790
rect 49470 11730 49510 11770
rect 49600 11730 49640 11770
rect 49860 11730 49900 11770
rect 50120 11730 50160 11770
rect 50250 11730 50290 11770
rect 50610 11790 50670 11810
rect 50710 11810 50730 11830
rect 51000 11810 51040 11920
rect 51310 11830 51390 11850
rect 51310 11810 51330 11830
rect 50710 11790 51330 11810
rect 51370 11810 51390 11830
rect 51790 11830 51870 11850
rect 51790 11810 51810 11830
rect 51370 11790 51430 11810
rect 50610 11770 51430 11790
rect 50610 11730 50650 11770
rect 50740 11730 50780 11770
rect 51000 11730 51040 11770
rect 51260 11730 51300 11770
rect 51390 11730 51430 11770
rect 51750 11790 51810 11810
rect 51850 11810 51870 11830
rect 52140 11810 52180 11920
rect 52450 11830 52530 11850
rect 52450 11810 52470 11830
rect 51850 11790 52470 11810
rect 52510 11810 52530 11830
rect 52510 11790 52570 11810
rect 51750 11770 52570 11790
rect 51750 11730 51790 11770
rect 51880 11730 51920 11770
rect 52140 11730 52180 11770
rect 52400 11730 52440 11770
rect 52530 11730 52570 11770
rect 49450 11710 49530 11730
rect 49450 11670 49470 11710
rect 49510 11670 49530 11710
rect 49450 11610 49530 11670
rect 49450 11570 49470 11610
rect 49510 11570 49530 11610
rect 49450 11550 49530 11570
rect 49580 11710 49660 11730
rect 49580 11670 49600 11710
rect 49640 11670 49660 11710
rect 49580 11610 49660 11670
rect 49580 11570 49600 11610
rect 49640 11570 49660 11610
rect 49580 11550 49660 11570
rect 49710 11710 49790 11730
rect 49710 11670 49730 11710
rect 49770 11670 49790 11710
rect 49710 11610 49790 11670
rect 49710 11570 49730 11610
rect 49770 11570 49790 11610
rect 49710 11550 49790 11570
rect 49840 11710 49920 11730
rect 49840 11670 49860 11710
rect 49900 11670 49920 11710
rect 49840 11610 49920 11670
rect 49840 11570 49860 11610
rect 49900 11570 49920 11610
rect 49840 11550 49920 11570
rect 49970 11710 50050 11730
rect 49970 11670 49990 11710
rect 50030 11670 50050 11710
rect 49970 11610 50050 11670
rect 49970 11570 49990 11610
rect 50030 11570 50050 11610
rect 49970 11550 50050 11570
rect 50100 11710 50190 11730
rect 50100 11670 50120 11710
rect 50160 11670 50190 11710
rect 50100 11610 50190 11670
rect 50100 11570 50120 11610
rect 50160 11570 50190 11610
rect 50100 11550 50190 11570
rect 50230 11710 50310 11730
rect 50230 11670 50250 11710
rect 50290 11670 50310 11710
rect 50230 11610 50310 11670
rect 50230 11570 50250 11610
rect 50290 11570 50310 11610
rect 50230 11550 50310 11570
rect 50490 11710 50670 11730
rect 50490 11670 50510 11710
rect 50550 11670 50610 11710
rect 50650 11670 50670 11710
rect 50490 11610 50670 11670
rect 50490 11570 50510 11610
rect 50550 11570 50610 11610
rect 50650 11570 50670 11610
rect 50490 11550 50670 11570
rect 50720 11710 50800 11730
rect 50720 11670 50740 11710
rect 50780 11670 50800 11710
rect 50720 11610 50800 11670
rect 50720 11570 50740 11610
rect 50780 11570 50800 11610
rect 50720 11550 50800 11570
rect 50850 11710 50930 11730
rect 50850 11670 50870 11710
rect 50910 11670 50930 11710
rect 50850 11610 50930 11670
rect 50850 11570 50870 11610
rect 50910 11570 50930 11610
rect 50850 11550 50930 11570
rect 50980 11710 51060 11730
rect 50980 11670 51000 11710
rect 51040 11670 51060 11710
rect 50980 11610 51060 11670
rect 50980 11570 51000 11610
rect 51040 11570 51060 11610
rect 50980 11550 51060 11570
rect 51110 11710 51190 11730
rect 51110 11670 51130 11710
rect 51170 11670 51190 11710
rect 51110 11610 51190 11670
rect 51110 11570 51130 11610
rect 51170 11570 51190 11610
rect 51110 11550 51190 11570
rect 51240 11710 51320 11730
rect 51240 11670 51260 11710
rect 51300 11670 51320 11710
rect 51240 11610 51320 11670
rect 51240 11570 51260 11610
rect 51300 11570 51320 11610
rect 51240 11550 51320 11570
rect 51370 11710 51550 11730
rect 51370 11670 51390 11710
rect 51430 11670 51490 11710
rect 51530 11670 51550 11710
rect 51370 11610 51550 11670
rect 51370 11570 51390 11610
rect 51430 11570 51490 11610
rect 51530 11570 51550 11610
rect 51370 11550 51550 11570
rect 51630 11710 51810 11730
rect 51630 11670 51650 11710
rect 51690 11670 51750 11710
rect 51790 11670 51810 11710
rect 51630 11610 51810 11670
rect 51630 11570 51650 11610
rect 51690 11570 51750 11610
rect 51790 11570 51810 11610
rect 51630 11550 51810 11570
rect 51860 11710 51940 11730
rect 51860 11670 51880 11710
rect 51920 11670 51940 11710
rect 51860 11610 51940 11670
rect 51860 11570 51880 11610
rect 51920 11570 51940 11610
rect 51860 11550 51940 11570
rect 51990 11710 52070 11730
rect 51990 11670 52010 11710
rect 52050 11670 52070 11710
rect 51990 11610 52070 11670
rect 51990 11570 52010 11610
rect 52050 11570 52070 11610
rect 51990 11550 52070 11570
rect 52120 11710 52200 11730
rect 52120 11670 52140 11710
rect 52180 11670 52200 11710
rect 52120 11610 52200 11670
rect 52120 11570 52140 11610
rect 52180 11570 52200 11610
rect 52120 11550 52200 11570
rect 52250 11710 52330 11730
rect 52250 11670 52270 11710
rect 52310 11670 52330 11710
rect 52250 11610 52330 11670
rect 52250 11570 52270 11610
rect 52310 11570 52330 11610
rect 52250 11550 52330 11570
rect 52380 11710 52460 11730
rect 52380 11670 52400 11710
rect 52440 11670 52460 11710
rect 52380 11610 52460 11670
rect 52380 11570 52400 11610
rect 52440 11570 52460 11610
rect 52380 11550 52460 11570
rect 52510 11710 52690 11730
rect 52510 11670 52530 11710
rect 52570 11670 52630 11710
rect 52670 11670 52690 11710
rect 52510 11610 52690 11670
rect 52510 11570 52530 11610
rect 52570 11570 52630 11610
rect 52670 11570 52690 11610
rect 52510 11550 52690 11570
rect 53067 13110 53090 13130
rect 49620 11490 49700 11510
rect 49620 11450 49640 11490
rect 49680 11450 49700 11490
rect 49620 11430 49700 11450
rect 50060 11490 50140 11510
rect 50060 11450 50080 11490
rect 50120 11450 50140 11490
rect 50060 11430 50140 11450
rect 50850 11480 50930 11500
rect 50850 11440 50870 11480
rect 50910 11440 50930 11480
rect 50850 11420 50930 11440
rect 51900 11490 51980 11510
rect 51900 11450 51920 11490
rect 51960 11450 51980 11490
rect 51900 11430 51980 11450
rect 52030 11340 52070 11550
rect 52250 11340 52290 11550
rect 52740 11490 52820 11510
rect 52740 11450 52760 11490
rect 52800 11450 52820 11490
rect 53033 11497 53067 11559
rect 53451 11497 53485 11559
rect 53033 11463 53129 11497
rect 53389 11463 53485 11497
rect 52740 11430 52820 11450
rect 52030 11320 52110 11340
rect 51900 11270 51980 11290
rect 51900 11230 51920 11270
rect 51960 11230 51980 11270
rect 51900 11210 51980 11230
rect 52030 11280 52050 11320
rect 52090 11280 52110 11320
rect 52030 11260 52110 11280
rect 52230 11320 52310 11340
rect 52230 11280 52250 11320
rect 52290 11280 52310 11320
rect 52230 11260 52310 11280
rect 53560 11320 53640 11340
rect 53560 11280 53580 11320
rect 53620 11280 53640 11320
rect 53560 11260 53640 11280
rect 49710 11150 49790 11170
rect 49710 11110 49730 11150
rect 49770 11110 49790 11150
rect 49710 11090 49790 11110
rect 50760 11150 50840 11170
rect 50760 11110 50780 11150
rect 50820 11110 50840 11150
rect 50760 11090 50840 11110
rect 51200 11150 51280 11170
rect 51200 11110 51220 11150
rect 51260 11110 51280 11150
rect 51200 11090 51280 11110
rect 52030 11050 52070 11260
rect 52250 11050 52290 11260
rect 52740 11150 52820 11170
rect 52740 11110 52760 11150
rect 52800 11110 52820 11150
rect 52740 11090 52820 11110
rect 53033 11101 53129 11135
rect 53389 11101 53485 11135
rect 49350 11030 49530 11050
rect 49350 10990 49370 11030
rect 49410 10990 49470 11030
rect 49510 10990 49530 11030
rect 49350 10970 49530 10990
rect 49580 11030 49660 11050
rect 49580 10990 49600 11030
rect 49640 10990 49660 11030
rect 49580 10970 49660 10990
rect 49710 11030 49790 11050
rect 49710 10990 49730 11030
rect 49770 10990 49790 11030
rect 49710 10970 49790 10990
rect 49840 11030 49920 11050
rect 49840 10990 49860 11030
rect 49900 10990 49920 11030
rect 49840 10970 49920 10990
rect 49970 11030 50050 11050
rect 49970 10990 49990 11030
rect 50030 10990 50050 11030
rect 49970 10970 50050 10990
rect 50100 11030 50180 11050
rect 50100 10990 50120 11030
rect 50160 10990 50180 11030
rect 50100 10970 50180 10990
rect 50230 11030 50410 11050
rect 50230 10990 50250 11030
rect 50290 10990 50350 11030
rect 50390 10990 50410 11030
rect 50230 10970 50410 10990
rect 50590 11030 50670 11050
rect 50590 10990 50610 11030
rect 50650 10990 50670 11030
rect 50590 10970 50670 10990
rect 50720 11030 50800 11050
rect 50720 10990 50740 11030
rect 50780 10990 50800 11030
rect 50720 10970 50800 10990
rect 50850 11030 50930 11050
rect 50850 10990 50870 11030
rect 50910 10990 50930 11030
rect 50850 10970 50930 10990
rect 50980 11030 51060 11050
rect 50980 10990 51000 11030
rect 51040 10990 51060 11030
rect 50980 10970 51060 10990
rect 51110 11030 51190 11050
rect 51110 10990 51130 11030
rect 51170 10990 51190 11030
rect 51110 10970 51190 10990
rect 51240 11030 51320 11050
rect 51240 10990 51260 11030
rect 51300 10990 51320 11030
rect 51240 10970 51320 10990
rect 51370 11030 51450 11050
rect 51370 10990 51390 11030
rect 51430 10990 51450 11030
rect 51370 10970 51450 10990
rect 51630 11030 51810 11050
rect 51630 10990 51650 11030
rect 51690 10990 51750 11030
rect 51790 10990 51810 11030
rect 51630 10970 51810 10990
rect 51860 11030 51940 11050
rect 51860 10990 51880 11030
rect 51920 10990 51940 11030
rect 51860 10970 51940 10990
rect 51990 11030 52070 11050
rect 51990 10990 52010 11030
rect 52050 10990 52070 11030
rect 51990 10970 52070 10990
rect 52120 11030 52200 11050
rect 52120 10990 52140 11030
rect 52180 10990 52200 11030
rect 52120 10970 52200 10990
rect 52250 11030 52330 11050
rect 52250 10990 52270 11030
rect 52310 10990 52330 11030
rect 52250 10970 52330 10990
rect 52380 11030 52460 11050
rect 52380 10990 52400 11030
rect 52440 10990 52460 11030
rect 52380 10970 52460 10990
rect 52510 11030 52690 11050
rect 52510 10990 52530 11030
rect 52570 10990 52630 11030
rect 52670 10990 52690 11030
rect 52510 10970 52690 10990
rect 53033 11039 53067 11101
rect 49470 10930 49510 10970
rect 49600 10930 49640 10970
rect 49860 10930 49900 10970
rect 50120 10930 50160 10970
rect 50250 10930 50290 10970
rect 49470 10910 50290 10930
rect 49470 10890 49530 10910
rect 49510 10860 49530 10890
rect 49580 10890 50180 10910
rect 49580 10860 49600 10890
rect 49510 10840 49600 10860
rect 49860 10780 49900 10890
rect 50160 10860 50180 10890
rect 50230 10890 50290 10910
rect 50610 10930 50650 10970
rect 50740 10930 50780 10970
rect 51000 10930 51040 10970
rect 51260 10930 51300 10970
rect 51390 10930 51430 10970
rect 50610 10910 51430 10930
rect 50610 10890 50670 10910
rect 50230 10860 50250 10890
rect 50160 10840 50250 10860
rect 50650 10870 50670 10890
rect 50710 10890 51330 10910
rect 50710 10870 50730 10890
rect 50650 10850 50730 10870
rect 50980 10870 51060 10890
rect 50980 10830 51000 10870
rect 51040 10830 51060 10870
rect 51310 10870 51330 10890
rect 51370 10890 51430 10910
rect 51750 10930 51790 10970
rect 51880 10930 51920 10970
rect 52140 10930 52180 10970
rect 52400 10930 52440 10970
rect 52530 10930 52570 10970
rect 51750 10910 52570 10930
rect 51370 10870 51390 10890
rect 51750 10880 51810 10910
rect 51310 10850 51390 10870
rect 51790 10870 51810 10880
rect 51850 10880 52470 10910
rect 51850 10870 51870 10880
rect 51790 10850 51870 10870
rect 50980 10810 51060 10830
rect 52140 10780 52180 10880
rect 52450 10870 52470 10880
rect 52510 10880 52570 10910
rect 52510 10870 52530 10880
rect 52450 10850 52530 10870
rect 49840 10760 49920 10780
rect 49840 10720 49860 10760
rect 49900 10720 49920 10760
rect 49840 10700 49920 10720
rect 52120 10760 52200 10780
rect 52120 10720 52140 10760
rect 52180 10720 52200 10760
rect 52120 10700 52200 10720
rect 50980 10650 51060 10670
rect 49400 10610 49480 10630
rect 49400 10570 49420 10610
rect 49460 10570 49480 10610
rect 50980 10610 51000 10650
rect 51040 10610 51060 10650
rect 50980 10590 51060 10610
rect 49400 10550 49480 10570
rect 49820 10550 51060 10590
rect 51400 10610 51480 10630
rect 51400 10570 51420 10610
rect 51460 10570 51480 10610
rect 51400 10550 51480 10570
rect 49420 10510 49460 10550
rect 49820 10510 49860 10550
rect 51020 10510 51060 10550
rect 51420 10510 51460 10550
rect 49300 10490 49480 10510
rect 49300 10440 49320 10490
rect 49360 10440 49420 10490
rect 49460 10440 49480 10490
rect 49300 10350 49480 10440
rect 49300 10300 49320 10350
rect 49360 10300 49420 10350
rect 49460 10300 49480 10350
rect 49300 10280 49480 10300
rect 49600 10490 49680 10510
rect 49600 10440 49620 10490
rect 49660 10440 49680 10490
rect 49600 10350 49680 10440
rect 49600 10300 49620 10350
rect 49660 10300 49680 10350
rect 49600 10280 49680 10300
rect 49800 10490 49880 10510
rect 49800 10440 49820 10490
rect 49860 10440 49880 10490
rect 49800 10350 49880 10440
rect 49800 10300 49820 10350
rect 49860 10300 49880 10350
rect 49800 10280 49880 10300
rect 50000 10490 50080 10510
rect 50000 10440 50020 10490
rect 50060 10440 50080 10490
rect 50000 10350 50080 10440
rect 50000 10300 50020 10350
rect 50060 10300 50080 10350
rect 50000 10280 50080 10300
rect 50200 10490 50280 10510
rect 50200 10440 50220 10490
rect 50260 10440 50280 10490
rect 50200 10350 50280 10440
rect 50200 10300 50220 10350
rect 50260 10300 50280 10350
rect 50200 10280 50280 10300
rect 50400 10490 50480 10510
rect 50400 10440 50420 10490
rect 50460 10440 50480 10490
rect 50400 10350 50480 10440
rect 50400 10300 50420 10350
rect 50460 10300 50480 10350
rect 50400 10280 50480 10300
rect 50600 10490 50680 10510
rect 50600 10440 50620 10490
rect 50660 10440 50680 10490
rect 50600 10350 50680 10440
rect 50600 10300 50620 10350
rect 50660 10300 50680 10350
rect 50600 10280 50680 10300
rect 50800 10490 50880 10510
rect 50800 10440 50820 10490
rect 50860 10440 50880 10490
rect 50800 10350 50880 10440
rect 50800 10300 50820 10350
rect 50860 10300 50880 10350
rect 50800 10280 50880 10300
rect 51000 10490 51080 10510
rect 51000 10440 51020 10490
rect 51060 10440 51080 10490
rect 51000 10350 51080 10440
rect 51000 10300 51020 10350
rect 51060 10300 51080 10350
rect 51000 10280 51080 10300
rect 51200 10490 51280 10510
rect 51200 10440 51220 10490
rect 51260 10440 51280 10490
rect 51200 10350 51280 10440
rect 51200 10300 51220 10350
rect 51260 10300 51280 10350
rect 51200 10280 51280 10300
rect 51400 10490 51580 10510
rect 51400 10440 51420 10490
rect 51460 10440 51520 10490
rect 51560 10440 51580 10490
rect 51400 10350 51580 10440
rect 51400 10300 51420 10350
rect 51460 10300 51520 10350
rect 51560 10300 51580 10350
rect 51400 10280 51580 10300
rect 50220 10240 50260 10280
rect 50620 10240 50660 10280
rect 50200 10220 50680 10240
rect 50200 10180 50220 10220
rect 50260 10180 50620 10220
rect 50660 10180 50680 10220
rect 50200 10160 50680 10180
rect 49140 10040 49260 10050
rect 50590 10040 50680 10160
rect 49140 10030 49294 10040
rect 49140 9990 49160 10030
rect 49200 10024 49294 10030
rect 49200 9990 49260 10024
rect 49140 9974 49294 9990
rect 50534 10024 50680 10040
rect 50568 9990 50680 10024
rect 50534 9974 50680 9990
rect 49140 9970 49260 9974
rect 50560 9970 50680 9974
rect 53010 9640 53033 9660
rect 53451 11039 53485 11101
rect 53067 9640 53090 9660
rect 53010 9600 53030 9640
rect 53070 9600 53090 9640
rect 53010 9580 53033 9600
rect 53067 9580 53090 9600
rect 53033 9227 53067 9289
rect 53451 9227 53485 9289
rect 53033 9193 53129 9227
rect 53389 9193 53485 9227
<< viali >>
rect 53240 13510 53278 13598
rect 53230 13450 53290 13510
rect 53240 13201 53278 13450
rect 53030 13130 53033 13170
rect 53033 13130 53067 13170
rect 53067 13130 53070 13170
rect 50340 12740 50380 12780
rect 50740 12740 50780 12780
rect 49540 12620 49580 12660
rect 49540 12520 49580 12560
rect 49540 12420 49580 12460
rect 49540 12320 49580 12360
rect 49540 12220 49580 12260
rect 49740 12620 49780 12660
rect 49740 12520 49780 12560
rect 49740 12420 49780 12460
rect 49740 12320 49780 12360
rect 49740 12220 49780 12260
rect 49940 12620 49980 12660
rect 49940 12520 49980 12560
rect 49940 12420 49980 12460
rect 49940 12320 49980 12360
rect 49940 12220 49980 12260
rect 50140 12620 50180 12660
rect 50140 12520 50180 12560
rect 50140 12420 50180 12460
rect 50140 12320 50180 12360
rect 50140 12220 50180 12260
rect 50340 12620 50380 12660
rect 50340 12520 50380 12560
rect 50340 12420 50380 12460
rect 50340 12320 50380 12360
rect 50340 12220 50380 12260
rect 50540 12620 50580 12660
rect 50540 12520 50580 12560
rect 50540 12420 50580 12460
rect 50540 12320 50580 12360
rect 50540 12220 50580 12260
rect 50740 12620 50780 12660
rect 50740 12520 50780 12560
rect 50740 12420 50780 12460
rect 50740 12320 50780 12360
rect 50740 12220 50780 12260
rect 50940 12620 50980 12660
rect 50940 12520 50980 12560
rect 50940 12420 50980 12460
rect 50940 12320 50980 12360
rect 50940 12220 50980 12260
rect 51140 12620 51180 12660
rect 51140 12520 51180 12560
rect 51140 12420 51180 12460
rect 51140 12320 51180 12360
rect 51140 12220 51180 12260
rect 51340 12620 51380 12660
rect 51340 12520 51380 12560
rect 51340 12420 51380 12460
rect 51340 12320 51380 12360
rect 51340 12220 51380 12260
rect 51540 12620 51580 12660
rect 51540 12520 51580 12560
rect 51540 12420 51580 12460
rect 51540 12320 51580 12360
rect 51540 12220 51580 12260
rect 49540 12100 49580 12140
rect 51540 12100 51580 12140
rect 51020 11940 51060 11980
rect 52140 11940 52180 11980
rect 49940 11830 49980 11870
rect 49470 11670 49510 11710
rect 49470 11570 49510 11610
rect 49600 11670 49640 11710
rect 49600 11570 49640 11610
rect 49730 11670 49770 11710
rect 49730 11570 49770 11610
rect 49860 11670 49900 11710
rect 49860 11570 49900 11610
rect 49990 11670 50030 11710
rect 49990 11570 50030 11610
rect 50120 11670 50160 11710
rect 50120 11570 50160 11610
rect 50250 11670 50290 11710
rect 50250 11570 50290 11610
rect 50610 11670 50650 11710
rect 50610 11570 50650 11610
rect 50740 11670 50780 11710
rect 50740 11570 50780 11610
rect 50870 11670 50910 11710
rect 50870 11570 50910 11610
rect 51000 11670 51040 11710
rect 51000 11570 51040 11610
rect 51130 11670 51170 11710
rect 51130 11570 51170 11610
rect 51260 11670 51300 11710
rect 51260 11570 51300 11610
rect 51390 11670 51430 11710
rect 51390 11570 51430 11610
rect 53230 11610 53290 12020
rect 49640 11450 49680 11490
rect 50080 11450 50120 11490
rect 50870 11440 50910 11480
rect 51920 11450 51960 11490
rect 52760 11450 52800 11490
rect 51920 11230 51960 11270
rect 52050 11280 52090 11320
rect 52250 11280 52290 11320
rect 53580 11280 53620 11320
rect 49730 11110 49770 11150
rect 50780 11110 50820 11150
rect 51220 11110 51260 11150
rect 52760 11110 52800 11150
rect 49470 10990 49510 11030
rect 49600 10990 49640 11030
rect 49730 10990 49770 11030
rect 49860 10990 49900 11030
rect 49990 10990 50030 11030
rect 50120 10990 50160 11030
rect 50250 10990 50290 11030
rect 50610 10990 50650 11030
rect 50740 10990 50780 11030
rect 50870 10990 50910 11030
rect 51000 10990 51040 11030
rect 51130 10990 51170 11030
rect 51260 10990 51300 11030
rect 51390 10990 51430 11030
rect 51000 10830 51040 10870
rect 49860 10720 49900 10760
rect 52140 10720 52180 10760
rect 49420 10570 49460 10610
rect 51000 10610 51040 10650
rect 51420 10570 51460 10610
rect 49620 10440 49660 10490
rect 49620 10300 49660 10350
rect 50020 10440 50060 10490
rect 50020 10300 50060 10350
rect 50420 10440 50460 10490
rect 50420 10300 50460 10350
rect 50820 10440 50860 10490
rect 50820 10300 50860 10350
rect 51220 10440 51260 10490
rect 51220 10300 51260 10350
rect 49160 9990 49200 10030
rect 53230 10590 53290 10980
rect 53030 9600 53033 9640
rect 53033 9600 53067 9640
rect 53067 9600 53070 9640
rect 53240 9350 53278 9747
<< metal1 >>
rect 53234 13598 53284 13610
rect 53234 13530 53240 13598
rect 53210 13510 53240 13530
rect 53278 13530 53284 13598
rect 53278 13510 53310 13530
rect 53210 13450 53230 13510
rect 53290 13450 53310 13510
rect 53210 13430 53240 13450
rect 53234 13201 53240 13430
rect 53278 13430 53310 13450
rect 53278 13201 53284 13430
rect 53010 13180 53090 13190
rect 53234 13189 53284 13201
rect 53010 13120 53020 13180
rect 53080 13120 53090 13180
rect 53010 13110 53090 13120
rect 49140 12790 49220 12800
rect 49140 12730 49150 12790
rect 49210 12730 49220 12790
rect 49030 11410 49110 11420
rect 49030 11350 49040 11410
rect 49100 11350 49110 11410
rect 49030 11340 49110 11350
rect 48920 11250 49000 11260
rect 48920 11190 48930 11250
rect 48990 11190 49000 11250
rect 48920 11180 49000 11190
rect 49140 10030 49220 12730
rect 50320 12790 50400 12800
rect 50320 12730 50330 12790
rect 50390 12730 50400 12790
rect 49520 12660 49600 12680
rect 49520 12620 49540 12660
rect 49580 12620 49600 12660
rect 49520 12560 49600 12620
rect 49520 12520 49540 12560
rect 49580 12520 49600 12560
rect 49520 12460 49600 12520
rect 49520 12420 49540 12460
rect 49580 12420 49600 12460
rect 49520 12360 49600 12420
rect 49520 12320 49540 12360
rect 49580 12320 49600 12360
rect 49520 12260 49600 12320
rect 49520 12220 49540 12260
rect 49580 12220 49600 12260
rect 49520 12200 49600 12220
rect 49720 12660 49800 12680
rect 49720 12620 49740 12660
rect 49780 12620 49800 12660
rect 49720 12560 49800 12620
rect 49720 12520 49740 12560
rect 49780 12520 49800 12560
rect 49720 12460 49800 12520
rect 49720 12420 49740 12460
rect 49780 12420 49800 12460
rect 49720 12360 49800 12420
rect 49720 12320 49740 12360
rect 49780 12320 49800 12360
rect 49720 12260 49800 12320
rect 49720 12220 49740 12260
rect 49780 12220 49800 12260
rect 49520 12140 49600 12160
rect 49520 12100 49540 12140
rect 49580 12100 49600 12140
rect 49520 11990 49600 12100
rect 49520 11930 49530 11990
rect 49590 11930 49600 11990
rect 49520 11920 49600 11930
rect 49720 11990 49800 12220
rect 49720 11930 49730 11990
rect 49790 11930 49800 11990
rect 49720 11920 49800 11930
rect 49920 12660 50000 12680
rect 49920 12620 49940 12660
rect 49980 12620 50000 12660
rect 49920 12560 50000 12620
rect 49920 12520 49940 12560
rect 49980 12520 50000 12560
rect 49920 12460 50000 12520
rect 49920 12420 49940 12460
rect 49980 12420 50000 12460
rect 49920 12360 50000 12420
rect 49920 12320 49940 12360
rect 49980 12320 50000 12360
rect 49920 12260 50000 12320
rect 49920 12220 49940 12260
rect 49980 12220 50000 12260
rect 49920 12130 50000 12220
rect 49920 12070 49930 12130
rect 49990 12070 50000 12130
rect 49920 11880 50000 12070
rect 50120 12660 50200 12680
rect 50120 12620 50140 12660
rect 50180 12620 50200 12660
rect 50120 12560 50200 12620
rect 50120 12520 50140 12560
rect 50180 12520 50200 12560
rect 50120 12460 50200 12520
rect 50120 12420 50140 12460
rect 50180 12420 50200 12460
rect 50120 12360 50200 12420
rect 50120 12320 50140 12360
rect 50180 12320 50200 12360
rect 50120 12260 50200 12320
rect 50120 12220 50140 12260
rect 50180 12220 50200 12260
rect 50120 11990 50200 12220
rect 50320 12660 50400 12730
rect 50720 12790 50800 12800
rect 50720 12730 50730 12790
rect 50790 12730 50800 12790
rect 50320 12620 50340 12660
rect 50380 12620 50400 12660
rect 50320 12560 50400 12620
rect 50320 12520 50340 12560
rect 50380 12520 50400 12560
rect 50320 12460 50400 12520
rect 50320 12420 50340 12460
rect 50380 12420 50400 12460
rect 50320 12360 50400 12420
rect 50320 12320 50340 12360
rect 50380 12320 50400 12360
rect 50320 12260 50400 12320
rect 50320 12220 50340 12260
rect 50380 12220 50400 12260
rect 50320 12200 50400 12220
rect 50520 12660 50600 12680
rect 50520 12620 50540 12660
rect 50580 12620 50600 12660
rect 50520 12560 50600 12620
rect 50520 12520 50540 12560
rect 50580 12520 50600 12560
rect 50520 12460 50600 12520
rect 50520 12420 50540 12460
rect 50580 12420 50600 12460
rect 50520 12360 50600 12420
rect 50520 12320 50540 12360
rect 50580 12320 50600 12360
rect 50520 12260 50600 12320
rect 50520 12220 50540 12260
rect 50580 12220 50600 12260
rect 50120 11930 50130 11990
rect 50190 11930 50200 11990
rect 50120 11920 50200 11930
rect 50520 11990 50600 12220
rect 50720 12660 50800 12730
rect 50720 12620 50740 12660
rect 50780 12620 50800 12660
rect 50720 12560 50800 12620
rect 50720 12520 50740 12560
rect 50780 12520 50800 12560
rect 50720 12460 50800 12520
rect 50720 12420 50740 12460
rect 50780 12420 50800 12460
rect 50720 12360 50800 12420
rect 50720 12320 50740 12360
rect 50780 12320 50800 12360
rect 50720 12260 50800 12320
rect 50720 12220 50740 12260
rect 50780 12220 50800 12260
rect 50720 12200 50800 12220
rect 50920 12660 51000 12680
rect 50920 12620 50940 12660
rect 50980 12620 51000 12660
rect 50920 12560 51000 12620
rect 50920 12520 50940 12560
rect 50980 12520 51000 12560
rect 50920 12460 51000 12520
rect 50920 12420 50940 12460
rect 50980 12420 51000 12460
rect 50920 12360 51000 12420
rect 50920 12320 50940 12360
rect 50980 12320 51000 12360
rect 50920 12260 51000 12320
rect 50920 12220 50940 12260
rect 50980 12220 51000 12260
rect 50520 11930 50530 11990
rect 50590 11930 50600 11990
rect 50520 11920 50600 11930
rect 50920 12000 51000 12220
rect 51120 12660 51200 12680
rect 51120 12620 51140 12660
rect 51180 12620 51200 12660
rect 51120 12560 51200 12620
rect 51120 12520 51140 12560
rect 51180 12520 51200 12560
rect 51120 12460 51200 12520
rect 51120 12420 51140 12460
rect 51180 12420 51200 12460
rect 51120 12360 51200 12420
rect 51120 12320 51140 12360
rect 51180 12320 51200 12360
rect 51120 12260 51200 12320
rect 51120 12220 51140 12260
rect 51180 12220 51200 12260
rect 51120 12130 51200 12220
rect 51120 12070 51130 12130
rect 51190 12070 51200 12130
rect 51120 12060 51200 12070
rect 51320 12660 51400 12680
rect 51320 12620 51340 12660
rect 51380 12620 51400 12660
rect 51320 12560 51400 12620
rect 51320 12520 51340 12560
rect 51380 12520 51400 12560
rect 51320 12460 51400 12520
rect 51320 12420 51340 12460
rect 51380 12420 51400 12460
rect 51320 12360 51400 12420
rect 51320 12320 51340 12360
rect 51380 12320 51400 12360
rect 51320 12260 51400 12320
rect 51320 12220 51340 12260
rect 51380 12220 51400 12260
rect 50920 11990 51080 12000
rect 50920 11930 50930 11990
rect 50990 11930 51010 11990
rect 51070 11930 51080 11990
rect 50920 11920 51080 11930
rect 51320 11990 51400 12220
rect 51320 11930 51330 11990
rect 51390 11930 51400 11990
rect 51320 11920 51400 11930
rect 51520 12660 51600 12680
rect 51520 12620 51540 12660
rect 51580 12620 51600 12660
rect 51520 12560 51600 12620
rect 51520 12520 51540 12560
rect 51580 12520 51600 12560
rect 51520 12460 51600 12520
rect 51520 12420 51540 12460
rect 51580 12420 51600 12460
rect 51520 12360 51600 12420
rect 51520 12320 51540 12360
rect 51580 12320 51600 12360
rect 51520 12260 51600 12320
rect 51520 12220 51540 12260
rect 51580 12220 51600 12260
rect 51520 12140 51600 12220
rect 51520 12100 51540 12140
rect 51580 12100 51600 12140
rect 51520 11990 51600 12100
rect 53220 12020 53300 12040
rect 51520 11930 51530 11990
rect 51590 11930 51600 11990
rect 51520 11920 51600 11930
rect 52120 11990 52200 12000
rect 52120 11930 52130 11990
rect 52190 11930 52200 11990
rect 52120 11920 52200 11930
rect 49920 11820 49930 11880
rect 49990 11820 50000 11880
rect 49920 11810 50000 11820
rect 49450 11710 49530 11730
rect 49450 11670 49470 11710
rect 49510 11670 49530 11710
rect 49450 11610 49530 11670
rect 49450 11570 49470 11610
rect 49510 11570 49530 11610
rect 49450 11550 49530 11570
rect 49580 11710 49660 11730
rect 49580 11670 49600 11710
rect 49640 11670 49660 11710
rect 49580 11610 49660 11670
rect 49580 11570 49600 11610
rect 49640 11570 49660 11610
rect 49580 11550 49660 11570
rect 49710 11710 49790 11730
rect 49710 11670 49730 11710
rect 49770 11670 49790 11710
rect 49710 11610 49790 11670
rect 49710 11570 49730 11610
rect 49770 11570 49790 11610
rect 49710 11550 49790 11570
rect 49840 11710 49920 11730
rect 49840 11670 49860 11710
rect 49900 11670 49920 11710
rect 49840 11610 49920 11670
rect 49840 11570 49860 11610
rect 49900 11570 49920 11610
rect 49840 11550 49920 11570
rect 49970 11710 50050 11730
rect 49970 11670 49990 11710
rect 50030 11670 50050 11710
rect 49970 11610 50050 11670
rect 49970 11570 49990 11610
rect 50030 11570 50050 11610
rect 49970 11550 50050 11570
rect 50100 11710 50180 11730
rect 50100 11670 50120 11710
rect 50160 11670 50180 11710
rect 50100 11610 50180 11670
rect 50100 11570 50120 11610
rect 50160 11570 50180 11610
rect 50100 11550 50180 11570
rect 50230 11710 50310 11730
rect 50230 11670 50250 11710
rect 50290 11670 50310 11710
rect 50230 11610 50310 11670
rect 50230 11570 50250 11610
rect 50290 11570 50310 11610
rect 50230 11550 50310 11570
rect 50590 11710 50670 11730
rect 50590 11670 50610 11710
rect 50650 11670 50670 11710
rect 50590 11610 50670 11670
rect 50590 11570 50610 11610
rect 50650 11570 50670 11610
rect 50590 11550 50670 11570
rect 50720 11710 50800 11730
rect 50720 11670 50740 11710
rect 50780 11670 50800 11710
rect 50720 11610 50800 11670
rect 50720 11570 50740 11610
rect 50780 11570 50800 11610
rect 50720 11550 50800 11570
rect 50850 11710 50930 11730
rect 50850 11670 50870 11710
rect 50910 11670 50930 11710
rect 50850 11610 50930 11670
rect 50850 11570 50870 11610
rect 50910 11570 50930 11610
rect 49620 11500 49700 11510
rect 49620 11440 49630 11500
rect 49690 11440 49700 11500
rect 49620 11430 49700 11440
rect 49730 11170 49770 11550
rect 49990 11330 50030 11550
rect 50060 11500 50140 11510
rect 50060 11440 50070 11500
rect 50130 11440 50140 11500
rect 50060 11430 50140 11440
rect 50850 11480 50930 11570
rect 50980 11710 51060 11730
rect 50980 11670 51000 11710
rect 51040 11670 51060 11710
rect 50980 11610 51060 11670
rect 50980 11570 51000 11610
rect 51040 11570 51060 11610
rect 50980 11550 51060 11570
rect 51110 11710 51190 11730
rect 51110 11670 51130 11710
rect 51170 11670 51190 11710
rect 51110 11610 51190 11670
rect 51110 11570 51130 11610
rect 51170 11570 51190 11610
rect 51110 11550 51190 11570
rect 51240 11710 51320 11730
rect 51240 11670 51260 11710
rect 51300 11670 51320 11710
rect 51240 11610 51320 11670
rect 51240 11570 51260 11610
rect 51300 11570 51320 11610
rect 51240 11550 51320 11570
rect 51370 11710 51450 11730
rect 51370 11670 51390 11710
rect 51430 11670 51450 11710
rect 51370 11610 51450 11670
rect 51370 11570 51390 11610
rect 51430 11570 51450 11610
rect 51370 11550 51450 11570
rect 53220 11610 53230 12020
rect 53290 11610 53300 12020
rect 50850 11440 50870 11480
rect 50910 11440 50930 11480
rect 49970 11270 49980 11330
rect 50040 11270 50050 11330
rect 49710 11150 49790 11170
rect 49710 11110 49730 11150
rect 49770 11110 49790 11150
rect 49450 11030 49530 11050
rect 49450 10990 49470 11030
rect 49510 10990 49530 11030
rect 49450 10970 49530 10990
rect 49580 11030 49660 11050
rect 49580 10990 49600 11030
rect 49640 10990 49660 11030
rect 49580 10970 49660 10990
rect 49710 11030 49790 11110
rect 49990 11090 50030 11270
rect 50080 11240 50120 11430
rect 50850 11420 50930 11440
rect 51130 11490 51170 11550
rect 51900 11500 51980 11510
rect 51130 11480 51210 11490
rect 51130 11420 51140 11480
rect 51200 11420 51210 11480
rect 51900 11440 51910 11500
rect 51970 11440 51980 11500
rect 51900 11430 51980 11440
rect 52740 11500 52820 11510
rect 52740 11440 52750 11500
rect 52810 11440 52820 11500
rect 52740 11430 52820 11440
rect 53220 11500 53300 11610
rect 53220 11440 53230 11500
rect 53290 11440 53300 11500
rect 53220 11430 53300 11440
rect 53540 11580 53650 11600
rect 53540 11510 53560 11580
rect 53630 11510 53650 11580
rect 50720 11350 50730 11410
rect 50790 11350 50800 11410
rect 50060 11230 50140 11240
rect 50060 11170 50070 11230
rect 50130 11170 50140 11230
rect 50060 11160 50140 11170
rect 50760 11170 50800 11350
rect 50760 11160 50840 11170
rect 50760 11100 50770 11160
rect 50830 11100 50840 11160
rect 50760 11090 50840 11100
rect 49710 10990 49730 11030
rect 49770 10990 49790 11030
rect 49710 10970 49790 10990
rect 49840 11030 49920 11050
rect 49840 10990 49860 11030
rect 49900 10990 49920 11030
rect 49840 10970 49920 10990
rect 49970 11030 50050 11090
rect 50870 11050 50910 11420
rect 51130 11410 51210 11420
rect 51130 11050 51170 11410
rect 52030 11330 52110 11340
rect 51900 11280 51980 11290
rect 51900 11220 51910 11280
rect 51970 11220 51980 11280
rect 52030 11270 52040 11330
rect 52100 11270 52110 11330
rect 52030 11260 52110 11270
rect 52230 11330 52310 11340
rect 52230 11270 52240 11330
rect 52300 11270 52310 11330
rect 52230 11260 52310 11270
rect 53540 11330 53650 11510
rect 53540 11270 53570 11330
rect 53630 11270 53650 11330
rect 51900 11210 51980 11220
rect 51200 11160 51280 11170
rect 51200 11100 51210 11160
rect 51270 11100 51280 11160
rect 51200 11090 51280 11100
rect 52740 11160 52820 11170
rect 52740 11100 52750 11160
rect 52810 11100 52820 11160
rect 52740 11090 52820 11100
rect 53220 11160 53300 11170
rect 53220 11100 53230 11160
rect 53290 11100 53300 11160
rect 49970 10990 49990 11030
rect 50030 10990 50050 11030
rect 49970 10970 50050 10990
rect 50100 11030 50180 11050
rect 50100 10990 50120 11030
rect 50160 10990 50180 11030
rect 50100 10970 50180 10990
rect 50230 11030 50310 11050
rect 50230 10990 50250 11030
rect 50290 10990 50310 11030
rect 50230 10970 50310 10990
rect 50590 11030 50670 11050
rect 50590 10990 50610 11030
rect 50650 10990 50670 11030
rect 50590 10970 50670 10990
rect 50720 11030 50800 11050
rect 50720 10990 50740 11030
rect 50780 10990 50800 11030
rect 50720 10970 50800 10990
rect 50850 11030 50930 11050
rect 50850 10990 50870 11030
rect 50910 10990 50930 11030
rect 50850 10970 50930 10990
rect 50980 11030 51060 11050
rect 50980 10990 51000 11030
rect 51040 10990 51060 11030
rect 50980 10970 51060 10990
rect 51110 11030 51190 11050
rect 51110 10990 51130 11030
rect 51170 10990 51190 11030
rect 51110 10970 51190 10990
rect 51240 11030 51320 11050
rect 51240 10990 51260 11030
rect 51300 10990 51320 11030
rect 51240 10970 51320 10990
rect 51370 11030 51450 11050
rect 51370 10990 51390 11030
rect 51430 10990 51450 11030
rect 51370 10970 51450 10990
rect 53220 10980 53300 11100
rect 53540 11070 53650 11270
rect 53540 11000 53560 11070
rect 53630 11000 53650 11070
rect 53540 10980 53650 11000
rect 50980 10880 51060 10890
rect 50980 10820 50990 10880
rect 51050 10820 51060 10880
rect 49400 10770 49480 10780
rect 49400 10710 49410 10770
rect 49470 10710 49480 10770
rect 49400 10610 49480 10710
rect 49400 10570 49420 10610
rect 49460 10570 49480 10610
rect 49400 10550 49480 10570
rect 49600 10770 49680 10780
rect 49600 10710 49610 10770
rect 49670 10710 49680 10770
rect 49600 10490 49680 10710
rect 49840 10770 49920 10780
rect 49840 10710 49850 10770
rect 49910 10710 49920 10770
rect 49840 10700 49920 10710
rect 50000 10770 50080 10780
rect 50000 10710 50010 10770
rect 50070 10710 50080 10770
rect 49600 10440 49620 10490
rect 49660 10440 49680 10490
rect 49600 10350 49680 10440
rect 49600 10300 49620 10350
rect 49660 10300 49680 10350
rect 49600 10280 49680 10300
rect 50000 10490 50080 10710
rect 50000 10440 50020 10490
rect 50060 10440 50080 10490
rect 50000 10350 50080 10440
rect 50000 10300 50020 10350
rect 50060 10300 50080 10350
rect 50000 10280 50080 10300
rect 50400 10770 50480 10780
rect 50400 10710 50410 10770
rect 50470 10710 50480 10770
rect 50400 10490 50480 10710
rect 50400 10440 50420 10490
rect 50460 10440 50480 10490
rect 50400 10350 50480 10440
rect 50400 10300 50420 10350
rect 50460 10300 50480 10350
rect 50400 10280 50480 10300
rect 50800 10770 50880 10780
rect 50800 10710 50810 10770
rect 50870 10710 50880 10770
rect 50800 10490 50880 10710
rect 50980 10660 51060 10820
rect 50980 10600 50990 10660
rect 51050 10600 51060 10660
rect 50980 10590 51060 10600
rect 51200 10770 51280 10780
rect 51200 10710 51210 10770
rect 51270 10710 51280 10770
rect 50800 10440 50820 10490
rect 50860 10440 50880 10490
rect 50800 10350 50880 10440
rect 50800 10300 50820 10350
rect 50860 10300 50880 10350
rect 50800 10280 50880 10300
rect 51200 10490 51280 10710
rect 51400 10770 51480 10780
rect 51400 10710 51410 10770
rect 51470 10710 51480 10770
rect 51400 10610 51480 10710
rect 52120 10770 52200 10780
rect 52120 10710 52130 10770
rect 52190 10710 52200 10770
rect 52120 10700 52200 10710
rect 51400 10570 51420 10610
rect 51460 10570 51480 10610
rect 53220 10590 53230 10980
rect 53290 10590 53300 10980
rect 53220 10570 53300 10590
rect 51400 10550 51480 10570
rect 53234 10569 53284 10570
rect 51200 10440 51220 10490
rect 51260 10440 51280 10490
rect 51200 10350 51280 10440
rect 51200 10300 51220 10350
rect 51260 10300 51280 10350
rect 51200 10280 51280 10300
rect 49140 9990 49160 10030
rect 49200 9990 49220 10030
rect 49140 9970 49220 9990
rect 53210 9747 53310 9760
rect 53010 9650 53090 9660
rect 53010 9590 53020 9650
rect 53080 9590 53090 9650
rect 53010 9580 53090 9590
rect 53210 9350 53240 9747
rect 53278 9350 53310 9747
rect 53210 9140 53310 9350
rect 53210 9080 53230 9140
rect 53290 9080 53310 9140
rect 53210 9060 53310 9080
<< via1 >>
rect 53230 13450 53290 13510
rect 53020 13170 53080 13180
rect 53020 13130 53030 13170
rect 53030 13130 53070 13170
rect 53070 13130 53080 13170
rect 53020 13120 53080 13130
rect 49150 12730 49210 12790
rect 49040 11350 49100 11410
rect 48930 11190 48990 11250
rect 50330 12780 50390 12790
rect 50330 12740 50340 12780
rect 50340 12740 50380 12780
rect 50380 12740 50390 12780
rect 50330 12730 50390 12740
rect 49530 11930 49590 11990
rect 49730 11930 49790 11990
rect 49930 12070 49990 12130
rect 50730 12780 50790 12790
rect 50730 12740 50740 12780
rect 50740 12740 50780 12780
rect 50780 12740 50790 12780
rect 50730 12730 50790 12740
rect 50130 11930 50190 11990
rect 50530 11930 50590 11990
rect 51130 12070 51190 12130
rect 50930 11930 50990 11990
rect 51010 11980 51070 11990
rect 51010 11940 51020 11980
rect 51020 11940 51060 11980
rect 51060 11940 51070 11980
rect 51010 11930 51070 11940
rect 51330 11930 51390 11990
rect 51530 11930 51590 11990
rect 52130 11980 52190 11990
rect 52130 11940 52140 11980
rect 52140 11940 52180 11980
rect 52180 11940 52190 11980
rect 52130 11930 52190 11940
rect 49930 11870 49990 11880
rect 49930 11830 49940 11870
rect 49940 11830 49980 11870
rect 49980 11830 49990 11870
rect 49930 11820 49990 11830
rect 49630 11490 49690 11500
rect 49630 11450 49640 11490
rect 49640 11450 49680 11490
rect 49680 11450 49690 11490
rect 49630 11440 49690 11450
rect 50070 11490 50130 11500
rect 50070 11450 50080 11490
rect 50080 11450 50120 11490
rect 50120 11450 50130 11490
rect 50070 11440 50130 11450
rect 49980 11270 50040 11330
rect 51140 11420 51200 11480
rect 51910 11490 51970 11500
rect 51910 11450 51920 11490
rect 51920 11450 51960 11490
rect 51960 11450 51970 11490
rect 51910 11440 51970 11450
rect 52750 11490 52810 11500
rect 52750 11450 52760 11490
rect 52760 11450 52800 11490
rect 52800 11450 52810 11490
rect 52750 11440 52810 11450
rect 53230 11440 53290 11500
rect 53560 11510 53630 11580
rect 50730 11350 50790 11410
rect 50070 11170 50130 11230
rect 50770 11150 50830 11160
rect 50770 11110 50780 11150
rect 50780 11110 50820 11150
rect 50820 11110 50830 11150
rect 50770 11100 50830 11110
rect 51910 11270 51970 11280
rect 51910 11230 51920 11270
rect 51920 11230 51960 11270
rect 51960 11230 51970 11270
rect 51910 11220 51970 11230
rect 52040 11320 52100 11330
rect 52040 11280 52050 11320
rect 52050 11280 52090 11320
rect 52090 11280 52100 11320
rect 52040 11270 52100 11280
rect 52240 11320 52300 11330
rect 52240 11280 52250 11320
rect 52250 11280 52290 11320
rect 52290 11280 52300 11320
rect 52240 11270 52300 11280
rect 53570 11320 53630 11330
rect 53570 11280 53580 11320
rect 53580 11280 53620 11320
rect 53620 11280 53630 11320
rect 53570 11270 53630 11280
rect 51210 11150 51270 11160
rect 51210 11110 51220 11150
rect 51220 11110 51260 11150
rect 51260 11110 51270 11150
rect 51210 11100 51270 11110
rect 52750 11150 52810 11160
rect 52750 11110 52760 11150
rect 52760 11110 52800 11150
rect 52800 11110 52810 11150
rect 52750 11100 52810 11110
rect 53230 11100 53290 11160
rect 53560 11000 53630 11070
rect 50990 10870 51050 10880
rect 50990 10830 51000 10870
rect 51000 10830 51040 10870
rect 51040 10830 51050 10870
rect 50990 10820 51050 10830
rect 49410 10710 49470 10770
rect 49610 10710 49670 10770
rect 49850 10760 49910 10770
rect 49850 10720 49860 10760
rect 49860 10720 49900 10760
rect 49900 10720 49910 10760
rect 49850 10710 49910 10720
rect 50010 10710 50070 10770
rect 50410 10710 50470 10770
rect 50810 10710 50870 10770
rect 50990 10650 51050 10660
rect 50990 10610 51000 10650
rect 51000 10610 51040 10650
rect 51040 10610 51050 10650
rect 50990 10600 51050 10610
rect 51210 10710 51270 10770
rect 51410 10710 51470 10770
rect 52130 10760 52190 10770
rect 52130 10720 52140 10760
rect 52140 10720 52180 10760
rect 52180 10720 52190 10760
rect 52130 10710 52190 10720
rect 53020 9640 53080 9650
rect 53020 9600 53030 9640
rect 53030 9600 53070 9640
rect 53070 9600 53080 9640
rect 53020 9590 53080 9600
rect 53230 9080 53290 9140
<< metal2 >>
rect 53210 13510 53310 13530
rect 53210 13450 53230 13510
rect 53290 13450 53310 13510
rect 53210 13430 53310 13450
rect 48790 13180 53090 13190
rect 48790 13120 53020 13180
rect 53080 13120 53090 13180
rect 48790 13110 53090 13120
rect 49140 12790 50800 12800
rect 49140 12730 49150 12790
rect 49210 12730 50330 12790
rect 50390 12730 50730 12790
rect 50790 12730 50800 12790
rect 49140 12720 50800 12730
rect 49920 12130 51200 12140
rect 49920 12070 49930 12130
rect 49990 12070 51130 12130
rect 51190 12070 51200 12130
rect 49920 12060 51200 12070
rect 48790 11990 52200 12000
rect 48790 11930 49530 11990
rect 49590 11930 49730 11990
rect 49790 11930 50130 11990
rect 50190 11930 50530 11990
rect 50590 11930 50930 11990
rect 50990 11930 51010 11990
rect 51070 11930 51330 11990
rect 51390 11930 51530 11990
rect 51590 11930 52130 11990
rect 52190 11930 52200 11990
rect 48790 11920 52200 11930
rect 49920 11880 50000 11890
rect 49920 11820 49930 11880
rect 49990 11820 50000 11880
rect 49920 11810 50000 11820
rect 53540 11580 53650 11600
rect 53540 11510 53560 11580
rect 53630 11510 53650 11580
rect 49620 11500 49700 11510
rect 49620 11440 49630 11500
rect 49690 11440 49700 11500
rect 49030 11410 49110 11420
rect 49030 11350 49040 11410
rect 49100 11400 49110 11410
rect 49620 11400 49700 11440
rect 50060 11500 50140 11510
rect 50060 11440 50070 11500
rect 50130 11440 50140 11500
rect 51900 11500 51980 11510
rect 50060 11430 50140 11440
rect 51130 11480 51210 11490
rect 51130 11420 51140 11480
rect 51200 11470 51210 11480
rect 51900 11470 51910 11500
rect 51200 11440 51910 11470
rect 51970 11440 51980 11500
rect 51200 11430 51980 11440
rect 52740 11500 53300 11510
rect 52740 11440 52750 11500
rect 52810 11440 53230 11500
rect 53290 11440 53300 11500
rect 53540 11490 53650 11510
rect 52740 11430 53300 11440
rect 51200 11420 51210 11430
rect 51130 11410 51210 11420
rect 50720 11400 50730 11410
rect 49100 11360 50730 11400
rect 49100 11350 49110 11360
rect 50720 11350 50730 11360
rect 50790 11350 50800 11410
rect 49030 11340 49110 11350
rect 52030 11330 55950 11340
rect 49970 11270 49980 11330
rect 50040 11320 50050 11330
rect 50040 11280 51980 11320
rect 50040 11270 50050 11280
rect 48920 11250 49000 11260
rect 48920 11190 48930 11250
rect 48990 11240 49000 11250
rect 48990 11230 51280 11240
rect 48990 11200 50070 11230
rect 48990 11190 49000 11200
rect 48920 11180 49000 11190
rect 50060 11170 50070 11200
rect 50130 11200 51280 11230
rect 51900 11220 51910 11280
rect 51970 11220 51980 11280
rect 52030 11270 52040 11330
rect 52100 11270 52240 11330
rect 52300 11270 53570 11330
rect 53630 11270 55950 11330
rect 52030 11260 55950 11270
rect 51900 11210 51980 11220
rect 50130 11170 50140 11200
rect 50060 11160 50140 11170
rect 50760 11160 50840 11170
rect 50760 11100 50770 11160
rect 50830 11100 50840 11160
rect 50760 11090 50840 11100
rect 51200 11160 51280 11200
rect 51200 11100 51210 11160
rect 51270 11100 51280 11160
rect 51200 11090 51280 11100
rect 52740 11160 53300 11170
rect 52740 11100 52750 11160
rect 52810 11100 53230 11160
rect 53290 11100 53300 11160
rect 52740 11090 53300 11100
rect 53540 11070 53650 11090
rect 53540 11000 53560 11070
rect 53630 11000 53650 11070
rect 53540 10980 53650 11000
rect 50980 10880 51060 10890
rect 50980 10820 50990 10880
rect 51050 10820 51060 10880
rect 50980 10810 51060 10820
rect 48790 10770 52200 10780
rect 48790 10710 49410 10770
rect 49470 10710 49610 10770
rect 49670 10710 49850 10770
rect 49910 10710 50010 10770
rect 50070 10710 50410 10770
rect 50470 10710 50810 10770
rect 50870 10710 51210 10770
rect 51270 10710 51410 10770
rect 51470 10710 52130 10770
rect 52190 10710 52200 10770
rect 48790 10700 52200 10710
rect 50980 10660 51060 10670
rect 50980 10600 50990 10660
rect 51050 10600 51060 10660
rect 50980 10590 51060 10600
rect 48790 9650 53090 9660
rect 48790 9590 53020 9650
rect 53080 9590 53090 9650
rect 48790 9580 53090 9590
rect 53210 9140 53310 9160
rect 53210 9080 53230 9140
rect 53290 9080 53310 9140
rect 53210 9060 53310 9080
<< via2 >>
rect 53230 13450 53290 13510
rect 53560 11510 53630 11580
rect 53560 11000 53630 11070
rect 53230 9080 53290 9140
<< metal3 >>
rect 53210 13520 53310 13530
rect 53210 13510 55950 13520
rect 53210 13450 53230 13510
rect 53290 13450 55950 13510
rect 53210 13430 55950 13450
rect 53540 11580 53650 11600
rect 53540 11510 53560 11580
rect 53630 11510 53650 11580
rect 53540 11490 53650 11510
rect 53890 11460 55950 13430
rect 53540 11070 53650 11090
rect 53540 11000 53560 11070
rect 53630 11000 53650 11070
rect 53540 10980 53650 11000
rect 53210 9150 53310 9160
rect 53890 9150 55950 11120
rect 53210 9140 55950 9150
rect 53210 9080 53230 9140
rect 53290 9080 55950 9140
rect 53210 9060 55950 9080
<< via3 >>
rect 53560 11510 53630 11580
rect 53560 11000 53630 11070
<< mimcap >>
rect 53920 11580 55920 13490
rect 53920 11510 53940 11580
rect 54010 11510 55920 11580
rect 53920 11490 55920 11510
rect 53920 11070 55920 11090
rect 53920 11000 53940 11070
rect 54010 11000 55920 11070
rect 53920 9090 55920 11000
<< mimcapcontact >>
rect 53940 11510 54010 11580
rect 53940 11000 54010 11070
<< metal4 >>
rect 53540 11580 54020 11600
rect 53540 11510 53560 11580
rect 53630 11510 53940 11580
rect 54010 11510 54020 11580
rect 53540 11490 54020 11510
rect 53540 11070 54020 11090
rect 53540 11000 53560 11070
rect 53630 11000 53940 11070
rect 54010 11000 54020 11070
rect 53540 10980 54020 11000
<< end >>
