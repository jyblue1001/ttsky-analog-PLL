magic
tech sky130A
magscale 1 2
timestamp 1757396817
<< locali >>
rect 15100 14690 15180 14710
rect 15100 14650 15120 14690
rect 15160 14650 15180 14690
rect 15100 14630 15180 14650
<< viali >>
rect 15120 14650 15160 14690
<< metal1 >>
rect 26000 19900 26480 19910
rect 26000 19840 26010 19900
rect 26070 19840 26100 19900
rect 26160 19840 26200 19900
rect 26260 19840 26310 19900
rect 26370 19840 26410 19900
rect 26470 19840 26480 19900
rect 15100 14700 15180 14710
rect 15100 14640 15110 14700
rect 15170 14640 15180 14700
rect 15100 14630 15180 14640
rect 15710 14700 15790 14710
rect 15710 14640 15720 14700
rect 15780 14640 15790 14700
rect 15710 14250 15790 14640
rect 15710 14190 15720 14250
rect 15780 14190 15790 14250
rect 15710 14170 15790 14190
rect 15710 14110 15720 14170
rect 15780 14110 15790 14170
rect 15710 14100 15790 14110
rect 18040 13420 18280 13440
rect 18040 13360 18080 13420
rect 18140 13360 18180 13420
rect 18240 13360 18280 13420
rect 18040 13340 18280 13360
rect 18650 9300 18890 9310
rect 18650 9240 18660 9300
rect 18720 9240 18740 9300
rect 18800 9240 18820 9300
rect 18880 9240 18890 9300
rect 18650 9220 18890 9240
rect 18650 9160 18660 9220
rect 18720 9160 18740 9220
rect 18800 9160 18820 9220
rect 18880 9160 18890 9220
rect 18650 9140 18890 9160
rect 18650 9080 18660 9140
rect 18720 9080 18740 9140
rect 18800 9080 18820 9140
rect 18880 9080 18890 9140
rect 12050 7810 12130 7820
rect 12050 7750 12060 7810
rect 12120 7750 12130 7810
rect 11940 6430 12020 6440
rect 11940 6370 11950 6430
rect 12010 6370 12020 6430
rect 11940 1330 12020 6370
rect 12050 3340 12130 7750
rect 18650 7380 18890 9080
rect 18650 7320 18660 7380
rect 18720 7320 18740 7380
rect 18800 7320 18820 7380
rect 18880 7320 18890 7380
rect 18650 7310 18890 7320
rect 18920 7040 19000 11580
rect 19030 8770 19110 11740
rect 19030 8710 19040 8770
rect 19100 8710 19110 8770
rect 19030 8690 19110 8710
rect 19030 8630 19040 8690
rect 19100 8630 19110 8690
rect 19030 8610 19110 8630
rect 19030 8550 19040 8610
rect 19100 8550 19110 8610
rect 19030 8540 19110 8550
rect 26000 8770 26480 19840
rect 26000 8710 26010 8770
rect 26070 8710 26090 8770
rect 26150 8710 26170 8770
rect 26230 8710 26250 8770
rect 26310 8710 26330 8770
rect 26390 8710 26410 8770
rect 26470 8710 26480 8770
rect 26000 8690 26480 8710
rect 26000 8630 26010 8690
rect 26070 8630 26090 8690
rect 26150 8630 26170 8690
rect 26230 8630 26250 8690
rect 26310 8630 26330 8690
rect 26390 8630 26410 8690
rect 26470 8630 26480 8690
rect 26000 8610 26480 8630
rect 26000 8550 26010 8610
rect 26070 8550 26090 8610
rect 26150 8550 26170 8610
rect 26230 8550 26250 8610
rect 26310 8550 26330 8610
rect 26390 8550 26410 8610
rect 26470 8550 26480 8610
rect 19140 8500 19220 8510
rect 19140 8440 19150 8500
rect 19210 8440 19220 8500
rect 19140 7160 19220 8440
rect 19140 7100 19150 7160
rect 19210 7100 19220 7160
rect 19140 7090 19220 7100
rect 26000 7320 26480 8550
rect 26510 11730 26590 11740
rect 26510 11670 26520 11730
rect 26580 11670 26590 11730
rect 26510 8500 26590 11670
rect 26510 8440 26520 8500
rect 26580 8440 26590 8500
rect 26510 8430 26590 8440
rect 26000 7260 26010 7320
rect 26070 7260 26090 7320
rect 26150 7260 26170 7320
rect 26230 7260 26250 7320
rect 26310 7260 26330 7320
rect 26390 7260 26410 7320
rect 26470 7260 26480 7320
rect 18920 6980 18930 7040
rect 18990 6980 19000 7040
rect 18920 6970 19000 6980
rect 12050 3280 12060 3340
rect 12120 3280 12130 3340
rect 12050 3270 12130 3280
rect 26000 2280 26480 7260
rect 26000 2220 26010 2280
rect 26070 2220 26090 2280
rect 26150 2220 26170 2280
rect 26230 2220 26250 2280
rect 26310 2220 26330 2280
rect 26390 2220 26410 2280
rect 26470 2220 26480 2280
rect 26000 2210 26480 2220
rect 11940 1270 11950 1330
rect 12010 1270 12020 1330
rect 11940 1260 12020 1270
<< via1 >>
rect 26010 19840 26070 19900
rect 26100 19840 26160 19900
rect 26200 19840 26260 19900
rect 26310 19840 26370 19900
rect 26410 19840 26470 19900
rect 15110 14690 15170 14700
rect 15110 14650 15120 14690
rect 15120 14650 15160 14690
rect 15160 14650 15170 14690
rect 15110 14640 15170 14650
rect 15720 14640 15780 14700
rect 15720 14190 15780 14250
rect 15720 14110 15780 14170
rect 18080 13360 18140 13420
rect 18180 13360 18240 13420
rect 18660 9240 18720 9300
rect 18740 9240 18800 9300
rect 18820 9240 18880 9300
rect 18660 9160 18720 9220
rect 18740 9160 18800 9220
rect 18820 9160 18880 9220
rect 18660 9080 18720 9140
rect 18740 9080 18800 9140
rect 18820 9080 18880 9140
rect 12060 7750 12120 7810
rect 11950 6370 12010 6430
rect 18660 7320 18720 7380
rect 18740 7320 18800 7380
rect 18820 7320 18880 7380
rect 19040 8710 19100 8770
rect 19040 8630 19100 8690
rect 19040 8550 19100 8610
rect 26010 8710 26070 8770
rect 26090 8710 26150 8770
rect 26170 8710 26230 8770
rect 26250 8710 26310 8770
rect 26330 8710 26390 8770
rect 26410 8710 26470 8770
rect 26010 8630 26070 8690
rect 26090 8630 26150 8690
rect 26170 8630 26230 8690
rect 26250 8630 26310 8690
rect 26330 8630 26390 8690
rect 26410 8630 26470 8690
rect 26010 8550 26070 8610
rect 26090 8550 26150 8610
rect 26170 8550 26230 8610
rect 26250 8550 26310 8610
rect 26330 8550 26390 8610
rect 26410 8550 26470 8610
rect 19150 8440 19210 8500
rect 19150 7100 19210 7160
rect 26520 11670 26580 11730
rect 26520 8440 26580 8500
rect 26010 7260 26070 7320
rect 26090 7260 26150 7320
rect 26170 7260 26230 7320
rect 26250 7260 26310 7320
rect 26330 7260 26390 7320
rect 26410 7260 26470 7320
rect 18930 6980 18990 7040
rect 12060 3280 12120 3340
rect 26010 2220 26070 2280
rect 26090 2220 26150 2280
rect 26170 2220 26230 2280
rect 26250 2220 26310 2280
rect 26330 2220 26390 2280
rect 26410 2220 26470 2280
rect 11950 1270 12010 1330
<< metal2 >>
rect 7460 20280 7720 20290
rect 7460 20220 7470 20280
rect 7530 20220 7560 20280
rect 7620 20220 7650 20280
rect 7710 20220 7720 20280
rect 7460 20190 7720 20220
rect 7460 20130 7470 20190
rect 7530 20130 7560 20190
rect 7620 20130 7650 20190
rect 7710 20130 7720 20190
rect 7460 20100 7720 20130
rect 7460 20040 7470 20100
rect 7530 20040 7560 20100
rect 7620 20040 7650 20100
rect 7710 20040 7720 20100
rect 7460 20030 7720 20040
rect 26000 19900 26480 19920
rect 26000 19840 26010 19900
rect 26070 19840 26100 19900
rect 26160 19840 26200 19900
rect 26260 19840 26310 19900
rect 26370 19840 26410 19900
rect 26470 19840 26480 19900
rect 26000 19820 26480 19840
rect 18020 19520 18100 19600
rect 7460 19450 8790 19490
rect 7460 19390 7470 19450
rect 7530 19390 7560 19450
rect 7620 19390 7650 19450
rect 7710 19390 8790 19450
rect 7460 19350 8790 19390
rect 7460 19290 7470 19350
rect 7530 19290 7560 19350
rect 7620 19290 7650 19350
rect 7710 19290 8790 19350
rect 7460 19250 8790 19290
rect 18360 16380 18440 16460
rect 11220 14740 11300 14820
rect 15100 14700 15790 14710
rect 15100 14640 15110 14700
rect 15170 14640 15720 14700
rect 15780 14640 15790 14700
rect 15100 14630 15790 14640
rect 15550 14250 18580 14260
rect 15550 14190 15720 14250
rect 15780 14210 18580 14250
rect 15780 14190 18380 14210
rect 15550 14170 18380 14190
rect 15550 14110 15720 14170
rect 15780 14150 18380 14170
rect 18440 14150 18480 14210
rect 18540 14150 18580 14210
rect 15780 14110 18580 14150
rect 15550 14100 18580 14110
rect 14660 13900 18580 13940
rect 14660 13840 18380 13900
rect 18440 13840 18480 13900
rect 18540 13840 18580 13900
rect 14660 13800 18580 13840
rect 14660 13740 18380 13800
rect 18440 13740 18480 13800
rect 18540 13740 18580 13800
rect 14660 13700 18580 13740
rect 18340 13580 18790 13590
rect 18340 13520 18380 13580
rect 18440 13520 18480 13580
rect 18540 13520 18790 13580
rect 18340 13510 18790 13520
rect 18040 13420 18280 13440
rect 18040 13360 18080 13420
rect 18140 13360 18180 13420
rect 18240 13360 18280 13420
rect 18040 13340 18280 13360
rect 15640 13100 18280 13140
rect 15640 13040 18080 13100
rect 18140 13040 18180 13100
rect 18240 13040 18280 13100
rect 15640 13000 18280 13040
rect 15640 12940 18080 13000
rect 18140 12940 18180 13000
rect 18240 12940 18280 13000
rect 15640 12900 18280 12940
rect 18040 12400 18280 12410
rect 18040 12390 18790 12400
rect 18040 12330 18080 12390
rect 18140 12330 18180 12390
rect 18240 12330 18790 12390
rect 18040 12320 18790 12330
rect 18040 12310 18280 12320
rect 25950 11730 26590 11740
rect 25950 11670 26520 11730
rect 26580 11670 26590 11730
rect 25950 11660 26590 11670
rect 16040 11440 18280 11480
rect 16040 11380 18080 11440
rect 18140 11380 18180 11440
rect 18240 11380 18280 11440
rect 16040 11340 18280 11380
rect 16040 11280 18080 11340
rect 18140 11280 18180 11340
rect 18240 11280 18280 11340
rect 16040 11240 18280 11280
rect 10090 11140 10160 11210
rect 18340 11180 18580 11190
rect 18340 11170 18790 11180
rect 18340 11110 18380 11170
rect 18440 11110 18480 11170
rect 18540 11110 18790 11170
rect 18340 11100 18790 11110
rect 18340 11090 18580 11100
rect 12000 10730 12040 10770
rect 18340 10050 18790 10060
rect 16010 9990 18280 10030
rect 16010 9930 18080 9990
rect 18140 9930 18180 9990
rect 18240 9930 18280 9990
rect 18340 9990 18380 10050
rect 18440 9990 18480 10050
rect 18540 9990 18790 10050
rect 18340 9980 18790 9990
rect 16010 9890 18280 9930
rect 16010 9830 18080 9890
rect 18140 9830 18180 9890
rect 18240 9830 18280 9890
rect 16010 9790 18280 9830
rect 18040 9430 18280 9440
rect 14930 9420 18280 9430
rect 14930 9360 18080 9420
rect 18140 9360 18180 9420
rect 18240 9360 18280 9420
rect 14930 9350 18280 9360
rect 18040 9340 18280 9350
rect 10160 9240 10240 9320
rect 14820 9300 18890 9310
rect 14820 9240 18660 9300
rect 18720 9240 18740 9300
rect 18800 9240 18820 9300
rect 18880 9240 18890 9300
rect 14820 9220 18890 9240
rect 14820 9160 18660 9220
rect 18720 9160 18740 9220
rect 18800 9160 18820 9220
rect 18880 9160 18890 9220
rect 14820 9140 18890 9160
rect 14820 9080 18660 9140
rect 18720 9080 18740 9140
rect 18800 9080 18820 9140
rect 18880 9080 18890 9140
rect 14820 9070 18890 9080
rect 19030 8770 26480 8780
rect 19030 8710 19040 8770
rect 19100 8710 26010 8770
rect 26070 8710 26090 8770
rect 26150 8710 26170 8770
rect 26230 8710 26250 8770
rect 26310 8710 26330 8770
rect 26390 8710 26410 8770
rect 26470 8710 26480 8770
rect 19030 8690 26480 8710
rect 19030 8630 19040 8690
rect 19100 8630 26010 8690
rect 26070 8630 26090 8690
rect 26150 8630 26170 8690
rect 26230 8630 26250 8690
rect 26310 8630 26330 8690
rect 26390 8630 26410 8690
rect 26470 8630 26480 8690
rect 19030 8610 26480 8630
rect 19030 8550 19040 8610
rect 19100 8550 26010 8610
rect 26070 8550 26090 8610
rect 26150 8550 26170 8610
rect 26230 8550 26250 8610
rect 26310 8550 26330 8610
rect 26390 8550 26410 8610
rect 26470 8550 26480 8610
rect 19030 8540 26480 8550
rect 19140 8500 26590 8510
rect 19140 8440 19150 8500
rect 19210 8440 26520 8500
rect 26580 8440 26590 8500
rect 19140 8430 26590 8440
rect 12910 8350 13010 8390
rect 12910 8290 12930 8350
rect 12990 8290 13010 8350
rect 12910 8250 13010 8290
rect 12910 8190 12930 8250
rect 12990 8190 13010 8250
rect 12910 8150 13010 8190
rect 18340 8230 19340 8240
rect 18340 8170 18380 8230
rect 18440 8170 18480 8230
rect 18540 8170 19340 8230
rect 18340 8160 19340 8170
rect 12050 7810 13010 7820
rect 12050 7750 12060 7810
rect 12120 7750 13010 7810
rect 12050 7740 13010 7750
rect 18650 7380 18890 7390
rect 18650 7320 18660 7380
rect 18720 7320 18740 7380
rect 18800 7320 18820 7380
rect 18880 7320 18890 7380
rect 18650 7310 18890 7320
rect 24190 7320 26480 7330
rect 24190 7260 26010 7320
rect 26070 7260 26090 7320
rect 26150 7260 26170 7320
rect 26230 7260 26250 7320
rect 26310 7260 26330 7320
rect 26390 7260 26410 7320
rect 26470 7260 26480 7320
rect 24190 7250 26480 7260
rect 12910 7170 13010 7210
rect 12910 7110 12930 7170
rect 12990 7110 13010 7170
rect 12910 7070 13010 7110
rect 19140 7160 19220 7170
rect 19140 7100 19150 7160
rect 19210 7100 19220 7160
rect 19140 7090 19220 7100
rect 12910 7010 12930 7070
rect 12990 7010 13010 7070
rect 12910 6970 13010 7010
rect 18920 7040 19980 7050
rect 18920 6980 18930 7040
rect 18990 6980 19980 7040
rect 18920 6970 19980 6980
rect 11940 6430 13010 6440
rect 11940 6370 11950 6430
rect 12010 6370 13010 6430
rect 11940 6360 13010 6370
rect 19240 6390 19540 6400
rect 19240 6330 19280 6390
rect 19340 6330 19380 6390
rect 19440 6330 19540 6390
rect 19240 6320 19540 6330
rect 12910 5990 13010 6030
rect 12910 5930 12930 5990
rect 12990 5930 13010 5990
rect 12910 5890 13010 5930
rect 12910 5830 12930 5890
rect 12990 5830 13010 5890
rect 12910 5790 13010 5830
rect 22590 5690 22690 5730
rect 22590 5630 22610 5690
rect 22670 5650 22690 5690
rect 22670 5630 23580 5650
rect 22590 5590 23580 5630
rect 22590 5530 22610 5590
rect 22670 5570 23580 5590
rect 22670 5530 22690 5570
rect 22590 5490 22690 5530
rect 12160 3790 12260 3830
rect 12160 3730 12180 3790
rect 12240 3730 12260 3790
rect 12160 3690 12260 3730
rect 12160 3630 12180 3690
rect 12240 3630 12260 3690
rect 12160 3590 12260 3630
rect 25410 3400 26670 3420
rect 12050 3340 12130 3350
rect 12050 3280 12060 3340
rect 12120 3280 12130 3340
rect 12050 3270 12130 3280
rect 25410 3320 26550 3400
rect 26630 3320 26670 3400
rect 25410 3280 26670 3320
rect 25410 3200 26550 3280
rect 26630 3200 26670 3280
rect 25410 3180 26670 3200
rect 12160 3010 12260 3050
rect 12160 2950 12180 3010
rect 12240 2950 12260 3010
rect 12160 2910 12260 2950
rect 12160 2850 12180 2910
rect 12240 2850 12260 2910
rect 12160 2810 12260 2850
rect 24950 2220 26010 2280
rect 26070 2220 26090 2280
rect 26150 2220 26170 2280
rect 26230 2220 26250 2280
rect 26310 2220 26330 2280
rect 26390 2220 26410 2280
rect 26470 2220 26480 2280
rect 24950 2210 26480 2220
rect 22590 1610 22690 1650
rect 22590 1550 22610 1610
rect 22670 1570 22690 1610
rect 22670 1550 23310 1570
rect 22590 1510 23310 1550
rect 22590 1450 22610 1510
rect 22670 1490 23310 1510
rect 22670 1450 22690 1490
rect 22590 1410 22690 1450
rect 30370 1340 30530 1380
rect 11940 1330 30410 1340
rect 11940 1270 11950 1330
rect 12010 1270 30410 1330
rect 11940 1260 30410 1270
rect 30490 1260 30530 1340
rect 30370 1220 30530 1260
<< via2 >>
rect 7470 20220 7530 20280
rect 7560 20220 7620 20280
rect 7650 20220 7710 20280
rect 7470 20130 7530 20190
rect 7560 20130 7620 20190
rect 7650 20130 7710 20190
rect 7470 20040 7530 20100
rect 7560 20040 7620 20100
rect 7650 20040 7710 20100
rect 7470 19390 7530 19450
rect 7560 19390 7620 19450
rect 7650 19390 7710 19450
rect 7470 19290 7530 19350
rect 7560 19290 7620 19350
rect 7650 19290 7710 19350
rect 18380 14150 18440 14210
rect 18480 14150 18540 14210
rect 18380 13840 18440 13900
rect 18480 13840 18540 13900
rect 18380 13740 18440 13800
rect 18480 13740 18540 13800
rect 18380 13520 18440 13580
rect 18480 13520 18540 13580
rect 18080 13360 18140 13420
rect 18180 13360 18240 13420
rect 18080 13040 18140 13100
rect 18180 13040 18240 13100
rect 18080 12940 18140 13000
rect 18180 12940 18240 13000
rect 18080 12330 18140 12390
rect 18180 12330 18240 12390
rect 18080 11380 18140 11440
rect 18180 11380 18240 11440
rect 18080 11280 18140 11340
rect 18180 11280 18240 11340
rect 18380 11110 18440 11170
rect 18480 11110 18540 11170
rect 18080 9930 18140 9990
rect 18180 9930 18240 9990
rect 18380 9990 18440 10050
rect 18480 9990 18540 10050
rect 18080 9830 18140 9890
rect 18180 9830 18240 9890
rect 18080 9360 18140 9420
rect 18180 9360 18240 9420
rect 12930 8290 12990 8350
rect 12930 8190 12990 8250
rect 18380 8170 18440 8230
rect 18480 8170 18540 8230
rect 12930 7110 12990 7170
rect 12930 7010 12990 7070
rect 19280 6330 19340 6390
rect 19380 6330 19440 6390
rect 12930 5930 12990 5990
rect 12930 5830 12990 5890
rect 22610 5630 22670 5690
rect 22610 5530 22670 5590
rect 12180 3730 12240 3790
rect 12180 3630 12240 3690
rect 26550 3320 26630 3400
rect 26550 3200 26630 3280
rect 12180 2950 12240 3010
rect 12180 2850 12240 2910
rect 22610 1550 22670 1610
rect 22610 1450 22670 1510
rect 30410 1260 30490 1340
<< metal3 >>
rect 800 20280 7720 20290
rect 800 20250 7470 20280
rect 800 20170 810 20250
rect 890 20170 910 20250
rect 990 20170 1010 20250
rect 1090 20170 1110 20250
rect 1190 20220 7470 20250
rect 7530 20220 7560 20280
rect 7620 20220 7650 20280
rect 7710 20220 7720 20280
rect 1190 20190 7720 20220
rect 1190 20170 7470 20190
rect 800 20150 7470 20170
rect 800 20070 810 20150
rect 890 20070 910 20150
rect 990 20070 1010 20150
rect 1090 20070 1110 20150
rect 1190 20130 7470 20150
rect 7530 20130 7560 20190
rect 7620 20130 7650 20190
rect 7710 20130 7720 20190
rect 1190 20100 7720 20130
rect 1190 20070 7470 20100
rect 800 20040 7470 20070
rect 7530 20040 7560 20100
rect 7620 20040 7650 20100
rect 7710 20040 7720 20100
rect 800 20030 7720 20040
rect 800 19460 7720 19490
rect 800 19380 810 19460
rect 890 19380 910 19460
rect 990 19380 1010 19460
rect 1090 19380 1110 19460
rect 1190 19450 7720 19460
rect 1190 19390 7470 19450
rect 7530 19390 7560 19450
rect 7620 19390 7650 19450
rect 7710 19390 7720 19450
rect 1190 19380 7720 19390
rect 800 19360 7720 19380
rect 800 19280 810 19360
rect 890 19280 910 19360
rect 990 19280 1010 19360
rect 1090 19280 1110 19360
rect 1190 19350 7720 19360
rect 1190 19290 7470 19350
rect 7530 19290 7560 19350
rect 7620 19290 7650 19350
rect 7710 19290 7720 19350
rect 1190 19280 7720 19290
rect 800 19250 7720 19280
rect 18340 14210 18580 14260
rect 18340 14150 18380 14210
rect 18440 14150 18480 14210
rect 18540 14150 18580 14210
rect 18340 13900 18580 14150
rect 18340 13840 18380 13900
rect 18440 13840 18480 13900
rect 18540 13840 18580 13900
rect 18340 13800 18580 13840
rect 23680 13830 23770 13920
rect 18340 13740 18380 13800
rect 18440 13740 18480 13800
rect 18540 13740 18580 13800
rect 18340 13580 18580 13740
rect 18340 13520 18380 13580
rect 18440 13520 18480 13580
rect 18540 13520 18580 13580
rect 18040 13420 18280 13440
rect 18040 13360 18080 13420
rect 18140 13360 18180 13420
rect 18240 13360 18280 13420
rect 18040 13100 18280 13360
rect 18040 13040 18080 13100
rect 18140 13040 18180 13100
rect 18240 13040 18280 13100
rect 18040 13000 18280 13040
rect 18040 12940 18080 13000
rect 18140 12940 18180 13000
rect 18240 12940 18280 13000
rect 18040 12390 18280 12940
rect 18040 12330 18080 12390
rect 18140 12330 18180 12390
rect 18240 12330 18280 12390
rect 18040 11440 18280 12330
rect 18040 11380 18080 11440
rect 18140 11380 18180 11440
rect 18240 11380 18280 11440
rect 18040 11340 18280 11380
rect 18040 11280 18080 11340
rect 18140 11280 18180 11340
rect 18240 11280 18280 11340
rect 18040 9990 18280 11280
rect 18040 9930 18080 9990
rect 18140 9930 18180 9990
rect 18240 9930 18280 9990
rect 18040 9890 18280 9930
rect 18040 9830 18080 9890
rect 18140 9830 18180 9890
rect 18240 9830 18280 9890
rect 18040 9420 18280 9830
rect 18040 9360 18080 9420
rect 18140 9360 18180 9420
rect 18240 9360 18280 9420
rect 18040 9040 18280 9360
rect 200 9010 18280 9040
rect 200 8930 210 9010
rect 290 8930 310 9010
rect 390 8930 410 9010
rect 490 8930 510 9010
rect 590 8930 18280 9010
rect 200 8910 18280 8930
rect 200 8830 210 8910
rect 290 8830 310 8910
rect 390 8830 410 8910
rect 490 8830 510 8910
rect 590 8830 18280 8910
rect 200 8800 18280 8830
rect 18340 11170 18580 13520
rect 18340 11110 18380 11170
rect 18440 11110 18480 11170
rect 18540 11110 18580 11170
rect 18340 10050 18580 11110
rect 18340 9990 18380 10050
rect 18440 9990 18480 10050
rect 18540 9990 18580 10050
rect 18340 8740 18580 9990
rect 23670 9460 23760 9550
rect 800 8710 18580 8740
rect 800 8630 810 8710
rect 890 8630 910 8710
rect 990 8630 1010 8710
rect 1090 8630 1110 8710
rect 1190 8630 18580 8710
rect 800 8610 18580 8630
rect 800 8530 810 8610
rect 890 8530 910 8610
rect 990 8530 1010 8610
rect 1090 8530 1110 8610
rect 1190 8530 18580 8610
rect 800 8500 18580 8530
rect 800 8360 13010 8390
rect 800 8280 810 8360
rect 890 8280 910 8360
rect 990 8280 1010 8360
rect 1090 8280 1110 8360
rect 1190 8350 13010 8360
rect 1190 8290 12930 8350
rect 12990 8290 13010 8350
rect 1190 8280 13010 8290
rect 800 8260 13010 8280
rect 800 8180 810 8260
rect 890 8180 910 8260
rect 990 8180 1010 8260
rect 1090 8180 1110 8260
rect 1190 8250 13010 8260
rect 1190 8190 12930 8250
rect 12990 8190 13010 8250
rect 1190 8180 13010 8190
rect 800 8150 13010 8180
rect 18340 8230 18580 8500
rect 18340 8170 18380 8230
rect 18440 8170 18480 8230
rect 18540 8170 18580 8230
rect 18340 8160 18580 8170
rect 200 7180 13010 7210
rect 200 7100 210 7180
rect 290 7100 310 7180
rect 390 7100 410 7180
rect 490 7100 510 7180
rect 590 7170 13010 7180
rect 590 7110 12930 7170
rect 12990 7110 13010 7170
rect 590 7100 13010 7110
rect 200 7080 13010 7100
rect 200 7000 210 7080
rect 290 7000 310 7080
rect 390 7000 410 7080
rect 490 7000 510 7080
rect 590 7070 13010 7080
rect 590 7010 12930 7070
rect 12990 7010 13010 7070
rect 590 7000 13010 7010
rect 200 6970 13010 7000
rect 19240 6390 19480 6400
rect 19240 6330 19280 6390
rect 19340 6330 19380 6390
rect 19440 6330 19480 6390
rect 800 6000 13010 6030
rect 800 5920 810 6000
rect 890 5920 910 6000
rect 990 5920 1010 6000
rect 1090 5920 1110 6000
rect 1190 5990 13010 6000
rect 1190 5930 12930 5990
rect 12990 5930 13010 5990
rect 1190 5920 13010 5930
rect 800 5900 13010 5920
rect 800 5820 810 5900
rect 890 5820 910 5900
rect 990 5820 1010 5900
rect 1090 5820 1110 5900
rect 1190 5890 13010 5900
rect 1190 5830 12930 5890
rect 12990 5830 13010 5890
rect 1190 5820 13010 5830
rect 800 5790 13010 5820
rect 19240 5730 19480 6330
rect 200 5700 22690 5730
rect 200 5620 210 5700
rect 290 5620 310 5700
rect 390 5620 410 5700
rect 490 5620 510 5700
rect 590 5690 22690 5700
rect 590 5630 22610 5690
rect 22670 5630 22690 5690
rect 590 5620 22690 5630
rect 200 5600 22690 5620
rect 200 5520 210 5600
rect 290 5520 310 5600
rect 390 5520 410 5600
rect 490 5520 510 5600
rect 590 5590 22690 5600
rect 590 5530 22610 5590
rect 22670 5530 22690 5590
rect 590 5520 22690 5530
rect 200 5490 22690 5520
rect 200 3800 12260 3830
rect 200 3720 210 3800
rect 290 3720 310 3800
rect 390 3720 410 3800
rect 490 3720 510 3800
rect 590 3790 12260 3800
rect 590 3730 12180 3790
rect 12240 3730 12260 3790
rect 590 3720 12260 3730
rect 200 3700 12260 3720
rect 200 3620 210 3700
rect 290 3620 310 3700
rect 390 3620 410 3700
rect 490 3620 510 3700
rect 590 3690 12260 3700
rect 590 3630 12180 3690
rect 12240 3630 12260 3690
rect 590 3620 12260 3630
rect 200 3590 12260 3620
rect 26510 3400 26670 3420
rect 26510 3320 26550 3400
rect 26630 3320 26670 3400
rect 26510 3280 26670 3320
rect 26510 3200 26550 3280
rect 26630 3200 26670 3280
rect 26510 3180 26670 3200
rect 800 3020 12260 3050
rect 800 2940 810 3020
rect 890 2940 910 3020
rect 990 2940 1010 3020
rect 1090 2940 1110 3020
rect 1190 3010 12260 3020
rect 1190 2950 12180 3010
rect 12240 2950 12260 3010
rect 1190 2940 12260 2950
rect 800 2920 12260 2940
rect 800 2840 810 2920
rect 890 2840 910 2920
rect 990 2840 1010 2920
rect 1090 2840 1110 2920
rect 1190 2910 12260 2920
rect 1190 2850 12180 2910
rect 12240 2850 12260 2910
rect 1190 2840 12260 2850
rect 800 2810 12260 2840
rect 800 1620 22690 1650
rect 800 1540 810 1620
rect 890 1540 910 1620
rect 990 1540 1010 1620
rect 1090 1540 1110 1620
rect 1190 1610 22690 1620
rect 1190 1550 22610 1610
rect 22670 1550 22690 1610
rect 1190 1540 22690 1550
rect 800 1520 22690 1540
rect 800 1440 810 1520
rect 890 1440 910 1520
rect 990 1440 1010 1520
rect 1090 1440 1110 1520
rect 1190 1510 22690 1520
rect 1190 1450 22610 1510
rect 22670 1450 22690 1510
rect 1190 1440 22690 1450
rect 800 1410 22690 1440
rect 30370 1340 30530 1380
rect 30370 1260 30410 1340
rect 30490 1260 30530 1340
rect 30370 1220 30530 1260
<< via3 >>
rect 810 20170 890 20250
rect 910 20170 990 20250
rect 1010 20170 1090 20250
rect 1110 20170 1190 20250
rect 810 20070 890 20150
rect 910 20070 990 20150
rect 1010 20070 1090 20150
rect 1110 20070 1190 20150
rect 810 19380 890 19460
rect 910 19380 990 19460
rect 1010 19380 1090 19460
rect 1110 19380 1190 19460
rect 810 19280 890 19360
rect 910 19280 990 19360
rect 1010 19280 1090 19360
rect 1110 19280 1190 19360
rect 210 8930 290 9010
rect 310 8930 390 9010
rect 410 8930 490 9010
rect 510 8930 590 9010
rect 210 8830 290 8910
rect 310 8830 390 8910
rect 410 8830 490 8910
rect 510 8830 590 8910
rect 810 8630 890 8710
rect 910 8630 990 8710
rect 1010 8630 1090 8710
rect 1110 8630 1190 8710
rect 810 8530 890 8610
rect 910 8530 990 8610
rect 1010 8530 1090 8610
rect 1110 8530 1190 8610
rect 810 8280 890 8360
rect 910 8280 990 8360
rect 1010 8280 1090 8360
rect 1110 8280 1190 8360
rect 810 8180 890 8260
rect 910 8180 990 8260
rect 1010 8180 1090 8260
rect 1110 8180 1190 8260
rect 210 7100 290 7180
rect 310 7100 390 7180
rect 410 7100 490 7180
rect 510 7100 590 7180
rect 210 7000 290 7080
rect 310 7000 390 7080
rect 410 7000 490 7080
rect 510 7000 590 7080
rect 810 5920 890 6000
rect 910 5920 990 6000
rect 1010 5920 1090 6000
rect 1110 5920 1190 6000
rect 810 5820 890 5900
rect 910 5820 990 5900
rect 1010 5820 1090 5900
rect 1110 5820 1190 5900
rect 210 5620 290 5700
rect 310 5620 390 5700
rect 410 5620 490 5700
rect 510 5620 590 5700
rect 210 5520 290 5600
rect 310 5520 390 5600
rect 410 5520 490 5600
rect 510 5520 590 5600
rect 210 3720 290 3800
rect 310 3720 390 3800
rect 410 3720 490 3800
rect 510 3720 590 3800
rect 210 3620 290 3700
rect 310 3620 390 3700
rect 410 3620 490 3700
rect 510 3620 590 3700
rect 26550 3320 26630 3400
rect 26550 3200 26630 3280
rect 810 2940 890 3020
rect 910 2940 990 3020
rect 1010 2940 1090 3020
rect 1110 2940 1190 3020
rect 810 2840 890 2920
rect 910 2840 990 2920
rect 1010 2840 1090 2920
rect 1110 2840 1190 2920
rect 810 1540 890 1620
rect 910 1540 990 1620
rect 1010 1540 1090 1620
rect 1110 1540 1190 1620
rect 810 1440 890 1520
rect 910 1440 990 1520
rect 1010 1440 1090 1520
rect 1110 1440 1190 1520
rect 30410 1260 30490 1340
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 9010 600 44152
rect 200 8930 210 9010
rect 290 8930 310 9010
rect 390 8930 410 9010
rect 490 8930 510 9010
rect 590 8930 600 9010
rect 200 8910 600 8930
rect 200 8830 210 8910
rect 290 8830 310 8910
rect 390 8830 410 8910
rect 490 8830 510 8910
rect 590 8830 600 8910
rect 200 7180 600 8830
rect 200 7100 210 7180
rect 290 7100 310 7180
rect 390 7100 410 7180
rect 490 7100 510 7180
rect 590 7100 600 7180
rect 200 7080 600 7100
rect 200 7000 210 7080
rect 290 7000 310 7080
rect 390 7000 410 7080
rect 490 7000 510 7080
rect 590 7000 600 7080
rect 200 5700 600 7000
rect 200 5620 210 5700
rect 290 5620 310 5700
rect 390 5620 410 5700
rect 490 5620 510 5700
rect 590 5620 600 5700
rect 200 5600 600 5620
rect 200 5520 210 5600
rect 290 5520 310 5600
rect 390 5520 410 5600
rect 490 5520 510 5600
rect 590 5520 600 5600
rect 200 3800 600 5520
rect 200 3720 210 3800
rect 290 3720 310 3800
rect 390 3720 410 3800
rect 490 3720 510 3800
rect 590 3720 600 3800
rect 200 3700 600 3720
rect 200 3620 210 3700
rect 290 3620 310 3700
rect 390 3620 410 3700
rect 490 3620 510 3700
rect 590 3620 600 3700
rect 200 1000 600 3620
rect 800 20250 1200 44152
rect 800 20170 810 20250
rect 890 20170 910 20250
rect 990 20170 1010 20250
rect 1090 20170 1110 20250
rect 1190 20170 1200 20250
rect 800 20150 1200 20170
rect 800 20070 810 20150
rect 890 20070 910 20150
rect 990 20070 1010 20150
rect 1090 20070 1110 20150
rect 1190 20070 1200 20150
rect 800 19460 1200 20070
rect 800 19380 810 19460
rect 890 19380 910 19460
rect 990 19380 1010 19460
rect 1090 19380 1110 19460
rect 1190 19380 1200 19460
rect 800 19360 1200 19380
rect 800 19280 810 19360
rect 890 19280 910 19360
rect 990 19280 1010 19360
rect 1090 19280 1110 19360
rect 1190 19280 1200 19360
rect 800 8710 1200 19280
rect 800 8630 810 8710
rect 890 8630 910 8710
rect 990 8630 1010 8710
rect 1090 8630 1110 8710
rect 1190 8630 1200 8710
rect 800 8610 1200 8630
rect 800 8530 810 8610
rect 890 8530 910 8610
rect 990 8530 1010 8610
rect 1090 8530 1110 8610
rect 1190 8530 1200 8610
rect 800 8360 1200 8530
rect 800 8280 810 8360
rect 890 8280 910 8360
rect 990 8280 1010 8360
rect 1090 8280 1110 8360
rect 1190 8280 1200 8360
rect 800 8260 1200 8280
rect 800 8180 810 8260
rect 890 8180 910 8260
rect 990 8180 1010 8260
rect 1090 8180 1110 8260
rect 1190 8180 1200 8260
rect 800 6000 1200 8180
rect 800 5920 810 6000
rect 890 5920 910 6000
rect 990 5920 1010 6000
rect 1090 5920 1110 6000
rect 1190 5920 1200 6000
rect 800 5900 1200 5920
rect 800 5820 810 5900
rect 890 5820 910 5900
rect 990 5820 1010 5900
rect 1090 5820 1110 5900
rect 1190 5820 1200 5900
rect 800 3020 1200 5820
rect 800 2940 810 3020
rect 890 2940 910 3020
rect 990 2940 1010 3020
rect 1090 2940 1110 3020
rect 1190 2940 1200 3020
rect 800 2920 1200 2940
rect 800 2840 810 2920
rect 890 2840 910 2920
rect 990 2840 1010 2920
rect 1090 2840 1110 2920
rect 1190 2840 1200 2920
rect 800 1620 1200 2840
rect 800 1540 810 1620
rect 890 1540 910 1620
rect 990 1540 1010 1620
rect 1090 1540 1110 1620
rect 1190 1540 1200 1620
rect 800 1520 1200 1540
rect 800 1440 810 1520
rect 890 1440 910 1520
rect 990 1440 1010 1520
rect 1090 1440 1110 1520
rect 1190 1440 1200 1520
rect 800 1000 1200 1440
rect 26510 3400 26670 3420
rect 26510 3320 26550 3400
rect 26630 3320 26670 3400
rect 26510 3280 26670 3320
rect 26510 3200 26550 3280
rect 26630 3200 26670 3280
rect 26510 200 26670 3200
rect 30370 1340 30530 1380
rect 30370 1260 30410 1340
rect 30490 1260 30530 1340
rect 30370 200 30530 1260
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use bgr  bgr_0
timestamp 1757393620
transform 1 0 -30000 0 1 400
box 38567 8670 55880 19200
use cp_opamp  cp_opamp_0
timestamp 1757393692
transform 1 0 -30000 0 1 400
box 48790 9060 55950 13791
use divide_by_120  divide_by_120_0
timestamp 1757393171
transform 1 0 -30000 0 1 0
box 42130 2890 52810 3750
use loop_filter  loop_filter_0
timestamp 1757393363
transform 1 0 -40000 0 1 400
box 47720 19209 66090 32110
use pfd_cp  pfd_cp_0
timestamp 1757393487
transform 1 0 -30000 0 1 0
box 43010 5790 54190 8400
use vco  vco_0
timestamp 1757392821
transform 1 0 -20000 0 1 0
box 42810 1490 45410 5650
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal1 18650 7760 18650 7760 7 FreeSans 1600 0 -800 0 I_IN
flabel metal2 18400 16380 18400 16380 5 FreeSans 1600 0 0 -800 cap_res1
flabel metal2 18060 19520 18060 19520 5 FreeSans 1600 0 0 -800 cap_res2
flabel metal2 11260 14740 11260 14740 5 FreeSans 1600 0 0 -800 Vbe2
flabel metal1 26080 2390 26080 2390 3 FreeSans 1600 0 800 0 V_CONT
flabel metal3 23730 13920 23730 13920 1 FreeSans 1600 0 0 800 res1
flabel metal3 23720 9460 23720 9460 5 FreeSans 1600 0 0 -800 res2
flabel metal2 12020 10770 12020 10770 1 FreeSans 1600 0 0 800 V_TOP
flabel metal2 10200 9320 10200 9320 1 FreeSans 1600 0 0 800 V_CUR_REF_REG
flabel metal2 10130 11210 10130 11210 1 FreeSans 1600 0 0 800 V1
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
