magic
tech sky130A
magscale 1 2
timestamp 1757090368
<< nwell >>
rect 33050 3340 35360 5570
<< pwell >>
rect 33050 1840 35170 3260
<< nmos >>
rect 33278 2840 33310 3040
rect 33798 2840 33830 3040
rect 34318 2840 34350 3040
rect 33280 2360 33310 2660
rect 33800 2360 33830 2660
rect 34320 2360 34350 2660
rect 33280 1980 33310 2180
rect 33800 1980 33830 2180
rect 34320 1980 34350 2180
rect 34920 1980 34950 2180
<< pmos >>
rect 33280 5030 33580 5430
rect 33800 5030 34100 5430
rect 34320 5030 34620 5430
rect 34840 5030 35140 5430
rect 33280 4140 33310 4740
rect 33800 4140 33830 4740
rect 34320 4140 34350 4740
rect 33278 3560 33310 3960
rect 33798 3560 33830 3960
rect 34318 3560 34350 3960
<< ndiff >>
rect 33198 3010 33278 3040
rect 33198 2970 33218 3010
rect 33258 2970 33278 3010
rect 33198 2910 33278 2970
rect 33198 2870 33218 2910
rect 33258 2870 33278 2910
rect 33198 2840 33278 2870
rect 33310 3010 33390 3040
rect 33310 2970 33330 3010
rect 33370 2970 33390 3010
rect 33310 2910 33390 2970
rect 33310 2870 33330 2910
rect 33370 2870 33390 2910
rect 33310 2840 33390 2870
rect 33718 3010 33798 3040
rect 33718 2970 33738 3010
rect 33778 2970 33798 3010
rect 33718 2910 33798 2970
rect 33718 2870 33738 2910
rect 33778 2870 33798 2910
rect 33718 2840 33798 2870
rect 33830 3010 33910 3040
rect 33830 2970 33850 3010
rect 33890 2970 33910 3010
rect 33830 2910 33910 2970
rect 33830 2870 33850 2910
rect 33890 2870 33910 2910
rect 33830 2840 33910 2870
rect 34238 3010 34318 3040
rect 34238 2970 34258 3010
rect 34298 2970 34318 3010
rect 34238 2910 34318 2970
rect 34238 2870 34258 2910
rect 34298 2870 34318 2910
rect 34238 2840 34318 2870
rect 34350 3010 34430 3040
rect 34350 2970 34370 3010
rect 34410 2970 34430 3010
rect 34350 2910 34430 2970
rect 34350 2870 34370 2910
rect 34410 2870 34430 2910
rect 34350 2840 34430 2870
rect 33200 2630 33280 2660
rect 33200 2590 33220 2630
rect 33260 2590 33280 2630
rect 33200 2530 33280 2590
rect 33200 2490 33220 2530
rect 33260 2490 33280 2530
rect 33200 2430 33280 2490
rect 33200 2390 33220 2430
rect 33260 2390 33280 2430
rect 33200 2360 33280 2390
rect 33310 2630 33390 2660
rect 33310 2590 33330 2630
rect 33370 2590 33390 2630
rect 33310 2530 33390 2590
rect 33310 2490 33330 2530
rect 33370 2490 33390 2530
rect 33310 2430 33390 2490
rect 33310 2390 33330 2430
rect 33370 2390 33390 2430
rect 33310 2360 33390 2390
rect 33720 2630 33800 2660
rect 33720 2590 33740 2630
rect 33780 2590 33800 2630
rect 33720 2530 33800 2590
rect 33720 2490 33740 2530
rect 33780 2490 33800 2530
rect 33720 2430 33800 2490
rect 33720 2390 33740 2430
rect 33780 2390 33800 2430
rect 33720 2360 33800 2390
rect 33830 2630 33910 2660
rect 33830 2590 33850 2630
rect 33890 2590 33910 2630
rect 33830 2530 33910 2590
rect 33830 2490 33850 2530
rect 33890 2490 33910 2530
rect 33830 2430 33910 2490
rect 33830 2390 33850 2430
rect 33890 2390 33910 2430
rect 33830 2360 33910 2390
rect 34240 2630 34320 2660
rect 34240 2590 34260 2630
rect 34300 2590 34320 2630
rect 34240 2530 34320 2590
rect 34240 2490 34260 2530
rect 34300 2490 34320 2530
rect 34240 2430 34320 2490
rect 34240 2390 34260 2430
rect 34300 2390 34320 2430
rect 34240 2360 34320 2390
rect 34350 2630 34430 2660
rect 34350 2590 34370 2630
rect 34410 2590 34430 2630
rect 34350 2530 34430 2590
rect 34350 2490 34370 2530
rect 34410 2490 34430 2530
rect 34350 2430 34430 2490
rect 34350 2390 34370 2430
rect 34410 2390 34430 2430
rect 34350 2360 34430 2390
rect 33200 2150 33280 2180
rect 33200 2110 33220 2150
rect 33260 2110 33280 2150
rect 33200 2050 33280 2110
rect 33200 2010 33220 2050
rect 33260 2010 33280 2050
rect 33200 1980 33280 2010
rect 33310 2150 33390 2180
rect 33310 2110 33330 2150
rect 33370 2110 33390 2150
rect 33310 2050 33390 2110
rect 33310 2010 33330 2050
rect 33370 2010 33390 2050
rect 33310 1980 33390 2010
rect 33720 2150 33800 2180
rect 33720 2110 33740 2150
rect 33780 2110 33800 2150
rect 33720 2050 33800 2110
rect 33720 2010 33740 2050
rect 33780 2010 33800 2050
rect 33720 1980 33800 2010
rect 33830 2150 33910 2180
rect 33830 2110 33850 2150
rect 33890 2110 33910 2150
rect 33830 2050 33910 2110
rect 33830 2010 33850 2050
rect 33890 2010 33910 2050
rect 33830 1980 33910 2010
rect 34240 2150 34320 2180
rect 34240 2110 34260 2150
rect 34300 2110 34320 2150
rect 34240 2050 34320 2110
rect 34240 2010 34260 2050
rect 34300 2010 34320 2050
rect 34240 1980 34320 2010
rect 34350 2150 34430 2180
rect 34350 2110 34370 2150
rect 34410 2110 34430 2150
rect 34350 2050 34430 2110
rect 34350 2010 34370 2050
rect 34410 2010 34430 2050
rect 34350 1980 34430 2010
rect 34840 2150 34920 2180
rect 34840 2110 34860 2150
rect 34900 2110 34920 2150
rect 34840 2050 34920 2110
rect 34840 2010 34860 2050
rect 34900 2010 34920 2050
rect 34840 1980 34920 2010
rect 34950 2150 35030 2180
rect 34950 2110 34970 2150
rect 35010 2110 35030 2150
rect 34950 2050 35030 2110
rect 34950 2010 34970 2050
rect 35010 2010 35030 2050
rect 34950 1980 35030 2010
<< pdiff >>
rect 33200 5400 33280 5430
rect 33200 5360 33220 5400
rect 33260 5360 33280 5400
rect 33200 5300 33280 5360
rect 33200 5260 33220 5300
rect 33260 5260 33280 5300
rect 33200 5200 33280 5260
rect 33200 5160 33220 5200
rect 33260 5160 33280 5200
rect 33200 5100 33280 5160
rect 33200 5060 33220 5100
rect 33260 5060 33280 5100
rect 33200 5030 33280 5060
rect 33580 5400 33660 5430
rect 33580 5360 33600 5400
rect 33640 5360 33660 5400
rect 33580 5300 33660 5360
rect 33580 5260 33600 5300
rect 33640 5260 33660 5300
rect 33580 5200 33660 5260
rect 33580 5160 33600 5200
rect 33640 5160 33660 5200
rect 33580 5100 33660 5160
rect 33580 5060 33600 5100
rect 33640 5060 33660 5100
rect 33580 5030 33660 5060
rect 33720 5400 33800 5430
rect 33720 5360 33740 5400
rect 33780 5360 33800 5400
rect 33720 5300 33800 5360
rect 33720 5260 33740 5300
rect 33780 5260 33800 5300
rect 33720 5200 33800 5260
rect 33720 5160 33740 5200
rect 33780 5160 33800 5200
rect 33720 5100 33800 5160
rect 33720 5060 33740 5100
rect 33780 5060 33800 5100
rect 33720 5030 33800 5060
rect 34100 5400 34180 5430
rect 34100 5360 34120 5400
rect 34160 5360 34180 5400
rect 34100 5300 34180 5360
rect 34100 5260 34120 5300
rect 34160 5260 34180 5300
rect 34100 5200 34180 5260
rect 34100 5160 34120 5200
rect 34160 5160 34180 5200
rect 34100 5100 34180 5160
rect 34100 5060 34120 5100
rect 34160 5060 34180 5100
rect 34100 5030 34180 5060
rect 34240 5400 34320 5430
rect 34240 5360 34260 5400
rect 34300 5360 34320 5400
rect 34240 5300 34320 5360
rect 34240 5260 34260 5300
rect 34300 5260 34320 5300
rect 34240 5200 34320 5260
rect 34240 5160 34260 5200
rect 34300 5160 34320 5200
rect 34240 5100 34320 5160
rect 34240 5060 34260 5100
rect 34300 5060 34320 5100
rect 34240 5030 34320 5060
rect 34620 5400 34700 5430
rect 34620 5360 34640 5400
rect 34680 5360 34700 5400
rect 34620 5300 34700 5360
rect 34620 5260 34640 5300
rect 34680 5260 34700 5300
rect 34620 5200 34700 5260
rect 34620 5160 34640 5200
rect 34680 5160 34700 5200
rect 34620 5100 34700 5160
rect 34620 5060 34640 5100
rect 34680 5060 34700 5100
rect 34620 5030 34700 5060
rect 34760 5400 34840 5430
rect 34760 5360 34780 5400
rect 34820 5360 34840 5400
rect 34760 5300 34840 5360
rect 34760 5260 34780 5300
rect 34820 5260 34840 5300
rect 34760 5200 34840 5260
rect 34760 5160 34780 5200
rect 34820 5160 34840 5200
rect 34760 5100 34840 5160
rect 34760 5060 34780 5100
rect 34820 5060 34840 5100
rect 34760 5030 34840 5060
rect 35140 5400 35220 5430
rect 35140 5360 35160 5400
rect 35200 5360 35220 5400
rect 35140 5300 35220 5360
rect 35140 5260 35160 5300
rect 35200 5260 35220 5300
rect 35140 5200 35220 5260
rect 35140 5160 35160 5200
rect 35200 5160 35220 5200
rect 35140 5100 35220 5160
rect 35140 5060 35160 5100
rect 35200 5060 35220 5100
rect 35140 5030 35220 5060
rect 33200 4710 33280 4740
rect 33200 4670 33220 4710
rect 33260 4670 33280 4710
rect 33200 4610 33280 4670
rect 33200 4570 33220 4610
rect 33260 4570 33280 4610
rect 33200 4510 33280 4570
rect 33200 4470 33220 4510
rect 33260 4470 33280 4510
rect 33200 4410 33280 4470
rect 33200 4370 33220 4410
rect 33260 4370 33280 4410
rect 33200 4310 33280 4370
rect 33200 4270 33220 4310
rect 33260 4270 33280 4310
rect 33200 4210 33280 4270
rect 33200 4170 33220 4210
rect 33260 4170 33280 4210
rect 33200 4140 33280 4170
rect 33310 4710 33390 4740
rect 33310 4670 33330 4710
rect 33370 4670 33390 4710
rect 33310 4610 33390 4670
rect 33310 4570 33330 4610
rect 33370 4570 33390 4610
rect 33310 4510 33390 4570
rect 33310 4470 33330 4510
rect 33370 4470 33390 4510
rect 33310 4410 33390 4470
rect 33310 4370 33330 4410
rect 33370 4370 33390 4410
rect 33310 4310 33390 4370
rect 33310 4270 33330 4310
rect 33370 4270 33390 4310
rect 33310 4210 33390 4270
rect 33310 4170 33330 4210
rect 33370 4170 33390 4210
rect 33310 4140 33390 4170
rect 33720 4710 33800 4740
rect 33720 4670 33740 4710
rect 33780 4670 33800 4710
rect 33720 4610 33800 4670
rect 33720 4570 33740 4610
rect 33780 4570 33800 4610
rect 33720 4510 33800 4570
rect 33720 4470 33740 4510
rect 33780 4470 33800 4510
rect 33720 4410 33800 4470
rect 33720 4370 33740 4410
rect 33780 4370 33800 4410
rect 33720 4310 33800 4370
rect 33720 4270 33740 4310
rect 33780 4270 33800 4310
rect 33720 4210 33800 4270
rect 33720 4170 33740 4210
rect 33780 4170 33800 4210
rect 33720 4140 33800 4170
rect 33830 4710 33910 4740
rect 33830 4670 33850 4710
rect 33890 4670 33910 4710
rect 33830 4610 33910 4670
rect 33830 4570 33850 4610
rect 33890 4570 33910 4610
rect 33830 4510 33910 4570
rect 33830 4470 33850 4510
rect 33890 4470 33910 4510
rect 33830 4410 33910 4470
rect 33830 4370 33850 4410
rect 33890 4370 33910 4410
rect 33830 4310 33910 4370
rect 33830 4270 33850 4310
rect 33890 4270 33910 4310
rect 33830 4210 33910 4270
rect 33830 4170 33850 4210
rect 33890 4170 33910 4210
rect 33830 4140 33910 4170
rect 34240 4710 34320 4740
rect 34240 4670 34260 4710
rect 34300 4670 34320 4710
rect 34240 4610 34320 4670
rect 34240 4570 34260 4610
rect 34300 4570 34320 4610
rect 34240 4510 34320 4570
rect 34240 4470 34260 4510
rect 34300 4470 34320 4510
rect 34240 4410 34320 4470
rect 34240 4370 34260 4410
rect 34300 4370 34320 4410
rect 34240 4310 34320 4370
rect 34240 4270 34260 4310
rect 34300 4270 34320 4310
rect 34240 4210 34320 4270
rect 34240 4170 34260 4210
rect 34300 4170 34320 4210
rect 34240 4140 34320 4170
rect 34350 4710 34430 4740
rect 34350 4670 34370 4710
rect 34410 4670 34430 4710
rect 34350 4610 34430 4670
rect 34350 4570 34370 4610
rect 34410 4570 34430 4610
rect 34350 4510 34430 4570
rect 34350 4470 34370 4510
rect 34410 4470 34430 4510
rect 34350 4410 34430 4470
rect 34350 4370 34370 4410
rect 34410 4370 34430 4410
rect 34350 4310 34430 4370
rect 34350 4270 34370 4310
rect 34410 4270 34430 4310
rect 34350 4210 34430 4270
rect 34350 4170 34370 4210
rect 34410 4170 34430 4210
rect 34350 4140 34430 4170
rect 33198 3930 33278 3960
rect 33198 3890 33218 3930
rect 33258 3890 33278 3930
rect 33198 3830 33278 3890
rect 33198 3790 33218 3830
rect 33258 3790 33278 3830
rect 33198 3730 33278 3790
rect 33198 3690 33218 3730
rect 33258 3690 33278 3730
rect 33198 3630 33278 3690
rect 33198 3590 33218 3630
rect 33258 3590 33278 3630
rect 33198 3560 33278 3590
rect 33310 3930 33390 3960
rect 33310 3890 33330 3930
rect 33370 3890 33390 3930
rect 33310 3830 33390 3890
rect 33310 3790 33330 3830
rect 33370 3790 33390 3830
rect 33310 3730 33390 3790
rect 33310 3690 33330 3730
rect 33370 3690 33390 3730
rect 33310 3630 33390 3690
rect 33310 3590 33330 3630
rect 33370 3590 33390 3630
rect 33310 3560 33390 3590
rect 33718 3930 33798 3960
rect 33718 3890 33738 3930
rect 33778 3890 33798 3930
rect 33718 3830 33798 3890
rect 33718 3790 33738 3830
rect 33778 3790 33798 3830
rect 33718 3730 33798 3790
rect 33718 3690 33738 3730
rect 33778 3690 33798 3730
rect 33718 3630 33798 3690
rect 33718 3590 33738 3630
rect 33778 3590 33798 3630
rect 33718 3560 33798 3590
rect 33830 3930 33910 3960
rect 33830 3890 33850 3930
rect 33890 3890 33910 3930
rect 33830 3830 33910 3890
rect 33830 3790 33850 3830
rect 33890 3790 33910 3830
rect 33830 3730 33910 3790
rect 33830 3690 33850 3730
rect 33890 3690 33910 3730
rect 33830 3630 33910 3690
rect 33830 3590 33850 3630
rect 33890 3590 33910 3630
rect 33830 3560 33910 3590
rect 34238 3930 34318 3960
rect 34238 3890 34258 3930
rect 34298 3890 34318 3930
rect 34238 3830 34318 3890
rect 34238 3790 34258 3830
rect 34298 3790 34318 3830
rect 34238 3730 34318 3790
rect 34238 3690 34258 3730
rect 34298 3690 34318 3730
rect 34238 3630 34318 3690
rect 34238 3590 34258 3630
rect 34298 3590 34318 3630
rect 34238 3560 34318 3590
rect 34350 3930 34430 3960
rect 34350 3890 34370 3930
rect 34410 3890 34430 3930
rect 34350 3830 34430 3890
rect 34350 3790 34370 3830
rect 34410 3790 34430 3830
rect 34350 3730 34430 3790
rect 34350 3690 34370 3730
rect 34410 3690 34430 3730
rect 34350 3630 34430 3690
rect 34350 3590 34370 3630
rect 34410 3590 34430 3630
rect 34350 3560 34430 3590
<< ndiffc >>
rect 33218 2970 33258 3010
rect 33218 2870 33258 2910
rect 33330 2970 33370 3010
rect 33330 2870 33370 2910
rect 33738 2970 33778 3010
rect 33738 2870 33778 2910
rect 33850 2970 33890 3010
rect 33850 2870 33890 2910
rect 34258 2970 34298 3010
rect 34258 2870 34298 2910
rect 34370 2970 34410 3010
rect 34370 2870 34410 2910
rect 33220 2590 33260 2630
rect 33220 2490 33260 2530
rect 33220 2390 33260 2430
rect 33330 2590 33370 2630
rect 33330 2490 33370 2530
rect 33330 2390 33370 2430
rect 33740 2590 33780 2630
rect 33740 2490 33780 2530
rect 33740 2390 33780 2430
rect 33850 2590 33890 2630
rect 33850 2490 33890 2530
rect 33850 2390 33890 2430
rect 34260 2590 34300 2630
rect 34260 2490 34300 2530
rect 34260 2390 34300 2430
rect 34370 2590 34410 2630
rect 34370 2490 34410 2530
rect 34370 2390 34410 2430
rect 33220 2110 33260 2150
rect 33220 2010 33260 2050
rect 33330 2110 33370 2150
rect 33330 2010 33370 2050
rect 33740 2110 33780 2150
rect 33740 2010 33780 2050
rect 33850 2110 33890 2150
rect 33850 2010 33890 2050
rect 34260 2110 34300 2150
rect 34260 2010 34300 2050
rect 34370 2110 34410 2150
rect 34370 2010 34410 2050
rect 34860 2110 34900 2150
rect 34860 2010 34900 2050
rect 34970 2110 35010 2150
rect 34970 2010 35010 2050
<< pdiffc >>
rect 33220 5360 33260 5400
rect 33220 5260 33260 5300
rect 33220 5160 33260 5200
rect 33220 5060 33260 5100
rect 33600 5360 33640 5400
rect 33600 5260 33640 5300
rect 33600 5160 33640 5200
rect 33600 5060 33640 5100
rect 33740 5360 33780 5400
rect 33740 5260 33780 5300
rect 33740 5160 33780 5200
rect 33740 5060 33780 5100
rect 34120 5360 34160 5400
rect 34120 5260 34160 5300
rect 34120 5160 34160 5200
rect 34120 5060 34160 5100
rect 34260 5360 34300 5400
rect 34260 5260 34300 5300
rect 34260 5160 34300 5200
rect 34260 5060 34300 5100
rect 34640 5360 34680 5400
rect 34640 5260 34680 5300
rect 34640 5160 34680 5200
rect 34640 5060 34680 5100
rect 34780 5360 34820 5400
rect 34780 5260 34820 5300
rect 34780 5160 34820 5200
rect 34780 5060 34820 5100
rect 35160 5360 35200 5400
rect 35160 5260 35200 5300
rect 35160 5160 35200 5200
rect 35160 5060 35200 5100
rect 33220 4670 33260 4710
rect 33220 4570 33260 4610
rect 33220 4470 33260 4510
rect 33220 4370 33260 4410
rect 33220 4270 33260 4310
rect 33220 4170 33260 4210
rect 33330 4670 33370 4710
rect 33330 4570 33370 4610
rect 33330 4470 33370 4510
rect 33330 4370 33370 4410
rect 33330 4270 33370 4310
rect 33330 4170 33370 4210
rect 33740 4670 33780 4710
rect 33740 4570 33780 4610
rect 33740 4470 33780 4510
rect 33740 4370 33780 4410
rect 33740 4270 33780 4310
rect 33740 4170 33780 4210
rect 33850 4670 33890 4710
rect 33850 4570 33890 4610
rect 33850 4470 33890 4510
rect 33850 4370 33890 4410
rect 33850 4270 33890 4310
rect 33850 4170 33890 4210
rect 34260 4670 34300 4710
rect 34260 4570 34300 4610
rect 34260 4470 34300 4510
rect 34260 4370 34300 4410
rect 34260 4270 34300 4310
rect 34260 4170 34300 4210
rect 34370 4670 34410 4710
rect 34370 4570 34410 4610
rect 34370 4470 34410 4510
rect 34370 4370 34410 4410
rect 34370 4270 34410 4310
rect 34370 4170 34410 4210
rect 33218 3890 33258 3930
rect 33218 3790 33258 3830
rect 33218 3690 33258 3730
rect 33218 3590 33258 3630
rect 33330 3890 33370 3930
rect 33330 3790 33370 3830
rect 33330 3690 33370 3730
rect 33330 3590 33370 3630
rect 33738 3890 33778 3930
rect 33738 3790 33778 3830
rect 33738 3690 33778 3730
rect 33738 3590 33778 3630
rect 33850 3890 33890 3930
rect 33850 3790 33890 3830
rect 33850 3690 33890 3730
rect 33850 3590 33890 3630
rect 34258 3890 34298 3930
rect 34258 3790 34298 3830
rect 34258 3690 34298 3730
rect 34258 3590 34298 3630
rect 34370 3890 34410 3930
rect 34370 3790 34410 3830
rect 34370 3690 34410 3730
rect 34370 3590 34410 3630
<< psubdiff >>
rect 33090 3180 34230 3220
rect 34370 3180 35130 3220
rect 33090 2660 33130 3180
rect 35090 2660 35130 3180
rect 33090 1920 33130 2450
rect 35090 1920 35130 2450
rect 33090 1880 34230 1920
rect 34370 1880 35130 1920
<< nsubdiff >>
rect 33090 5490 34110 5530
rect 34270 5490 35150 5530
rect 35220 5490 35320 5530
rect 33090 5060 33130 5490
rect 35280 5060 35320 5490
rect 33090 3420 33130 4730
rect 35280 3420 35320 4730
rect 33090 3380 34110 3420
rect 34270 3380 35320 3420
<< psubdiffcont >>
rect 34230 3180 34370 3220
rect 33090 2450 33130 2660
rect 35090 2450 35130 2660
rect 34230 1880 34370 1920
<< nsubdiffcont >>
rect 34110 5490 34270 5530
rect 35150 5490 35220 5530
rect 33090 4730 33130 5060
rect 35280 4730 35320 5060
rect 34110 3380 34270 3420
<< poly >>
rect 33280 5430 33580 5460
rect 33800 5430 34100 5460
rect 34320 5430 34620 5460
rect 34840 5430 35140 5460
rect 33280 5000 33580 5030
rect 33800 5000 34100 5030
rect 34320 5000 34620 5030
rect 34840 5000 35140 5030
rect 33390 4980 33470 5000
rect 33390 4940 33410 4980
rect 33450 4940 33470 4980
rect 33390 4920 33470 4940
rect 33910 4980 33990 5000
rect 33910 4940 33930 4980
rect 33970 4940 33990 4980
rect 33910 4920 33990 4940
rect 34430 4980 34510 5000
rect 34430 4940 34450 4980
rect 34490 4940 34510 4980
rect 34430 4920 34510 4940
rect 34960 4980 35020 5000
rect 34960 4940 34970 4980
rect 35010 4940 35020 4980
rect 34960 4920 35020 4940
rect 33280 4740 33310 4770
rect 33800 4740 33830 4770
rect 34320 4740 34350 4770
rect 33280 4110 33310 4140
rect 33800 4110 33830 4140
rect 34320 4110 34350 4140
rect 33280 4092 33338 4110
rect 33280 4058 33292 4092
rect 33326 4058 33338 4092
rect 33280 4040 33338 4058
rect 33800 4092 33858 4110
rect 33800 4058 33812 4092
rect 33846 4058 33858 4092
rect 33800 4040 33858 4058
rect 34320 4092 34378 4110
rect 34320 4058 34332 4092
rect 34366 4058 34378 4092
rect 34320 4040 34378 4058
rect 33278 3960 33310 3990
rect 33798 3960 33830 3990
rect 34318 3960 34350 3990
rect 33278 3530 33310 3560
rect 33798 3530 33830 3560
rect 34318 3530 34350 3560
rect 33252 3512 33310 3530
rect 33252 3478 33264 3512
rect 33298 3478 33310 3512
rect 33252 3460 33310 3478
rect 33772 3512 33830 3530
rect 33772 3478 33784 3512
rect 33818 3478 33830 3512
rect 33772 3460 33830 3478
rect 34292 3512 34350 3530
rect 34292 3478 34304 3512
rect 34338 3478 34350 3512
rect 34292 3460 34350 3478
rect 33252 3122 33310 3140
rect 33252 3088 33264 3122
rect 33298 3088 33310 3122
rect 33252 3070 33310 3088
rect 33772 3122 33830 3140
rect 33772 3088 33784 3122
rect 33818 3088 33830 3122
rect 33772 3070 33830 3088
rect 34292 3122 34350 3140
rect 34292 3088 34304 3122
rect 34338 3088 34350 3122
rect 34292 3070 34350 3088
rect 33278 3040 33310 3070
rect 33798 3040 33830 3070
rect 34318 3040 34350 3070
rect 33278 2810 33310 2840
rect 33798 2810 33830 2840
rect 34318 2810 34350 2840
rect 33280 2742 33338 2760
rect 33280 2708 33292 2742
rect 33326 2708 33338 2742
rect 33280 2690 33338 2708
rect 33800 2742 33858 2760
rect 33800 2708 33812 2742
rect 33846 2708 33858 2742
rect 33800 2690 33858 2708
rect 34320 2742 34378 2760
rect 34320 2708 34332 2742
rect 34366 2708 34378 2742
rect 34320 2690 34378 2708
rect 33280 2660 33310 2690
rect 33800 2660 33830 2690
rect 34320 2660 34350 2690
rect 33280 2330 33310 2360
rect 33800 2330 33830 2360
rect 34320 2330 34350 2360
rect 33266 2262 33324 2280
rect 33266 2228 33278 2262
rect 33312 2228 33324 2262
rect 33266 2210 33324 2228
rect 33786 2262 33844 2280
rect 33786 2228 33798 2262
rect 33832 2228 33844 2262
rect 33786 2210 33844 2228
rect 34306 2262 34364 2280
rect 34306 2228 34318 2262
rect 34352 2228 34364 2262
rect 34306 2210 34364 2228
rect 34874 2262 34950 2280
rect 34874 2228 34886 2262
rect 34920 2228 34950 2262
rect 34874 2210 34950 2228
rect 33280 2180 33310 2210
rect 33800 2180 33830 2210
rect 34320 2180 34350 2210
rect 34920 2180 34950 2210
rect 33280 1950 33310 1980
rect 33800 1950 33830 1980
rect 34320 1950 34350 1980
rect 34920 1950 34950 1980
<< polycont >>
rect 33410 4940 33450 4980
rect 33930 4940 33970 4980
rect 34450 4940 34490 4980
rect 34970 4940 35010 4980
rect 33292 4058 33326 4092
rect 33812 4058 33846 4092
rect 34332 4058 34366 4092
rect 33264 3478 33298 3512
rect 33784 3478 33818 3512
rect 34304 3478 34338 3512
rect 33264 3088 33298 3122
rect 33784 3088 33818 3122
rect 34304 3088 34338 3122
rect 33292 2708 33326 2742
rect 33812 2708 33846 2742
rect 34332 2708 34366 2742
rect 33278 2228 33312 2262
rect 33798 2228 33832 2262
rect 34318 2228 34352 2262
rect 34886 2228 34920 2262
<< locali >>
rect 33580 5530 33660 5550
rect 34100 5530 34180 5550
rect 34620 5530 34700 5550
rect 35140 5530 35220 5550
rect 33090 5490 33600 5530
rect 33640 5490 34110 5530
rect 34270 5490 34640 5530
rect 34680 5490 35150 5530
rect 35220 5490 35320 5530
rect 33090 5060 33130 5490
rect 33580 5470 33660 5490
rect 34100 5470 34180 5490
rect 34620 5470 34700 5490
rect 35140 5470 35220 5490
rect 33210 5400 33270 5420
rect 33210 5360 33220 5400
rect 33260 5360 33270 5400
rect 33210 5300 33270 5360
rect 33210 5260 33220 5300
rect 33260 5260 33270 5300
rect 33210 5200 33270 5260
rect 33210 5160 33220 5200
rect 33260 5160 33270 5200
rect 33210 5100 33270 5160
rect 33210 5060 33220 5100
rect 33260 5060 33270 5100
rect 33210 5040 33270 5060
rect 33590 5400 33650 5420
rect 33590 5360 33600 5400
rect 33640 5360 33650 5400
rect 33590 5300 33650 5360
rect 33590 5260 33600 5300
rect 33640 5260 33650 5300
rect 33590 5200 33650 5260
rect 33590 5160 33600 5200
rect 33640 5160 33650 5200
rect 33590 5100 33650 5160
rect 33590 5060 33600 5100
rect 33640 5060 33650 5100
rect 33590 5040 33650 5060
rect 33730 5400 33790 5420
rect 33730 5360 33740 5400
rect 33780 5360 33790 5400
rect 33730 5300 33790 5360
rect 33730 5260 33740 5300
rect 33780 5260 33790 5300
rect 33730 5200 33790 5260
rect 33730 5160 33740 5200
rect 33780 5160 33790 5200
rect 33730 5100 33790 5160
rect 33730 5060 33740 5100
rect 33780 5060 33790 5100
rect 33730 5040 33790 5060
rect 34110 5400 34170 5420
rect 34110 5360 34120 5400
rect 34160 5360 34170 5400
rect 34110 5300 34170 5360
rect 34110 5260 34120 5300
rect 34160 5260 34170 5300
rect 34110 5200 34170 5260
rect 34110 5160 34120 5200
rect 34160 5160 34170 5200
rect 34110 5100 34170 5160
rect 34110 5060 34120 5100
rect 34160 5060 34170 5100
rect 34110 5040 34170 5060
rect 34250 5400 34310 5420
rect 34250 5360 34260 5400
rect 34300 5360 34310 5400
rect 34250 5300 34310 5360
rect 34250 5260 34260 5300
rect 34300 5260 34310 5300
rect 34250 5200 34310 5260
rect 34250 5160 34260 5200
rect 34300 5160 34310 5200
rect 34250 5100 34310 5160
rect 34250 5060 34260 5100
rect 34300 5060 34310 5100
rect 34250 5040 34310 5060
rect 34630 5400 34690 5420
rect 34630 5360 34640 5400
rect 34680 5360 34690 5400
rect 34630 5300 34690 5360
rect 34630 5260 34640 5300
rect 34680 5260 34690 5300
rect 34630 5200 34690 5260
rect 34630 5160 34640 5200
rect 34680 5160 34690 5200
rect 34630 5100 34690 5160
rect 34630 5060 34640 5100
rect 34680 5060 34690 5100
rect 34630 5040 34690 5060
rect 34770 5400 34830 5420
rect 34770 5360 34780 5400
rect 34820 5360 34830 5400
rect 34770 5300 34830 5360
rect 34770 5260 34780 5300
rect 34820 5260 34830 5300
rect 34770 5200 34830 5260
rect 34770 5160 34780 5200
rect 34820 5160 34830 5200
rect 34770 5100 34830 5160
rect 34770 5060 34780 5100
rect 34820 5060 34830 5100
rect 34770 5040 34830 5060
rect 35150 5400 35210 5420
rect 35150 5360 35160 5400
rect 35200 5360 35210 5400
rect 35150 5300 35210 5360
rect 35150 5260 35160 5300
rect 35200 5260 35210 5300
rect 35150 5200 35210 5260
rect 35150 5160 35160 5200
rect 35200 5160 35210 5200
rect 35150 5100 35210 5160
rect 35150 5060 35160 5100
rect 35200 5060 35210 5100
rect 35150 5040 35210 5060
rect 35280 5060 35320 5490
rect 33390 4980 33470 5000
rect 33390 4940 33410 4980
rect 33450 4940 33470 4980
rect 33390 4920 33470 4940
rect 33910 4980 33990 5000
rect 33910 4940 33930 4980
rect 33970 4940 33990 4980
rect 33910 4920 33990 4940
rect 34430 4980 34510 5000
rect 34430 4940 34450 4980
rect 34490 4940 34510 4980
rect 34430 4920 34510 4940
rect 34960 4980 35020 5000
rect 34960 4940 34970 4980
rect 35010 4940 35020 4980
rect 34960 4920 35020 4940
rect 33090 3420 33130 4730
rect 33210 4710 33270 4730
rect 33210 4670 33220 4710
rect 33260 4670 33270 4710
rect 33210 4610 33270 4670
rect 33210 4570 33220 4610
rect 33260 4570 33270 4610
rect 33210 4510 33270 4570
rect 33210 4470 33220 4510
rect 33260 4470 33270 4510
rect 33210 4410 33270 4470
rect 33210 4370 33220 4410
rect 33260 4370 33270 4410
rect 33210 4310 33270 4370
rect 33210 4270 33220 4310
rect 33260 4270 33270 4310
rect 33210 4210 33270 4270
rect 33210 4170 33220 4210
rect 33260 4170 33270 4210
rect 33210 4150 33270 4170
rect 33320 4710 33380 4730
rect 33320 4670 33330 4710
rect 33370 4670 33380 4710
rect 33320 4610 33380 4670
rect 33320 4570 33330 4610
rect 33370 4570 33380 4610
rect 33320 4510 33380 4570
rect 33320 4470 33330 4510
rect 33370 4470 33380 4510
rect 33320 4410 33380 4470
rect 33320 4370 33330 4410
rect 33370 4370 33380 4410
rect 33320 4310 33380 4370
rect 33320 4270 33330 4310
rect 33370 4270 33380 4310
rect 33320 4210 33380 4270
rect 33320 4170 33330 4210
rect 33370 4170 33380 4210
rect 33320 4150 33380 4170
rect 33730 4710 33790 4730
rect 33730 4670 33740 4710
rect 33780 4670 33790 4710
rect 33730 4610 33790 4670
rect 33730 4570 33740 4610
rect 33780 4570 33790 4610
rect 33730 4510 33790 4570
rect 33730 4470 33740 4510
rect 33780 4470 33790 4510
rect 33730 4410 33790 4470
rect 33730 4370 33740 4410
rect 33780 4370 33790 4410
rect 33730 4310 33790 4370
rect 33730 4270 33740 4310
rect 33780 4270 33790 4310
rect 33730 4210 33790 4270
rect 33730 4170 33740 4210
rect 33780 4170 33790 4210
rect 33730 4150 33790 4170
rect 33840 4710 33900 4730
rect 33840 4670 33850 4710
rect 33890 4670 33900 4710
rect 33840 4610 33900 4670
rect 33840 4570 33850 4610
rect 33890 4570 33900 4610
rect 33840 4510 33900 4570
rect 33840 4470 33850 4510
rect 33890 4470 33900 4510
rect 33840 4410 33900 4470
rect 33840 4370 33850 4410
rect 33890 4370 33900 4410
rect 33840 4310 33900 4370
rect 33840 4270 33850 4310
rect 33890 4270 33900 4310
rect 33840 4210 33900 4270
rect 33840 4170 33850 4210
rect 33890 4170 33900 4210
rect 33840 4150 33900 4170
rect 34250 4710 34310 4730
rect 34250 4670 34260 4710
rect 34300 4670 34310 4710
rect 34250 4610 34310 4670
rect 34250 4570 34260 4610
rect 34300 4570 34310 4610
rect 34250 4510 34310 4570
rect 34250 4470 34260 4510
rect 34300 4470 34310 4510
rect 34250 4410 34310 4470
rect 34250 4370 34260 4410
rect 34300 4370 34310 4410
rect 34250 4310 34310 4370
rect 34250 4270 34260 4310
rect 34300 4270 34310 4310
rect 34250 4210 34310 4270
rect 34250 4170 34260 4210
rect 34300 4170 34310 4210
rect 34250 4150 34310 4170
rect 34360 4710 34420 4730
rect 34360 4670 34370 4710
rect 34410 4670 34420 4710
rect 34360 4610 34420 4670
rect 34360 4570 34370 4610
rect 34410 4570 34420 4610
rect 34360 4510 34420 4570
rect 34360 4470 34370 4510
rect 34410 4470 34420 4510
rect 34360 4410 34420 4470
rect 34360 4370 34370 4410
rect 34410 4370 34420 4410
rect 34360 4310 34420 4370
rect 34360 4270 34370 4310
rect 34410 4270 34420 4310
rect 34360 4210 34420 4270
rect 34360 4170 34370 4210
rect 34410 4170 34420 4210
rect 34360 4150 34420 4170
rect 33280 4092 33338 4110
rect 33280 4058 33292 4092
rect 33326 4058 33338 4092
rect 33280 4040 33338 4058
rect 33800 4092 33858 4110
rect 33800 4058 33812 4092
rect 33846 4058 33858 4092
rect 33800 4040 33858 4058
rect 34320 4092 34378 4110
rect 34320 4058 34332 4092
rect 34366 4058 34378 4092
rect 34320 4040 34378 4058
rect 33208 3930 33268 3950
rect 33208 3890 33218 3930
rect 33258 3890 33268 3930
rect 33208 3830 33268 3890
rect 33208 3790 33218 3830
rect 33258 3790 33268 3830
rect 33208 3730 33268 3790
rect 33208 3690 33218 3730
rect 33258 3690 33268 3730
rect 33208 3630 33268 3690
rect 33208 3590 33218 3630
rect 33258 3590 33268 3630
rect 33208 3570 33268 3590
rect 33320 3930 33380 3950
rect 33320 3890 33330 3930
rect 33370 3890 33380 3930
rect 33320 3830 33380 3890
rect 33320 3790 33330 3830
rect 33370 3790 33380 3830
rect 33320 3730 33380 3790
rect 33320 3690 33330 3730
rect 33370 3690 33380 3730
rect 33320 3630 33380 3690
rect 33320 3590 33330 3630
rect 33370 3590 33380 3630
rect 33320 3570 33380 3590
rect 33728 3930 33788 3950
rect 33728 3890 33738 3930
rect 33778 3890 33788 3930
rect 33728 3830 33788 3890
rect 33728 3790 33738 3830
rect 33778 3790 33788 3830
rect 33728 3730 33788 3790
rect 33728 3690 33738 3730
rect 33778 3690 33788 3730
rect 33728 3630 33788 3690
rect 33728 3590 33738 3630
rect 33778 3590 33788 3630
rect 33728 3570 33788 3590
rect 33840 3930 33900 3950
rect 33840 3890 33850 3930
rect 33890 3890 33900 3930
rect 33840 3830 33900 3890
rect 33840 3790 33850 3830
rect 33890 3790 33900 3830
rect 33840 3730 33900 3790
rect 33840 3690 33850 3730
rect 33890 3690 33900 3730
rect 33840 3630 33900 3690
rect 33840 3590 33850 3630
rect 33890 3590 33900 3630
rect 33840 3570 33900 3590
rect 34248 3930 34308 3950
rect 34248 3890 34258 3930
rect 34298 3890 34308 3930
rect 34248 3830 34308 3890
rect 34248 3790 34258 3830
rect 34298 3790 34308 3830
rect 34248 3730 34308 3790
rect 34248 3690 34258 3730
rect 34298 3690 34308 3730
rect 34248 3630 34308 3690
rect 34248 3590 34258 3630
rect 34298 3590 34308 3630
rect 34248 3570 34308 3590
rect 34360 3930 34420 3950
rect 34360 3890 34370 3930
rect 34410 3890 34420 3930
rect 34360 3830 34420 3890
rect 34360 3790 34370 3830
rect 34410 3790 34420 3830
rect 34360 3730 34420 3790
rect 34360 3690 34370 3730
rect 34410 3690 34420 3730
rect 34360 3630 34420 3690
rect 34360 3590 34370 3630
rect 34410 3590 34420 3630
rect 34360 3570 34420 3590
rect 33252 3512 33310 3530
rect 33252 3478 33264 3512
rect 33298 3478 33310 3512
rect 33252 3460 33310 3478
rect 33772 3512 33830 3530
rect 33772 3478 33784 3512
rect 33818 3478 33830 3512
rect 33772 3460 33830 3478
rect 34292 3512 34350 3530
rect 34292 3478 34304 3512
rect 34338 3478 34350 3512
rect 34292 3460 34350 3478
rect 35280 3420 35320 4730
rect 33090 3380 34110 3420
rect 34270 3380 35320 3420
rect 33090 3180 34230 3220
rect 34370 3180 35130 3220
rect 33090 2660 33130 3180
rect 33252 3122 33310 3140
rect 33252 3088 33264 3122
rect 33298 3088 33310 3122
rect 33252 3070 33310 3088
rect 33772 3122 33830 3140
rect 33772 3088 33784 3122
rect 33818 3088 33830 3122
rect 33772 3070 33830 3088
rect 34292 3122 34350 3140
rect 34292 3088 34304 3122
rect 34338 3088 34350 3122
rect 34292 3070 34350 3088
rect 33208 3010 33268 3030
rect 33208 2970 33218 3010
rect 33258 2970 33268 3010
rect 33208 2910 33268 2970
rect 33208 2870 33218 2910
rect 33258 2870 33268 2910
rect 33208 2850 33268 2870
rect 33320 3010 33380 3030
rect 33320 2970 33330 3010
rect 33370 2970 33380 3010
rect 33320 2910 33380 2970
rect 33320 2870 33330 2910
rect 33370 2870 33380 2910
rect 33320 2850 33380 2870
rect 33728 3010 33788 3030
rect 33728 2970 33738 3010
rect 33778 2970 33788 3010
rect 33728 2910 33788 2970
rect 33728 2870 33738 2910
rect 33778 2870 33788 2910
rect 33728 2850 33788 2870
rect 33840 3010 33900 3030
rect 33840 2970 33850 3010
rect 33890 2970 33900 3010
rect 33840 2910 33900 2970
rect 33840 2870 33850 2910
rect 33890 2870 33900 2910
rect 33840 2850 33900 2870
rect 34248 3010 34308 3030
rect 34248 2970 34258 3010
rect 34298 2970 34308 3010
rect 34248 2910 34308 2970
rect 34248 2870 34258 2910
rect 34298 2870 34308 2910
rect 34248 2850 34308 2870
rect 34360 3010 34420 3030
rect 34360 2970 34370 3010
rect 34410 2970 34420 3010
rect 34360 2910 34420 2970
rect 34360 2870 34370 2910
rect 34410 2870 34420 2910
rect 34360 2850 34420 2870
rect 33280 2742 33338 2760
rect 33280 2708 33292 2742
rect 33326 2708 33338 2742
rect 33280 2690 33338 2708
rect 33800 2742 33858 2760
rect 33800 2708 33812 2742
rect 33846 2708 33858 2742
rect 33800 2690 33858 2708
rect 34320 2742 34378 2760
rect 34320 2708 34332 2742
rect 34366 2708 34378 2742
rect 34320 2690 34378 2708
rect 35090 2660 35130 3180
rect 33090 1920 33130 2450
rect 33210 2630 33270 2650
rect 33210 2590 33220 2630
rect 33260 2590 33270 2630
rect 33210 2530 33270 2590
rect 33210 2490 33220 2530
rect 33260 2490 33270 2530
rect 33210 2430 33270 2490
rect 33210 2390 33220 2430
rect 33260 2390 33270 2430
rect 33210 2370 33270 2390
rect 33320 2630 33380 2650
rect 33320 2590 33330 2630
rect 33370 2590 33380 2630
rect 33320 2530 33380 2590
rect 33320 2490 33330 2530
rect 33370 2490 33380 2530
rect 33320 2430 33380 2490
rect 33320 2390 33330 2430
rect 33370 2390 33380 2430
rect 33320 2370 33380 2390
rect 33730 2630 33790 2650
rect 33730 2590 33740 2630
rect 33780 2590 33790 2630
rect 33730 2530 33790 2590
rect 33730 2490 33740 2530
rect 33780 2490 33790 2530
rect 33730 2430 33790 2490
rect 33730 2390 33740 2430
rect 33780 2390 33790 2430
rect 33730 2370 33790 2390
rect 33840 2630 33900 2650
rect 33840 2590 33850 2630
rect 33890 2590 33900 2630
rect 33840 2530 33900 2590
rect 33840 2490 33850 2530
rect 33890 2490 33900 2530
rect 33840 2430 33900 2490
rect 33840 2390 33850 2430
rect 33890 2390 33900 2430
rect 33840 2370 33900 2390
rect 34250 2630 34310 2650
rect 34250 2590 34260 2630
rect 34300 2590 34310 2630
rect 34250 2530 34310 2590
rect 34250 2490 34260 2530
rect 34300 2490 34310 2530
rect 34250 2430 34310 2490
rect 34250 2390 34260 2430
rect 34300 2390 34310 2430
rect 34250 2370 34310 2390
rect 34360 2630 34420 2650
rect 34360 2590 34370 2630
rect 34410 2590 34420 2630
rect 34360 2530 34420 2590
rect 34360 2490 34370 2530
rect 34410 2490 34420 2530
rect 34360 2430 34420 2490
rect 34360 2390 34370 2430
rect 34410 2390 34420 2430
rect 34360 2370 34420 2390
rect 33266 2262 33324 2280
rect 33266 2228 33278 2262
rect 33312 2228 33324 2262
rect 33266 2210 33324 2228
rect 33786 2262 33844 2280
rect 33786 2228 33798 2262
rect 33832 2228 33844 2262
rect 33786 2210 33844 2228
rect 34306 2262 34364 2280
rect 34306 2228 34318 2262
rect 34352 2228 34364 2262
rect 34306 2210 34364 2228
rect 34874 2262 34932 2280
rect 34874 2228 34886 2262
rect 34920 2228 34932 2262
rect 34874 2210 34932 2228
rect 33210 2150 33270 2170
rect 33210 2110 33220 2150
rect 33260 2110 33270 2150
rect 33210 2050 33270 2110
rect 33210 2010 33220 2050
rect 33260 2010 33270 2050
rect 33210 1990 33270 2010
rect 33320 2150 33380 2170
rect 33320 2110 33330 2150
rect 33370 2110 33380 2150
rect 33320 2050 33380 2110
rect 33320 2010 33330 2050
rect 33370 2010 33380 2050
rect 33320 1990 33380 2010
rect 33730 2150 33790 2170
rect 33730 2110 33740 2150
rect 33780 2110 33790 2150
rect 33730 2050 33790 2110
rect 33730 2010 33740 2050
rect 33780 2010 33790 2050
rect 33730 1990 33790 2010
rect 33840 2150 33900 2170
rect 33840 2110 33850 2150
rect 33890 2110 33900 2150
rect 33840 2050 33900 2110
rect 33840 2010 33850 2050
rect 33890 2010 33900 2050
rect 33840 1990 33900 2010
rect 34250 2150 34310 2170
rect 34250 2110 34260 2150
rect 34300 2110 34310 2150
rect 34250 2050 34310 2110
rect 34250 2010 34260 2050
rect 34300 2010 34310 2050
rect 34250 1990 34310 2010
rect 34360 2150 34420 2170
rect 34360 2110 34370 2150
rect 34410 2110 34420 2150
rect 34360 2050 34420 2110
rect 34360 2010 34370 2050
rect 34410 2010 34420 2050
rect 34360 1990 34420 2010
rect 34850 2150 34910 2170
rect 34850 2110 34860 2150
rect 34900 2110 34910 2150
rect 34850 2050 34910 2110
rect 34850 2010 34860 2050
rect 34900 2010 34910 2050
rect 34850 1990 34910 2010
rect 34960 2150 35020 2170
rect 34960 2110 34970 2150
rect 35010 2110 35020 2150
rect 34960 2050 35020 2110
rect 34960 2010 34970 2050
rect 35010 2010 35020 2050
rect 34960 1990 35020 2010
rect 33310 1920 33390 1940
rect 33830 1920 33910 1940
rect 34350 1920 34430 1940
rect 34840 1920 34920 1940
rect 35090 1920 35130 2450
rect 33090 1880 33330 1920
rect 33370 1880 33850 1920
rect 33890 1880 34230 1920
rect 34410 1880 34860 1920
rect 34900 1880 35130 1920
rect 33310 1860 33390 1880
rect 33830 1860 33910 1880
rect 34350 1860 34430 1880
rect 34840 1860 34920 1880
<< viali >>
rect 33600 5490 33640 5530
rect 34120 5490 34160 5530
rect 34640 5490 34680 5530
rect 35160 5490 35200 5530
rect 33220 5360 33260 5400
rect 33220 5260 33260 5300
rect 33220 5160 33260 5200
rect 33220 5060 33260 5100
rect 33600 5360 33640 5400
rect 33600 5260 33640 5300
rect 33600 5160 33640 5200
rect 33600 5060 33640 5100
rect 33740 5360 33780 5400
rect 33740 5260 33780 5300
rect 33740 5160 33780 5200
rect 33740 5060 33780 5100
rect 34120 5360 34160 5400
rect 34120 5260 34160 5300
rect 34120 5160 34160 5200
rect 34120 5060 34160 5100
rect 34260 5360 34300 5400
rect 34260 5260 34300 5300
rect 34260 5160 34300 5200
rect 34260 5060 34300 5100
rect 34640 5360 34680 5400
rect 34640 5260 34680 5300
rect 34640 5160 34680 5200
rect 34640 5060 34680 5100
rect 34780 5360 34820 5400
rect 34780 5260 34820 5300
rect 34780 5160 34820 5200
rect 34780 5060 34820 5100
rect 35160 5360 35200 5400
rect 35160 5260 35200 5300
rect 35160 5160 35200 5200
rect 35160 5060 35200 5100
rect 33410 4940 33450 4980
rect 33930 4940 33970 4980
rect 34450 4940 34490 4980
rect 34970 4940 35010 4980
rect 33220 4670 33260 4710
rect 33220 4570 33260 4610
rect 33220 4470 33260 4510
rect 33220 4370 33260 4410
rect 33220 4270 33260 4310
rect 33220 4170 33260 4210
rect 33330 4670 33370 4710
rect 33330 4570 33370 4610
rect 33330 4470 33370 4510
rect 33330 4370 33370 4410
rect 33330 4270 33370 4310
rect 33330 4170 33370 4210
rect 33740 4670 33780 4710
rect 33740 4570 33780 4610
rect 33740 4470 33780 4510
rect 33740 4370 33780 4410
rect 33740 4270 33780 4310
rect 33740 4170 33780 4210
rect 33850 4670 33890 4710
rect 33850 4570 33890 4610
rect 33850 4470 33890 4510
rect 33850 4370 33890 4410
rect 33850 4270 33890 4310
rect 33850 4170 33890 4210
rect 34260 4670 34300 4710
rect 34260 4570 34300 4610
rect 34260 4470 34300 4510
rect 34260 4370 34300 4410
rect 34260 4270 34300 4310
rect 34260 4170 34300 4210
rect 34370 4670 34410 4710
rect 34370 4570 34410 4610
rect 34370 4470 34410 4510
rect 34370 4370 34410 4410
rect 34370 4270 34410 4310
rect 34370 4170 34410 4210
rect 33292 4058 33326 4092
rect 33812 4058 33846 4092
rect 34332 4058 34366 4092
rect 33218 3890 33258 3930
rect 33218 3790 33258 3830
rect 33218 3690 33258 3730
rect 33218 3590 33258 3630
rect 33330 3890 33370 3930
rect 33330 3790 33370 3830
rect 33330 3690 33370 3730
rect 33330 3590 33370 3630
rect 33738 3890 33778 3930
rect 33738 3790 33778 3830
rect 33738 3690 33778 3730
rect 33738 3590 33778 3630
rect 33850 3890 33890 3930
rect 33850 3790 33890 3830
rect 33850 3690 33890 3730
rect 33850 3590 33890 3630
rect 34258 3890 34298 3930
rect 34258 3790 34298 3830
rect 34258 3690 34298 3730
rect 34258 3590 34298 3630
rect 34370 3890 34410 3930
rect 34370 3790 34410 3830
rect 34370 3690 34410 3730
rect 34370 3590 34410 3630
rect 33264 3478 33298 3512
rect 33784 3478 33818 3512
rect 34304 3478 34338 3512
rect 33264 3088 33298 3122
rect 33784 3088 33818 3122
rect 34304 3088 34338 3122
rect 33218 2970 33258 3010
rect 33218 2870 33258 2910
rect 33330 2970 33370 3010
rect 33330 2870 33370 2910
rect 33738 2970 33778 3010
rect 33738 2870 33778 2910
rect 33850 2970 33890 3010
rect 33850 2870 33890 2910
rect 34258 2970 34298 3010
rect 34258 2870 34298 2910
rect 34370 2970 34410 3010
rect 34370 2870 34410 2910
rect 33292 2708 33326 2742
rect 33812 2708 33846 2742
rect 34332 2708 34366 2742
rect 33220 2590 33260 2630
rect 33220 2490 33260 2530
rect 33220 2390 33260 2430
rect 33330 2590 33370 2630
rect 33330 2490 33370 2530
rect 33330 2390 33370 2430
rect 33740 2590 33780 2630
rect 33740 2490 33780 2530
rect 33740 2390 33780 2430
rect 33850 2590 33890 2630
rect 33850 2490 33890 2530
rect 33850 2390 33890 2430
rect 34260 2590 34300 2630
rect 34260 2490 34300 2530
rect 34260 2390 34300 2430
rect 34370 2590 34410 2630
rect 34370 2490 34410 2530
rect 34370 2390 34410 2430
rect 33278 2228 33312 2262
rect 33798 2228 33832 2262
rect 34318 2228 34352 2262
rect 34886 2228 34920 2262
rect 33220 2110 33260 2150
rect 33220 2010 33260 2050
rect 33330 2110 33370 2150
rect 33330 2010 33370 2050
rect 33740 2110 33780 2150
rect 33740 2010 33780 2050
rect 33850 2110 33890 2150
rect 33850 2010 33890 2050
rect 34260 2110 34300 2150
rect 34260 2010 34300 2050
rect 34370 2110 34410 2150
rect 34370 2010 34410 2050
rect 34860 2110 34900 2150
rect 34860 2010 34900 2050
rect 34970 2110 35010 2150
rect 34970 2010 35010 2050
rect 33330 1880 33370 1920
rect 33850 1880 33890 1920
rect 34370 1880 34410 1920
rect 34860 1880 34900 1920
<< metal1 >>
rect 33580 5640 33660 5650
rect 33580 5580 33590 5640
rect 33650 5580 33660 5640
rect 33580 5530 33660 5580
rect 33580 5490 33600 5530
rect 33640 5490 33660 5530
rect 33580 5470 33660 5490
rect 34100 5640 34180 5650
rect 34100 5580 34110 5640
rect 34170 5580 34180 5640
rect 34100 5530 34180 5580
rect 34100 5490 34120 5530
rect 34160 5490 34180 5530
rect 34100 5470 34180 5490
rect 34620 5640 34700 5650
rect 34620 5580 34630 5640
rect 34690 5580 34700 5640
rect 34620 5530 34700 5580
rect 34620 5490 34640 5530
rect 34680 5490 34700 5530
rect 34620 5470 34700 5490
rect 35140 5640 35220 5650
rect 35140 5580 35150 5640
rect 35210 5580 35220 5640
rect 35140 5530 35220 5580
rect 35140 5490 35160 5530
rect 35200 5490 35220 5530
rect 35140 5470 35220 5490
rect 33210 5400 33270 5420
rect 33210 5360 33220 5400
rect 33260 5360 33270 5400
rect 33210 5300 33270 5360
rect 33210 5260 33220 5300
rect 33260 5260 33270 5300
rect 33210 5200 33270 5260
rect 33210 5160 33220 5200
rect 33260 5160 33270 5200
rect 33210 5100 33270 5160
rect 33210 5060 33220 5100
rect 33260 5060 33270 5100
rect 33210 4710 33270 5060
rect 33590 5400 33650 5470
rect 33590 5360 33600 5400
rect 33640 5360 33650 5400
rect 33590 5300 33650 5360
rect 33590 5260 33600 5300
rect 33640 5260 33650 5300
rect 33590 5200 33650 5260
rect 33590 5160 33600 5200
rect 33640 5160 33650 5200
rect 33590 5100 33650 5160
rect 33590 5060 33600 5100
rect 33640 5060 33650 5100
rect 33390 4990 33470 5000
rect 33390 4930 33400 4990
rect 33460 4930 33470 4990
rect 33390 4920 33470 4930
rect 33590 4820 33650 5060
rect 33730 5400 33790 5420
rect 33730 5360 33740 5400
rect 33780 5360 33790 5400
rect 33730 5300 33790 5360
rect 33730 5260 33740 5300
rect 33780 5260 33790 5300
rect 33730 5200 33790 5260
rect 33730 5160 33740 5200
rect 33780 5160 33790 5200
rect 33730 5100 33790 5160
rect 33730 5060 33740 5100
rect 33780 5060 33790 5100
rect 33310 4810 33390 4820
rect 33310 4750 33320 4810
rect 33380 4750 33390 4810
rect 33310 4740 33390 4750
rect 33580 4810 33660 4820
rect 33580 4750 33590 4810
rect 33650 4750 33660 4810
rect 33580 4740 33660 4750
rect 33210 4670 33220 4710
rect 33260 4670 33270 4710
rect 33210 4610 33270 4670
rect 33210 4570 33220 4610
rect 33260 4570 33270 4610
rect 33210 4510 33270 4570
rect 33210 4470 33220 4510
rect 33260 4470 33270 4510
rect 33210 4410 33270 4470
rect 33210 4370 33220 4410
rect 33260 4370 33270 4410
rect 33210 4310 33270 4370
rect 33210 4270 33220 4310
rect 33260 4270 33270 4310
rect 33210 4210 33270 4270
rect 33210 4170 33220 4210
rect 33260 4170 33270 4210
rect 33210 4150 33270 4170
rect 33320 4710 33380 4740
rect 33320 4670 33330 4710
rect 33370 4670 33380 4710
rect 33320 4610 33380 4670
rect 33320 4570 33330 4610
rect 33370 4570 33380 4610
rect 33320 4510 33380 4570
rect 33320 4470 33330 4510
rect 33370 4470 33380 4510
rect 33320 4410 33380 4470
rect 33320 4370 33330 4410
rect 33370 4370 33380 4410
rect 33320 4310 33380 4370
rect 33320 4270 33330 4310
rect 33370 4270 33380 4310
rect 33320 4220 33380 4270
rect 33730 4710 33790 5060
rect 34110 5400 34170 5470
rect 34110 5360 34120 5400
rect 34160 5360 34170 5400
rect 34110 5300 34170 5360
rect 34110 5260 34120 5300
rect 34160 5260 34170 5300
rect 34110 5200 34170 5260
rect 34110 5160 34120 5200
rect 34160 5160 34170 5200
rect 34110 5100 34170 5160
rect 34110 5060 34120 5100
rect 34160 5060 34170 5100
rect 33910 4990 33990 5000
rect 33910 4930 33920 4990
rect 33980 4930 33990 4990
rect 33910 4920 33990 4930
rect 34110 4820 34170 5060
rect 34250 5400 34310 5420
rect 34250 5360 34260 5400
rect 34300 5360 34310 5400
rect 34250 5300 34310 5360
rect 34250 5260 34260 5300
rect 34300 5260 34310 5300
rect 34250 5200 34310 5260
rect 34250 5160 34260 5200
rect 34300 5160 34310 5200
rect 34250 5100 34310 5160
rect 34250 5060 34260 5100
rect 34300 5060 34310 5100
rect 33830 4810 33910 4820
rect 33830 4750 33840 4810
rect 33900 4750 33910 4810
rect 33830 4740 33910 4750
rect 34100 4810 34180 4820
rect 34100 4750 34110 4810
rect 34170 4750 34180 4810
rect 34100 4740 34180 4750
rect 33730 4670 33740 4710
rect 33780 4670 33790 4710
rect 33730 4610 33790 4670
rect 33730 4570 33740 4610
rect 33780 4570 33790 4610
rect 33730 4510 33790 4570
rect 33730 4470 33740 4510
rect 33780 4470 33790 4510
rect 33730 4410 33790 4470
rect 33730 4370 33740 4410
rect 33780 4370 33790 4410
rect 33730 4310 33790 4370
rect 33730 4270 33740 4310
rect 33780 4270 33790 4310
rect 33320 4150 33380 4160
rect 33410 4220 33490 4230
rect 33410 4160 33420 4220
rect 33480 4160 33490 4220
rect 33410 4150 33490 4160
rect 33210 3950 33250 4150
rect 33280 4100 33338 4110
rect 33280 4048 33284 4100
rect 33336 4048 33338 4100
rect 33280 4040 33338 4048
rect 33208 3930 33268 3950
rect 33208 3890 33218 3930
rect 33258 3890 33268 3930
rect 33208 3830 33268 3890
rect 33208 3790 33218 3830
rect 33258 3790 33268 3830
rect 33208 3730 33268 3790
rect 33208 3690 33218 3730
rect 33258 3690 33268 3730
rect 33208 3630 33268 3690
rect 33208 3590 33218 3630
rect 33258 3590 33268 3630
rect 33208 3570 33268 3590
rect 33320 3930 33380 3950
rect 33320 3890 33330 3930
rect 33370 3890 33380 3930
rect 33320 3830 33380 3890
rect 33320 3790 33330 3830
rect 33370 3790 33380 3830
rect 33320 3730 33380 3790
rect 33320 3690 33330 3730
rect 33370 3690 33380 3730
rect 33320 3630 33380 3690
rect 33320 3590 33330 3630
rect 33370 3590 33380 3630
rect 33320 3560 33380 3590
rect 33252 3512 33310 3530
rect 33252 3478 33264 3512
rect 33298 3478 33310 3512
rect 33252 3460 33310 3478
rect 33260 3420 33310 3460
rect 32810 3410 33050 3420
rect 32810 3350 32820 3410
rect 32880 3350 32900 3410
rect 32960 3350 32980 3410
rect 33040 3350 33050 3410
rect 32810 3330 33050 3350
rect 32810 3270 32820 3330
rect 32880 3270 32900 3330
rect 32960 3270 32980 3330
rect 33040 3270 33050 3330
rect 32810 3250 33050 3270
rect 32810 3190 32820 3250
rect 32880 3190 32900 3250
rect 32960 3190 32980 3250
rect 33040 3190 33050 3250
rect 32810 1830 33050 3190
rect 33250 3410 33310 3420
rect 33250 3330 33310 3350
rect 33250 3250 33310 3270
rect 33250 3180 33310 3190
rect 33260 3140 33310 3180
rect 33252 3122 33310 3140
rect 33252 3088 33264 3122
rect 33298 3088 33310 3122
rect 33252 3070 33310 3088
rect 33340 3420 33380 3560
rect 33340 3410 33400 3420
rect 33340 3330 33400 3350
rect 33340 3250 33400 3270
rect 33340 3180 33400 3190
rect 33340 3030 33380 3180
rect 33170 3010 33268 3030
rect 33170 2970 33218 3010
rect 33258 2970 33268 3010
rect 33170 2910 33268 2970
rect 33170 2870 33218 2910
rect 33258 2870 33268 2910
rect 33170 2850 33268 2870
rect 33320 3010 33380 3030
rect 33320 2970 33330 3010
rect 33370 2970 33380 3010
rect 33320 2910 33380 2970
rect 33320 2870 33330 2910
rect 33370 2870 33380 2910
rect 33320 2850 33380 2870
rect 33170 2800 33212 2850
rect 33170 2650 33210 2800
rect 33430 2770 33490 4150
rect 33730 4210 33790 4270
rect 33730 4170 33740 4210
rect 33780 4170 33790 4210
rect 33730 4150 33790 4170
rect 33840 4710 33900 4740
rect 33840 4670 33850 4710
rect 33890 4670 33900 4710
rect 33840 4610 33900 4670
rect 33840 4570 33850 4610
rect 33890 4570 33900 4610
rect 33840 4510 33900 4570
rect 33840 4470 33850 4510
rect 33890 4470 33900 4510
rect 33840 4410 33900 4470
rect 33840 4370 33850 4410
rect 33890 4370 33900 4410
rect 33840 4310 33900 4370
rect 33840 4270 33850 4310
rect 33890 4270 33900 4310
rect 33840 4220 33900 4270
rect 34250 4710 34310 5060
rect 34630 5400 34690 5470
rect 34630 5360 34640 5400
rect 34680 5360 34690 5400
rect 34630 5300 34690 5360
rect 34630 5260 34640 5300
rect 34680 5260 34690 5300
rect 34630 5200 34690 5260
rect 34630 5160 34640 5200
rect 34680 5160 34690 5200
rect 34630 5100 34690 5160
rect 34630 5060 34640 5100
rect 34680 5060 34690 5100
rect 34430 4990 34510 5000
rect 34430 4930 34440 4990
rect 34500 4930 34510 4990
rect 34430 4920 34510 4930
rect 34630 4820 34690 5060
rect 34770 5400 34830 5420
rect 34770 5360 34780 5400
rect 34820 5360 34830 5400
rect 34770 5300 34830 5360
rect 34770 5260 34780 5300
rect 34820 5260 34830 5300
rect 34770 5200 34830 5260
rect 34770 5160 34780 5200
rect 34820 5160 34830 5200
rect 34770 5100 34830 5160
rect 34770 5060 34780 5100
rect 34820 5060 34830 5100
rect 34770 4990 34830 5060
rect 35150 5400 35210 5470
rect 35150 5360 35160 5400
rect 35200 5360 35210 5400
rect 35150 5300 35210 5360
rect 35150 5260 35160 5300
rect 35200 5260 35210 5300
rect 35150 5200 35210 5260
rect 35150 5160 35160 5200
rect 35200 5160 35210 5200
rect 35150 5100 35210 5160
rect 35150 5060 35160 5100
rect 35200 5060 35210 5100
rect 35150 5040 35210 5060
rect 34770 4920 34830 4930
rect 34960 4990 35020 5000
rect 34350 4810 34430 4820
rect 34350 4750 34360 4810
rect 34420 4750 34430 4810
rect 34350 4740 34430 4750
rect 34620 4810 34700 4820
rect 34620 4750 34630 4810
rect 34690 4750 34700 4810
rect 34620 4740 34700 4750
rect 34250 4670 34260 4710
rect 34300 4670 34310 4710
rect 34250 4610 34310 4670
rect 34250 4570 34260 4610
rect 34300 4570 34310 4610
rect 34250 4510 34310 4570
rect 34250 4470 34260 4510
rect 34300 4470 34310 4510
rect 34250 4410 34310 4470
rect 34250 4370 34260 4410
rect 34300 4370 34310 4410
rect 34250 4310 34310 4370
rect 34250 4270 34260 4310
rect 34300 4270 34310 4310
rect 33840 4150 33900 4160
rect 33930 4220 34010 4230
rect 33930 4160 33940 4220
rect 34000 4160 34010 4220
rect 33930 4150 34010 4160
rect 33410 2760 33490 2770
rect 33280 2750 33338 2760
rect 33280 2698 33284 2750
rect 33336 2698 33338 2750
rect 33280 2690 33338 2698
rect 33410 2700 33420 2760
rect 33480 2700 33490 2760
rect 33410 2690 33490 2700
rect 33520 4100 33600 4110
rect 33520 4040 33530 4100
rect 33590 4040 33600 4100
rect 33170 2630 33270 2650
rect 33170 2590 33220 2630
rect 33260 2590 33270 2630
rect 33170 2530 33270 2590
rect 33170 2490 33220 2530
rect 33260 2490 33270 2530
rect 33170 2430 33270 2490
rect 33170 2390 33220 2430
rect 33260 2390 33270 2430
rect 33170 2370 33270 2390
rect 33320 2640 33420 2650
rect 33380 2580 33420 2640
rect 33320 2530 33420 2580
rect 33520 2640 33600 4040
rect 33730 3950 33770 4150
rect 33800 4100 33858 4110
rect 33800 4048 33804 4100
rect 33856 4048 33858 4100
rect 33800 4040 33858 4048
rect 33728 3930 33788 3950
rect 33728 3890 33738 3930
rect 33778 3890 33788 3930
rect 33728 3830 33788 3890
rect 33728 3790 33738 3830
rect 33778 3790 33788 3830
rect 33728 3730 33788 3790
rect 33728 3690 33738 3730
rect 33778 3690 33788 3730
rect 33728 3630 33788 3690
rect 33728 3590 33738 3630
rect 33778 3590 33788 3630
rect 33728 3570 33788 3590
rect 33840 3930 33900 3950
rect 33840 3890 33850 3930
rect 33890 3890 33900 3930
rect 33840 3830 33900 3890
rect 33840 3790 33850 3830
rect 33890 3790 33900 3830
rect 33840 3730 33900 3790
rect 33840 3690 33850 3730
rect 33890 3690 33900 3730
rect 33840 3630 33900 3690
rect 33840 3590 33850 3630
rect 33890 3590 33900 3630
rect 33840 3560 33900 3590
rect 33772 3512 33830 3530
rect 33772 3478 33784 3512
rect 33818 3478 33830 3512
rect 33772 3460 33830 3478
rect 33780 3420 33830 3460
rect 33770 3410 33830 3420
rect 33770 3330 33830 3350
rect 33770 3250 33830 3270
rect 33770 3180 33830 3190
rect 33780 3140 33830 3180
rect 33772 3122 33830 3140
rect 33772 3088 33784 3122
rect 33818 3088 33830 3122
rect 33772 3070 33830 3088
rect 33860 3420 33900 3560
rect 33860 3410 33920 3420
rect 33860 3330 33920 3350
rect 33860 3250 33920 3270
rect 33860 3180 33920 3190
rect 33860 3030 33900 3180
rect 33520 2580 33530 2640
rect 33590 2580 33600 2640
rect 33520 2570 33600 2580
rect 33690 3010 33788 3030
rect 33690 2970 33738 3010
rect 33778 2970 33788 3010
rect 33690 2910 33788 2970
rect 33690 2870 33738 2910
rect 33778 2870 33788 2910
rect 33690 2850 33788 2870
rect 33840 3010 33900 3030
rect 33840 2970 33850 3010
rect 33890 2970 33900 3010
rect 33840 2910 33900 2970
rect 33840 2870 33850 2910
rect 33890 2870 33900 2910
rect 33840 2850 33900 2870
rect 33690 2800 33732 2850
rect 33690 2650 33730 2800
rect 33950 2770 34010 4150
rect 34250 4210 34310 4270
rect 34250 4170 34260 4210
rect 34300 4170 34310 4210
rect 34250 4150 34310 4170
rect 34360 4710 34420 4740
rect 34360 4670 34370 4710
rect 34410 4670 34420 4710
rect 34360 4610 34420 4670
rect 34360 4570 34370 4610
rect 34410 4570 34420 4610
rect 34360 4510 34420 4570
rect 34360 4470 34370 4510
rect 34410 4470 34420 4510
rect 34360 4410 34420 4470
rect 34360 4370 34370 4410
rect 34410 4370 34420 4410
rect 34360 4310 34420 4370
rect 34360 4270 34370 4310
rect 34410 4270 34420 4310
rect 34360 4220 34420 4270
rect 34360 4150 34420 4160
rect 34450 4220 34530 4230
rect 34450 4160 34460 4220
rect 34520 4160 34530 4220
rect 34450 4150 34530 4160
rect 33930 2760 34010 2770
rect 33800 2750 33858 2760
rect 33800 2698 33804 2750
rect 33856 2698 33858 2750
rect 33800 2690 33858 2698
rect 33930 2700 33940 2760
rect 34000 2700 34010 2760
rect 33930 2690 34010 2700
rect 34040 4100 34120 4110
rect 34040 4040 34050 4100
rect 34110 4040 34120 4100
rect 33690 2630 33790 2650
rect 33690 2590 33740 2630
rect 33780 2590 33790 2630
rect 33320 2490 33330 2530
rect 33370 2490 33420 2530
rect 33320 2430 33420 2490
rect 33320 2390 33330 2430
rect 33370 2390 33420 2430
rect 33320 2370 33420 2390
rect 33170 2170 33210 2370
rect 33266 2270 33324 2280
rect 33266 2218 33270 2270
rect 33322 2218 33324 2270
rect 33266 2210 33324 2218
rect 33380 2170 33420 2370
rect 33170 2150 33270 2170
rect 33170 2110 33220 2150
rect 33260 2110 33270 2150
rect 33170 2050 33270 2110
rect 33170 2010 33220 2050
rect 33260 2010 33270 2050
rect 33170 1990 33270 2010
rect 33320 2150 33420 2170
rect 33320 2110 33330 2150
rect 33370 2110 33420 2150
rect 33320 2050 33420 2110
rect 33320 2010 33330 2050
rect 33370 2010 33420 2050
rect 33320 1990 33420 2010
rect 33690 2530 33790 2590
rect 33690 2490 33740 2530
rect 33780 2490 33790 2530
rect 33690 2430 33790 2490
rect 33690 2390 33740 2430
rect 33780 2390 33790 2430
rect 33690 2370 33790 2390
rect 33840 2640 33940 2650
rect 33900 2580 33940 2640
rect 33840 2530 33940 2580
rect 34040 2640 34120 4040
rect 34250 3950 34290 4150
rect 34320 4100 34378 4110
rect 34320 4048 34324 4100
rect 34376 4048 34378 4100
rect 34320 4040 34378 4048
rect 34248 3930 34308 3950
rect 34248 3890 34258 3930
rect 34298 3890 34308 3930
rect 34248 3830 34308 3890
rect 34248 3790 34258 3830
rect 34298 3790 34308 3830
rect 34248 3730 34308 3790
rect 34248 3690 34258 3730
rect 34298 3690 34308 3730
rect 34248 3630 34308 3690
rect 34248 3590 34258 3630
rect 34298 3590 34308 3630
rect 34248 3570 34308 3590
rect 34360 3930 34420 3950
rect 34360 3890 34370 3930
rect 34410 3890 34420 3930
rect 34360 3830 34420 3890
rect 34360 3790 34370 3830
rect 34410 3790 34420 3830
rect 34360 3730 34420 3790
rect 34360 3690 34370 3730
rect 34410 3690 34420 3730
rect 34360 3630 34420 3690
rect 34360 3590 34370 3630
rect 34410 3590 34420 3630
rect 34360 3560 34420 3590
rect 34292 3512 34350 3530
rect 34292 3478 34304 3512
rect 34338 3478 34350 3512
rect 34292 3460 34350 3478
rect 34300 3420 34350 3460
rect 34290 3410 34350 3420
rect 34290 3330 34350 3350
rect 34290 3250 34350 3270
rect 34290 3180 34350 3190
rect 34300 3140 34350 3180
rect 34292 3122 34350 3140
rect 34292 3088 34304 3122
rect 34338 3088 34350 3122
rect 34292 3070 34350 3088
rect 34380 3420 34420 3560
rect 34380 3410 34440 3420
rect 34380 3330 34440 3350
rect 34380 3250 34440 3270
rect 34380 3180 34440 3190
rect 34380 3030 34420 3180
rect 34040 2580 34050 2640
rect 34110 2580 34120 2640
rect 34040 2570 34120 2580
rect 34210 3010 34308 3030
rect 34210 2970 34258 3010
rect 34298 2970 34308 3010
rect 34210 2910 34308 2970
rect 34210 2870 34258 2910
rect 34298 2870 34308 2910
rect 34210 2850 34308 2870
rect 34360 3010 34420 3030
rect 34360 2970 34370 3010
rect 34410 2970 34420 3010
rect 34360 2910 34420 2970
rect 34360 2870 34370 2910
rect 34410 2870 34420 2910
rect 34360 2850 34420 2870
rect 34210 2800 34252 2850
rect 34210 2650 34250 2800
rect 34470 2770 34530 4150
rect 34450 2760 34530 2770
rect 34320 2750 34378 2760
rect 34320 2698 34324 2750
rect 34376 2698 34378 2750
rect 34320 2690 34378 2698
rect 34450 2700 34460 2760
rect 34520 2700 34530 2760
rect 34450 2690 34530 2700
rect 34560 4100 34640 4110
rect 34560 4040 34570 4100
rect 34630 4040 34640 4100
rect 34210 2630 34310 2650
rect 34210 2590 34260 2630
rect 34300 2590 34310 2630
rect 33840 2490 33850 2530
rect 33890 2490 33940 2530
rect 33840 2430 33940 2490
rect 33840 2390 33850 2430
rect 33890 2390 33940 2430
rect 33840 2370 33940 2390
rect 33690 2170 33730 2370
rect 33786 2270 33844 2280
rect 33786 2218 33790 2270
rect 33842 2218 33844 2270
rect 33786 2210 33844 2218
rect 33900 2170 33940 2370
rect 33690 2150 33790 2170
rect 33690 2110 33740 2150
rect 33780 2110 33790 2150
rect 33690 2050 33790 2110
rect 33690 2010 33740 2050
rect 33780 2010 33790 2050
rect 33690 1990 33790 2010
rect 33840 2150 33940 2170
rect 33840 2110 33850 2150
rect 33890 2110 33940 2150
rect 33840 2050 33940 2110
rect 33840 2010 33850 2050
rect 33890 2010 33940 2050
rect 33840 1990 33940 2010
rect 34210 2530 34310 2590
rect 34210 2490 34260 2530
rect 34300 2490 34310 2530
rect 34210 2430 34310 2490
rect 34210 2390 34260 2430
rect 34300 2390 34310 2430
rect 34210 2370 34310 2390
rect 34360 2640 34460 2650
rect 34420 2580 34460 2640
rect 34360 2530 34460 2580
rect 34560 2640 34640 4040
rect 34560 2580 34570 2640
rect 34630 2580 34640 2640
rect 34560 2570 34640 2580
rect 34360 2490 34370 2530
rect 34410 2490 34460 2530
rect 34360 2430 34460 2490
rect 34360 2390 34370 2430
rect 34410 2390 34460 2430
rect 34360 2370 34460 2390
rect 34210 2170 34250 2370
rect 34306 2270 34364 2280
rect 34306 2218 34310 2270
rect 34362 2218 34364 2270
rect 34306 2210 34364 2218
rect 34420 2170 34460 2370
rect 34874 2270 34932 2280
rect 34874 2218 34876 2270
rect 34928 2218 34932 2270
rect 34874 2210 34932 2218
rect 34210 2150 34310 2170
rect 34210 2110 34260 2150
rect 34300 2110 34310 2150
rect 34210 2050 34310 2110
rect 34210 2010 34260 2050
rect 34300 2010 34310 2050
rect 34210 1990 34310 2010
rect 34360 2150 34460 2170
rect 34360 2110 34370 2150
rect 34410 2110 34460 2150
rect 34360 2050 34460 2110
rect 34360 2010 34370 2050
rect 34410 2010 34460 2050
rect 34360 1990 34460 2010
rect 34850 2150 34910 2170
rect 34850 2110 34860 2150
rect 34900 2110 34910 2150
rect 34850 2050 34910 2110
rect 34850 2010 34860 2050
rect 34900 2010 34910 2050
rect 33320 1940 33380 1990
rect 33840 1940 33900 1990
rect 34360 1940 34420 1990
rect 34850 1940 34910 2010
rect 34960 2150 35020 4930
rect 34960 2110 34970 2150
rect 35010 2110 35020 2150
rect 34960 2050 35020 2110
rect 34960 2010 34970 2050
rect 35010 2010 35020 2050
rect 34960 1990 35020 2010
rect 35170 3410 35410 3420
rect 35170 3350 35180 3410
rect 35240 3350 35260 3410
rect 35320 3350 35340 3410
rect 35400 3350 35410 3410
rect 35170 3330 35410 3350
rect 35170 3270 35180 3330
rect 35240 3270 35260 3330
rect 35320 3270 35340 3330
rect 35400 3270 35410 3330
rect 35170 3250 35410 3270
rect 35170 3190 35180 3250
rect 35240 3190 35260 3250
rect 35320 3190 35340 3250
rect 35400 3190 35410 3250
rect 32810 1770 32820 1830
rect 32880 1770 32900 1830
rect 32960 1770 32980 1830
rect 33040 1770 33050 1830
rect 32810 1750 33050 1770
rect 32810 1690 32820 1750
rect 32880 1690 32900 1750
rect 32960 1690 32980 1750
rect 33040 1690 33050 1750
rect 32810 1670 33050 1690
rect 32810 1610 32820 1670
rect 32880 1610 32900 1670
rect 32960 1610 32980 1670
rect 33040 1610 33050 1670
rect 32810 1600 33050 1610
rect 33310 1920 33390 1940
rect 33310 1880 33330 1920
rect 33370 1880 33390 1920
rect 33310 1560 33390 1880
rect 33310 1500 33320 1560
rect 33380 1500 33390 1560
rect 33310 1490 33390 1500
rect 33830 1920 33910 1940
rect 33830 1880 33850 1920
rect 33890 1880 33910 1920
rect 33830 1560 33910 1880
rect 33830 1500 33840 1560
rect 33900 1500 33910 1560
rect 33830 1490 33910 1500
rect 34350 1920 34430 1940
rect 34350 1880 34370 1920
rect 34410 1880 34430 1920
rect 34350 1560 34430 1880
rect 34350 1500 34360 1560
rect 34420 1500 34430 1560
rect 34350 1490 34430 1500
rect 34840 1920 34920 1940
rect 34840 1880 34860 1920
rect 34900 1880 34920 1920
rect 34840 1560 34920 1880
rect 35170 1830 35410 3190
rect 35170 1770 35180 1830
rect 35240 1770 35260 1830
rect 35320 1770 35340 1830
rect 35400 1770 35410 1830
rect 35170 1750 35410 1770
rect 35170 1690 35180 1750
rect 35240 1690 35260 1750
rect 35320 1690 35340 1750
rect 35400 1690 35410 1750
rect 35170 1670 35410 1690
rect 35170 1610 35180 1670
rect 35240 1610 35260 1670
rect 35320 1610 35340 1670
rect 35400 1610 35410 1670
rect 35170 1600 35410 1610
rect 34840 1500 34850 1560
rect 34910 1500 34920 1560
rect 34840 1490 34920 1500
<< via1 >>
rect 33590 5580 33650 5640
rect 34110 5580 34170 5640
rect 34630 5580 34690 5640
rect 35150 5580 35210 5640
rect 33400 4980 33460 4990
rect 33400 4940 33410 4980
rect 33410 4940 33450 4980
rect 33450 4940 33460 4980
rect 33400 4930 33460 4940
rect 33320 4750 33380 4810
rect 33590 4750 33650 4810
rect 33920 4980 33980 4990
rect 33920 4940 33930 4980
rect 33930 4940 33970 4980
rect 33970 4940 33980 4980
rect 33920 4930 33980 4940
rect 33840 4750 33900 4810
rect 34110 4750 34170 4810
rect 33320 4210 33380 4220
rect 33320 4170 33330 4210
rect 33330 4170 33370 4210
rect 33370 4170 33380 4210
rect 33320 4160 33380 4170
rect 33420 4160 33480 4220
rect 33284 4092 33336 4100
rect 33284 4058 33292 4092
rect 33292 4058 33326 4092
rect 33326 4058 33336 4092
rect 33284 4048 33336 4058
rect 32820 3350 32880 3410
rect 32900 3350 32960 3410
rect 32980 3350 33040 3410
rect 32820 3270 32880 3330
rect 32900 3270 32960 3330
rect 32980 3270 33040 3330
rect 32820 3190 32880 3250
rect 32900 3190 32960 3250
rect 32980 3190 33040 3250
rect 33250 3350 33310 3410
rect 33250 3270 33310 3330
rect 33250 3190 33310 3250
rect 33340 3350 33400 3410
rect 33340 3270 33400 3330
rect 33340 3190 33400 3250
rect 34440 4980 34500 4990
rect 34440 4940 34450 4980
rect 34450 4940 34490 4980
rect 34490 4940 34500 4980
rect 34440 4930 34500 4940
rect 34770 4930 34830 4990
rect 34960 4980 35020 4990
rect 34960 4940 34970 4980
rect 34970 4940 35010 4980
rect 35010 4940 35020 4980
rect 34960 4930 35020 4940
rect 34360 4750 34420 4810
rect 34630 4750 34690 4810
rect 33840 4210 33900 4220
rect 33840 4170 33850 4210
rect 33850 4170 33890 4210
rect 33890 4170 33900 4210
rect 33840 4160 33900 4170
rect 33940 4160 34000 4220
rect 33284 2742 33336 2750
rect 33284 2708 33292 2742
rect 33292 2708 33326 2742
rect 33326 2708 33336 2742
rect 33284 2698 33336 2708
rect 33420 2700 33480 2760
rect 33530 4040 33590 4100
rect 33320 2630 33380 2640
rect 33320 2590 33330 2630
rect 33330 2590 33370 2630
rect 33370 2590 33380 2630
rect 33320 2580 33380 2590
rect 33804 4092 33856 4100
rect 33804 4058 33812 4092
rect 33812 4058 33846 4092
rect 33846 4058 33856 4092
rect 33804 4048 33856 4058
rect 33770 3350 33830 3410
rect 33770 3270 33830 3330
rect 33770 3190 33830 3250
rect 33860 3350 33920 3410
rect 33860 3270 33920 3330
rect 33860 3190 33920 3250
rect 33530 2580 33590 2640
rect 34360 4210 34420 4220
rect 34360 4170 34370 4210
rect 34370 4170 34410 4210
rect 34410 4170 34420 4210
rect 34360 4160 34420 4170
rect 34460 4160 34520 4220
rect 33804 2742 33856 2750
rect 33804 2708 33812 2742
rect 33812 2708 33846 2742
rect 33846 2708 33856 2742
rect 33804 2698 33856 2708
rect 33940 2700 34000 2760
rect 34050 4040 34110 4100
rect 33270 2262 33322 2270
rect 33270 2228 33278 2262
rect 33278 2228 33312 2262
rect 33312 2228 33322 2262
rect 33270 2218 33322 2228
rect 33840 2630 33900 2640
rect 33840 2590 33850 2630
rect 33850 2590 33890 2630
rect 33890 2590 33900 2630
rect 33840 2580 33900 2590
rect 34324 4092 34376 4100
rect 34324 4058 34332 4092
rect 34332 4058 34366 4092
rect 34366 4058 34376 4092
rect 34324 4048 34376 4058
rect 34290 3350 34350 3410
rect 34290 3270 34350 3330
rect 34290 3190 34350 3250
rect 34380 3350 34440 3410
rect 34380 3270 34440 3330
rect 34380 3190 34440 3250
rect 34050 2580 34110 2640
rect 34324 2742 34376 2750
rect 34324 2708 34332 2742
rect 34332 2708 34366 2742
rect 34366 2708 34376 2742
rect 34324 2698 34376 2708
rect 34460 2700 34520 2760
rect 34570 4040 34630 4100
rect 33790 2262 33842 2270
rect 33790 2228 33798 2262
rect 33798 2228 33832 2262
rect 33832 2228 33842 2262
rect 33790 2218 33842 2228
rect 34360 2630 34420 2640
rect 34360 2590 34370 2630
rect 34370 2590 34410 2630
rect 34410 2590 34420 2630
rect 34360 2580 34420 2590
rect 34570 2580 34630 2640
rect 34310 2262 34362 2270
rect 34310 2228 34318 2262
rect 34318 2228 34352 2262
rect 34352 2228 34362 2262
rect 34310 2218 34362 2228
rect 34876 2262 34928 2270
rect 34876 2228 34886 2262
rect 34886 2228 34920 2262
rect 34920 2228 34928 2262
rect 34876 2218 34928 2228
rect 35180 3350 35240 3410
rect 35260 3350 35320 3410
rect 35340 3350 35400 3410
rect 35180 3270 35240 3330
rect 35260 3270 35320 3330
rect 35340 3270 35400 3330
rect 35180 3190 35240 3250
rect 35260 3190 35320 3250
rect 35340 3190 35400 3250
rect 32820 1770 32880 1830
rect 32900 1770 32960 1830
rect 32980 1770 33040 1830
rect 32820 1690 32880 1750
rect 32900 1690 32960 1750
rect 32980 1690 33040 1750
rect 32820 1610 32880 1670
rect 32900 1610 32960 1670
rect 32980 1610 33040 1670
rect 33320 1500 33380 1560
rect 33840 1500 33900 1560
rect 34360 1500 34420 1560
rect 35180 1770 35240 1830
rect 35260 1770 35320 1830
rect 35340 1770 35400 1830
rect 35180 1690 35240 1750
rect 35260 1690 35320 1750
rect 35340 1690 35400 1750
rect 35180 1610 35240 1670
rect 35260 1610 35320 1670
rect 35340 1610 35400 1670
rect 34850 1500 34910 1560
<< metal2 >>
rect 33580 5640 35220 5650
rect 33580 5580 33590 5640
rect 33650 5580 34110 5640
rect 34170 5580 34630 5640
rect 34690 5580 35150 5640
rect 35210 5580 35220 5640
rect 33580 5570 35220 5580
rect 33390 4990 35020 5000
rect 33390 4930 33400 4990
rect 33460 4930 33920 4990
rect 33980 4930 34440 4990
rect 34500 4930 34770 4990
rect 34830 4930 34960 4990
rect 33390 4920 35020 4930
rect 33310 4810 33660 4820
rect 33310 4750 33320 4810
rect 33380 4750 33590 4810
rect 33650 4750 33660 4810
rect 33310 4740 33660 4750
rect 33830 4810 34180 4820
rect 33830 4750 33840 4810
rect 33900 4750 34110 4810
rect 34170 4750 34180 4810
rect 33830 4740 34180 4750
rect 34350 4810 34700 4820
rect 34350 4750 34360 4810
rect 34420 4750 34630 4810
rect 34690 4750 34700 4810
rect 34350 4740 34700 4750
rect 33320 4220 33490 4230
rect 33380 4160 33420 4220
rect 33480 4160 33490 4220
rect 33320 4150 33490 4160
rect 33840 4220 34010 4230
rect 33900 4160 33940 4220
rect 34000 4160 34010 4220
rect 33840 4150 34010 4160
rect 34360 4220 34530 4230
rect 34420 4160 34460 4220
rect 34520 4160 34530 4220
rect 34360 4150 34530 4160
rect 33280 4100 33600 4110
rect 33280 4048 33284 4100
rect 33336 4048 33530 4100
rect 33280 4040 33530 4048
rect 33590 4040 33600 4100
rect 33800 4100 34120 4110
rect 33800 4048 33804 4100
rect 33856 4048 34050 4100
rect 33800 4040 34050 4048
rect 34110 4040 34120 4100
rect 34320 4100 34640 4110
rect 34320 4048 34324 4100
rect 34376 4048 34570 4100
rect 34320 4040 34570 4048
rect 34630 4040 34640 4100
rect 33520 4030 33600 4040
rect 34040 4030 34120 4040
rect 34560 4030 34640 4040
rect 32810 3410 33310 3420
rect 32810 3350 32820 3410
rect 32880 3350 32900 3410
rect 32960 3350 32980 3410
rect 33040 3350 33250 3410
rect 32810 3330 33310 3350
rect 32810 3270 32820 3330
rect 32880 3270 32900 3330
rect 32960 3270 32980 3330
rect 33040 3270 33250 3330
rect 32810 3250 33310 3270
rect 32810 3190 32820 3250
rect 32880 3190 32900 3250
rect 32960 3190 32980 3250
rect 33040 3190 33250 3250
rect 32810 3180 33310 3190
rect 33340 3410 33830 3420
rect 33400 3350 33770 3410
rect 33340 3330 33830 3350
rect 33400 3270 33770 3330
rect 33340 3250 33830 3270
rect 33400 3190 33770 3250
rect 33340 3180 33830 3190
rect 33860 3410 34350 3420
rect 33920 3350 34290 3410
rect 33860 3330 34350 3350
rect 33920 3270 34290 3330
rect 33860 3250 34350 3270
rect 33920 3190 34290 3250
rect 33860 3180 34350 3190
rect 34380 3410 35410 3420
rect 34440 3350 35180 3410
rect 35240 3350 35260 3410
rect 35320 3350 35340 3410
rect 35400 3350 35410 3410
rect 34380 3330 35410 3350
rect 34440 3270 35180 3330
rect 35240 3270 35260 3330
rect 35320 3270 35340 3330
rect 35400 3270 35410 3330
rect 34380 3250 35410 3270
rect 34440 3190 35180 3250
rect 35240 3190 35260 3250
rect 35320 3190 35340 3250
rect 35400 3190 35410 3250
rect 34380 3180 35410 3190
rect 33410 2760 33490 2770
rect 33930 2760 34010 2770
rect 34450 2760 34530 2770
rect 33280 2750 33420 2760
rect 33280 2698 33284 2750
rect 33336 2700 33420 2750
rect 33480 2700 33490 2760
rect 33336 2698 33490 2700
rect 33280 2690 33490 2698
rect 33800 2750 33940 2760
rect 33800 2698 33804 2750
rect 33856 2700 33940 2750
rect 34000 2700 34010 2760
rect 33856 2698 34010 2700
rect 33800 2690 34010 2698
rect 34320 2750 34460 2760
rect 34320 2698 34324 2750
rect 34376 2700 34460 2750
rect 34520 2700 34530 2760
rect 34376 2698 34530 2700
rect 34320 2690 34530 2698
rect 33320 2640 33600 2650
rect 33380 2580 33530 2640
rect 33590 2580 33600 2640
rect 33320 2570 33600 2580
rect 33840 2640 34120 2650
rect 33900 2580 34050 2640
rect 34110 2580 34120 2640
rect 33840 2570 34120 2580
rect 34360 2640 34640 2650
rect 34420 2580 34570 2640
rect 34630 2580 34640 2640
rect 34360 2570 34640 2580
rect 33265 2270 34950 2280
rect 33265 2218 33270 2270
rect 33322 2218 33790 2270
rect 33842 2218 34310 2270
rect 34362 2218 34876 2270
rect 34928 2218 34950 2270
rect 33265 2210 34950 2218
rect 32810 1830 35410 1840
rect 32810 1770 32820 1830
rect 32880 1770 32900 1830
rect 32960 1770 32980 1830
rect 33040 1770 35180 1830
rect 35240 1770 35260 1830
rect 35320 1770 35340 1830
rect 35400 1770 35410 1830
rect 32810 1750 35410 1770
rect 32810 1690 32820 1750
rect 32880 1690 32900 1750
rect 32960 1690 32980 1750
rect 33040 1690 35180 1750
rect 35240 1690 35260 1750
rect 35320 1690 35340 1750
rect 35400 1690 35410 1750
rect 32810 1670 35410 1690
rect 32810 1610 32820 1670
rect 32880 1610 32900 1670
rect 32960 1610 32980 1670
rect 33040 1610 35180 1670
rect 35240 1610 35260 1670
rect 35320 1610 35340 1670
rect 35400 1610 35410 1670
rect 32810 1600 35410 1610
rect 33310 1560 34920 1570
rect 33310 1500 33320 1560
rect 33380 1500 33840 1560
rect 33900 1500 34360 1560
rect 34420 1500 34850 1560
rect 34910 1500 34920 1560
rect 33310 1490 34920 1500
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
