magic
tech sky130A
magscale 1 2
timestamp 1757210648
<< nwell >>
rect 8567 16457 9091 18625
rect 9347 14887 9871 18631
rect 10127 16111 10983 18633
rect 15447 16111 16303 18633
rect 16557 15777 17081 18631
rect 17347 16457 17871 18625
rect 11367 14117 15189 14641
rect 10400 11180 13130 11460
rect 13430 11180 16160 11460
rect 11500 9620 15060 10300
rect 15360 9820 16130 10100
rect 11510 9020 13150 9300
rect 13410 9020 15050 9300
<< pwell >>
rect 13240 18810 13320 19090
rect 11250 18657 12590 18810
rect 11250 17623 11403 18657
rect 12437 17623 12590 18657
rect 11250 17470 12590 17623
rect 12610 18657 13950 18810
rect 12610 17623 12763 18657
rect 13797 17623 13950 18657
rect 12610 17470 13950 17623
rect 13970 18657 15310 18810
rect 13970 17623 14123 18657
rect 15157 17623 15310 18657
rect 13970 17470 15310 17623
rect 11250 17297 12590 17450
rect 11250 16263 11403 17297
rect 12437 16263 12590 17297
rect 11250 16110 12590 16263
rect 12610 17297 13950 17450
rect 12610 16263 12763 17297
rect 13797 16263 13950 17297
rect 12610 16110 13950 16263
rect 13970 17297 15310 17450
rect 13970 16263 14123 17297
rect 15157 16263 15310 17297
rect 13970 16110 15310 16263
rect 11250 15937 12590 16090
rect 11250 14903 11403 15937
rect 12437 14903 12590 15937
rect 11250 14750 12590 14903
rect 12610 15937 13950 16090
rect 12610 14903 12763 15937
rect 13797 14903 13950 15937
rect 12610 14750 13950 14903
rect 13970 15937 15310 16090
rect 13970 14903 14123 15937
rect 15157 14903 15310 15937
rect 13970 14750 15310 14903
<< nbase >>
rect 11403 17623 12437 18657
rect 12763 17623 13797 18657
rect 14123 17623 15157 18657
rect 11403 16263 12437 17297
rect 12763 16263 13797 17297
rect 14123 16263 15157 17297
rect 11403 14903 12437 15937
rect 12763 14903 13797 15937
rect 14123 14903 15157 15937
<< nmos >>
rect 11240 13680 13240 13880
rect 13320 13680 15320 13880
rect 10820 12770 11820 13270
rect 12060 12770 13060 13270
rect 13500 12770 14500 13270
rect 14740 12770 15740 13270
rect 11440 12160 11480 12260
rect 11560 12160 11600 12260
rect 11680 12160 11720 12260
rect 11800 12160 11840 12260
rect 11920 12160 11960 12260
rect 12040 12160 12080 12260
rect 12160 12160 12200 12260
rect 12280 12160 12320 12260
rect 12400 12160 12440 12260
rect 12520 12160 12560 12260
rect 14000 12160 14040 12260
rect 14120 12160 14160 12260
rect 14240 12160 14280 12260
rect 14360 12160 14400 12260
rect 14480 12160 14520 12260
rect 14600 12160 14640 12260
rect 14720 12160 14760 12260
rect 14840 12160 14880 12260
rect 14960 12160 15000 12260
rect 15080 12160 15120 12260
<< pmos >>
rect 10600 11220 10640 11420
rect 10720 11220 10760 11420
rect 10840 11220 10880 11420
rect 10960 11220 11000 11420
rect 11080 11220 11120 11420
rect 11200 11220 11240 11420
rect 11320 11220 11360 11420
rect 11440 11220 11480 11420
rect 11560 11220 11600 11420
rect 11680 11220 11720 11420
rect 11800 11220 11840 11420
rect 11920 11220 11960 11420
rect 12040 11220 12080 11420
rect 12160 11220 12200 11420
rect 12280 11220 12320 11420
rect 12400 11220 12440 11420
rect 12520 11220 12560 11420
rect 12640 11220 12680 11420
rect 12760 11220 12800 11420
rect 12880 11220 12920 11420
rect 13640 11220 13680 11420
rect 13760 11220 13800 11420
rect 13880 11220 13920 11420
rect 14000 11220 14040 11420
rect 14120 11220 14160 11420
rect 14240 11220 14280 11420
rect 14360 11220 14400 11420
rect 14480 11220 14520 11420
rect 14600 11220 14640 11420
rect 14720 11220 14760 11420
rect 14840 11220 14880 11420
rect 14960 11220 15000 11420
rect 15080 11220 15120 11420
rect 15200 11220 15240 11420
rect 15320 11220 15360 11420
rect 15440 11220 15480 11420
rect 15560 11220 15600 11420
rect 15680 11220 15720 11420
rect 15800 11220 15840 11420
rect 15920 11220 15960 11420
rect 11700 9660 11800 10260
rect 11880 9660 11980 10260
rect 12060 9660 12160 10260
rect 12240 9660 12340 10260
rect 12420 9660 12520 10260
rect 12600 9660 12700 10260
rect 12780 9660 12880 10260
rect 12960 9660 13060 10260
rect 13140 9660 13240 10260
rect 13320 9660 13420 10260
rect 13500 9660 13600 10260
rect 13680 9660 13780 10260
rect 13860 9660 13960 10260
rect 14040 9660 14140 10260
rect 14220 9660 14320 10260
rect 14400 9660 14500 10260
rect 14580 9660 14680 10260
rect 14760 9660 14860 10260
rect 15570 9860 15600 10060
rect 15680 9860 15710 10060
rect 15790 9860 15820 10060
rect 15900 9860 15930 10060
rect 11710 9060 11740 9260
rect 11820 9060 11850 9260
rect 11930 9060 11960 9260
rect 12040 9060 12070 9260
rect 12150 9060 12180 9260
rect 12260 9060 12290 9260
rect 12370 9060 12400 9260
rect 12480 9060 12510 9260
rect 12590 9060 12620 9260
rect 12700 9060 12730 9260
rect 12810 9060 12840 9260
rect 12920 9060 12950 9260
rect 13610 9060 13640 9260
rect 13720 9060 13750 9260
rect 13830 9060 13860 9260
rect 13940 9060 13970 9260
rect 14050 9060 14080 9260
rect 14160 9060 14190 9260
rect 14270 9060 14300 9260
rect 14380 9060 14410 9260
rect 14490 9060 14520 9260
rect 14600 9060 14630 9260
rect 14710 9060 14740 9260
rect 14820 9060 14850 9260
<< ndiff >>
rect 11160 13850 11240 13880
rect 11160 13810 11180 13850
rect 11220 13810 11240 13850
rect 11160 13750 11240 13810
rect 11160 13710 11180 13750
rect 11220 13710 11240 13750
rect 11160 13680 11240 13710
rect 13240 13850 13320 13880
rect 13240 13810 13260 13850
rect 13300 13810 13320 13850
rect 13240 13750 13320 13810
rect 13240 13710 13260 13750
rect 13300 13710 13320 13750
rect 13240 13680 13320 13710
rect 15320 13850 15400 13880
rect 15320 13810 15340 13850
rect 15380 13810 15400 13850
rect 15320 13750 15400 13810
rect 15320 13710 15340 13750
rect 15380 13710 15400 13750
rect 15320 13680 15400 13710
rect 10740 13240 10820 13270
rect 10740 13200 10760 13240
rect 10800 13200 10820 13240
rect 10740 13140 10820 13200
rect 10740 13100 10760 13140
rect 10800 13100 10820 13140
rect 10740 13040 10820 13100
rect 10740 13000 10760 13040
rect 10800 13000 10820 13040
rect 10740 12940 10820 13000
rect 10740 12900 10760 12940
rect 10800 12900 10820 12940
rect 10740 12840 10820 12900
rect 10740 12800 10760 12840
rect 10800 12800 10820 12840
rect 10740 12770 10820 12800
rect 11820 13240 11900 13270
rect 11980 13240 12060 13270
rect 11820 13200 11840 13240
rect 11880 13200 11900 13240
rect 11980 13200 12000 13240
rect 12040 13200 12060 13240
rect 11820 13140 11900 13200
rect 11980 13140 12060 13200
rect 11820 13100 11840 13140
rect 11880 13100 11900 13140
rect 11980 13100 12000 13140
rect 12040 13100 12060 13140
rect 11820 13040 11900 13100
rect 11980 13040 12060 13100
rect 11820 13000 11840 13040
rect 11880 13000 11900 13040
rect 11980 13000 12000 13040
rect 12040 13000 12060 13040
rect 11820 12940 11900 13000
rect 11980 12940 12060 13000
rect 11820 12900 11840 12940
rect 11880 12900 11900 12940
rect 11980 12900 12000 12940
rect 12040 12900 12060 12940
rect 11820 12840 11900 12900
rect 11980 12840 12060 12900
rect 11820 12800 11840 12840
rect 11880 12800 11900 12840
rect 11980 12800 12000 12840
rect 12040 12800 12060 12840
rect 11820 12770 11900 12800
rect 11980 12770 12060 12800
rect 13060 13240 13140 13270
rect 13060 13200 13080 13240
rect 13120 13200 13140 13240
rect 13060 13140 13140 13200
rect 13060 13100 13080 13140
rect 13120 13100 13140 13140
rect 13060 13040 13140 13100
rect 13060 13000 13080 13040
rect 13120 13000 13140 13040
rect 13060 12940 13140 13000
rect 13060 12900 13080 12940
rect 13120 12900 13140 12940
rect 13060 12840 13140 12900
rect 13060 12800 13080 12840
rect 13120 12800 13140 12840
rect 13060 12770 13140 12800
rect 13420 13240 13500 13270
rect 13420 13200 13440 13240
rect 13480 13200 13500 13240
rect 13420 13140 13500 13200
rect 13420 13100 13440 13140
rect 13480 13100 13500 13140
rect 13420 13040 13500 13100
rect 13420 13000 13440 13040
rect 13480 13000 13500 13040
rect 13420 12940 13500 13000
rect 13420 12900 13440 12940
rect 13480 12900 13500 12940
rect 13420 12840 13500 12900
rect 13420 12800 13440 12840
rect 13480 12800 13500 12840
rect 13420 12770 13500 12800
rect 14500 13240 14580 13270
rect 14660 13240 14740 13270
rect 14500 13200 14520 13240
rect 14560 13200 14580 13240
rect 14660 13200 14680 13240
rect 14720 13200 14740 13240
rect 14500 13140 14580 13200
rect 14660 13140 14740 13200
rect 14500 13100 14520 13140
rect 14560 13100 14580 13140
rect 14660 13100 14680 13140
rect 14720 13100 14740 13140
rect 14500 13040 14580 13100
rect 14660 13040 14740 13100
rect 14500 13000 14520 13040
rect 14560 13000 14580 13040
rect 14660 13000 14680 13040
rect 14720 13000 14740 13040
rect 14500 12940 14580 13000
rect 14660 12940 14740 13000
rect 14500 12900 14520 12940
rect 14560 12900 14580 12940
rect 14660 12900 14680 12940
rect 14720 12900 14740 12940
rect 14500 12840 14580 12900
rect 14660 12840 14740 12900
rect 14500 12800 14520 12840
rect 14560 12800 14580 12840
rect 14660 12800 14680 12840
rect 14720 12800 14740 12840
rect 14500 12770 14580 12800
rect 14660 12770 14740 12800
rect 15740 13240 15820 13270
rect 15740 13200 15760 13240
rect 15800 13200 15820 13240
rect 15740 13140 15820 13200
rect 15740 13100 15760 13140
rect 15800 13100 15820 13140
rect 15740 13040 15820 13100
rect 15740 13000 15760 13040
rect 15800 13000 15820 13040
rect 15740 12940 15820 13000
rect 15740 12900 15760 12940
rect 15800 12900 15820 12940
rect 15740 12840 15820 12900
rect 15740 12800 15760 12840
rect 15800 12800 15820 12840
rect 15740 12770 15820 12800
rect 11360 12230 11440 12260
rect 11360 12190 11380 12230
rect 11420 12190 11440 12230
rect 11360 12160 11440 12190
rect 11480 12230 11560 12260
rect 11480 12190 11500 12230
rect 11540 12190 11560 12230
rect 11480 12160 11560 12190
rect 11600 12230 11680 12260
rect 11600 12190 11620 12230
rect 11660 12190 11680 12230
rect 11600 12160 11680 12190
rect 11720 12230 11800 12260
rect 11720 12190 11740 12230
rect 11780 12190 11800 12230
rect 11720 12160 11800 12190
rect 11840 12230 11920 12260
rect 11840 12190 11860 12230
rect 11900 12190 11920 12230
rect 11840 12160 11920 12190
rect 11960 12230 12040 12260
rect 11960 12190 11980 12230
rect 12020 12190 12040 12230
rect 11960 12160 12040 12190
rect 12080 12230 12160 12260
rect 12080 12190 12100 12230
rect 12140 12190 12160 12230
rect 12080 12160 12160 12190
rect 12200 12230 12280 12260
rect 12200 12190 12220 12230
rect 12260 12190 12280 12230
rect 12200 12160 12280 12190
rect 12320 12230 12400 12260
rect 12320 12190 12340 12230
rect 12380 12190 12400 12230
rect 12320 12160 12400 12190
rect 12440 12230 12520 12260
rect 12440 12190 12460 12230
rect 12500 12190 12520 12230
rect 12440 12160 12520 12190
rect 12560 12230 12640 12260
rect 12560 12190 12580 12230
rect 12620 12190 12640 12230
rect 12560 12160 12640 12190
rect 13920 12230 14000 12260
rect 13920 12190 13940 12230
rect 13980 12190 14000 12230
rect 13920 12160 14000 12190
rect 14040 12230 14120 12260
rect 14040 12190 14060 12230
rect 14100 12190 14120 12230
rect 14040 12160 14120 12190
rect 14160 12230 14240 12260
rect 14160 12190 14180 12230
rect 14220 12190 14240 12230
rect 14160 12160 14240 12190
rect 14280 12230 14360 12260
rect 14280 12190 14300 12230
rect 14340 12190 14360 12230
rect 14280 12160 14360 12190
rect 14400 12230 14480 12260
rect 14400 12190 14420 12230
rect 14460 12190 14480 12230
rect 14400 12160 14480 12190
rect 14520 12230 14600 12260
rect 14520 12190 14540 12230
rect 14580 12190 14600 12230
rect 14520 12160 14600 12190
rect 14640 12230 14720 12260
rect 14640 12190 14660 12230
rect 14700 12190 14720 12230
rect 14640 12160 14720 12190
rect 14760 12230 14840 12260
rect 14760 12190 14780 12230
rect 14820 12190 14840 12230
rect 14760 12160 14840 12190
rect 14880 12230 14960 12260
rect 14880 12190 14900 12230
rect 14940 12190 14960 12230
rect 14880 12160 14960 12190
rect 15000 12230 15080 12260
rect 15000 12190 15020 12230
rect 15060 12190 15080 12230
rect 15000 12160 15080 12190
rect 15120 12230 15200 12260
rect 15120 12190 15140 12230
rect 15180 12190 15200 12230
rect 15120 12160 15200 12190
<< pdiff >>
rect 11580 18426 12260 18480
rect 11580 18392 11632 18426
rect 11666 18392 11722 18426
rect 11756 18392 11812 18426
rect 11846 18392 11902 18426
rect 11936 18392 11992 18426
rect 12026 18392 12082 18426
rect 12116 18392 12172 18426
rect 12206 18392 12260 18426
rect 11580 18336 12260 18392
rect 11580 18302 11632 18336
rect 11666 18302 11722 18336
rect 11756 18302 11812 18336
rect 11846 18302 11902 18336
rect 11936 18302 11992 18336
rect 12026 18302 12082 18336
rect 12116 18302 12172 18336
rect 12206 18302 12260 18336
rect 11580 18246 12260 18302
rect 11580 18212 11632 18246
rect 11666 18212 11722 18246
rect 11756 18212 11812 18246
rect 11846 18212 11902 18246
rect 11936 18212 11992 18246
rect 12026 18212 12082 18246
rect 12116 18212 12172 18246
rect 12206 18212 12260 18246
rect 11580 18156 12260 18212
rect 11580 18122 11632 18156
rect 11666 18122 11722 18156
rect 11756 18122 11812 18156
rect 11846 18122 11902 18156
rect 11936 18122 11992 18156
rect 12026 18122 12082 18156
rect 12116 18122 12172 18156
rect 12206 18122 12260 18156
rect 11580 18066 12260 18122
rect 11580 18032 11632 18066
rect 11666 18032 11722 18066
rect 11756 18032 11812 18066
rect 11846 18032 11902 18066
rect 11936 18032 11992 18066
rect 12026 18032 12082 18066
rect 12116 18032 12172 18066
rect 12206 18032 12260 18066
rect 11580 17976 12260 18032
rect 11580 17942 11632 17976
rect 11666 17942 11722 17976
rect 11756 17942 11812 17976
rect 11846 17942 11902 17976
rect 11936 17942 11992 17976
rect 12026 17942 12082 17976
rect 12116 17942 12172 17976
rect 12206 17942 12260 17976
rect 11580 17886 12260 17942
rect 11580 17852 11632 17886
rect 11666 17852 11722 17886
rect 11756 17852 11812 17886
rect 11846 17852 11902 17886
rect 11936 17852 11992 17886
rect 12026 17852 12082 17886
rect 12116 17852 12172 17886
rect 12206 17852 12260 17886
rect 11580 17800 12260 17852
rect 12940 18426 13620 18480
rect 12940 18392 12992 18426
rect 13026 18392 13082 18426
rect 13116 18392 13172 18426
rect 13206 18392 13262 18426
rect 13296 18392 13352 18426
rect 13386 18392 13442 18426
rect 13476 18392 13532 18426
rect 13566 18392 13620 18426
rect 12940 18336 13620 18392
rect 12940 18302 12992 18336
rect 13026 18302 13082 18336
rect 13116 18302 13172 18336
rect 13206 18302 13262 18336
rect 13296 18302 13352 18336
rect 13386 18302 13442 18336
rect 13476 18302 13532 18336
rect 13566 18302 13620 18336
rect 12940 18246 13620 18302
rect 12940 18212 12992 18246
rect 13026 18212 13082 18246
rect 13116 18212 13172 18246
rect 13206 18212 13262 18246
rect 13296 18212 13352 18246
rect 13386 18212 13442 18246
rect 13476 18212 13532 18246
rect 13566 18212 13620 18246
rect 12940 18156 13620 18212
rect 12940 18122 12992 18156
rect 13026 18122 13082 18156
rect 13116 18122 13172 18156
rect 13206 18122 13262 18156
rect 13296 18122 13352 18156
rect 13386 18122 13442 18156
rect 13476 18122 13532 18156
rect 13566 18122 13620 18156
rect 12940 18066 13620 18122
rect 12940 18032 12992 18066
rect 13026 18032 13082 18066
rect 13116 18032 13172 18066
rect 13206 18032 13262 18066
rect 13296 18032 13352 18066
rect 13386 18032 13442 18066
rect 13476 18032 13532 18066
rect 13566 18032 13620 18066
rect 12940 17976 13620 18032
rect 12940 17942 12992 17976
rect 13026 17942 13082 17976
rect 13116 17942 13172 17976
rect 13206 17942 13262 17976
rect 13296 17942 13352 17976
rect 13386 17942 13442 17976
rect 13476 17942 13532 17976
rect 13566 17942 13620 17976
rect 12940 17886 13620 17942
rect 12940 17852 12992 17886
rect 13026 17852 13082 17886
rect 13116 17852 13172 17886
rect 13206 17852 13262 17886
rect 13296 17852 13352 17886
rect 13386 17852 13442 17886
rect 13476 17852 13532 17886
rect 13566 17852 13620 17886
rect 12940 17800 13620 17852
rect 14300 18426 14980 18480
rect 14300 18392 14352 18426
rect 14386 18392 14442 18426
rect 14476 18392 14532 18426
rect 14566 18392 14622 18426
rect 14656 18392 14712 18426
rect 14746 18392 14802 18426
rect 14836 18392 14892 18426
rect 14926 18392 14980 18426
rect 14300 18336 14980 18392
rect 14300 18302 14352 18336
rect 14386 18302 14442 18336
rect 14476 18302 14532 18336
rect 14566 18302 14622 18336
rect 14656 18302 14712 18336
rect 14746 18302 14802 18336
rect 14836 18302 14892 18336
rect 14926 18302 14980 18336
rect 14300 18246 14980 18302
rect 14300 18212 14352 18246
rect 14386 18212 14442 18246
rect 14476 18212 14532 18246
rect 14566 18212 14622 18246
rect 14656 18212 14712 18246
rect 14746 18212 14802 18246
rect 14836 18212 14892 18246
rect 14926 18212 14980 18246
rect 14300 18156 14980 18212
rect 14300 18122 14352 18156
rect 14386 18122 14442 18156
rect 14476 18122 14532 18156
rect 14566 18122 14622 18156
rect 14656 18122 14712 18156
rect 14746 18122 14802 18156
rect 14836 18122 14892 18156
rect 14926 18122 14980 18156
rect 14300 18066 14980 18122
rect 14300 18032 14352 18066
rect 14386 18032 14442 18066
rect 14476 18032 14532 18066
rect 14566 18032 14622 18066
rect 14656 18032 14712 18066
rect 14746 18032 14802 18066
rect 14836 18032 14892 18066
rect 14926 18032 14980 18066
rect 14300 17976 14980 18032
rect 14300 17942 14352 17976
rect 14386 17942 14442 17976
rect 14476 17942 14532 17976
rect 14566 17942 14622 17976
rect 14656 17942 14712 17976
rect 14746 17942 14802 17976
rect 14836 17942 14892 17976
rect 14926 17942 14980 17976
rect 14300 17886 14980 17942
rect 14300 17852 14352 17886
rect 14386 17852 14442 17886
rect 14476 17852 14532 17886
rect 14566 17852 14622 17886
rect 14656 17852 14712 17886
rect 14746 17852 14802 17886
rect 14836 17852 14892 17886
rect 14926 17852 14980 17886
rect 14300 17800 14980 17852
rect 11580 17066 12260 17120
rect 11580 17032 11632 17066
rect 11666 17032 11722 17066
rect 11756 17032 11812 17066
rect 11846 17032 11902 17066
rect 11936 17032 11992 17066
rect 12026 17032 12082 17066
rect 12116 17032 12172 17066
rect 12206 17032 12260 17066
rect 11580 16976 12260 17032
rect 11580 16942 11632 16976
rect 11666 16942 11722 16976
rect 11756 16942 11812 16976
rect 11846 16942 11902 16976
rect 11936 16942 11992 16976
rect 12026 16942 12082 16976
rect 12116 16942 12172 16976
rect 12206 16942 12260 16976
rect 11580 16886 12260 16942
rect 11580 16852 11632 16886
rect 11666 16852 11722 16886
rect 11756 16852 11812 16886
rect 11846 16852 11902 16886
rect 11936 16852 11992 16886
rect 12026 16852 12082 16886
rect 12116 16852 12172 16886
rect 12206 16852 12260 16886
rect 11580 16796 12260 16852
rect 11580 16762 11632 16796
rect 11666 16762 11722 16796
rect 11756 16762 11812 16796
rect 11846 16762 11902 16796
rect 11936 16762 11992 16796
rect 12026 16762 12082 16796
rect 12116 16762 12172 16796
rect 12206 16762 12260 16796
rect 11580 16706 12260 16762
rect 11580 16672 11632 16706
rect 11666 16672 11722 16706
rect 11756 16672 11812 16706
rect 11846 16672 11902 16706
rect 11936 16672 11992 16706
rect 12026 16672 12082 16706
rect 12116 16672 12172 16706
rect 12206 16672 12260 16706
rect 11580 16616 12260 16672
rect 11580 16582 11632 16616
rect 11666 16582 11722 16616
rect 11756 16582 11812 16616
rect 11846 16582 11902 16616
rect 11936 16582 11992 16616
rect 12026 16582 12082 16616
rect 12116 16582 12172 16616
rect 12206 16582 12260 16616
rect 11580 16526 12260 16582
rect 11580 16492 11632 16526
rect 11666 16492 11722 16526
rect 11756 16492 11812 16526
rect 11846 16492 11902 16526
rect 11936 16492 11992 16526
rect 12026 16492 12082 16526
rect 12116 16492 12172 16526
rect 12206 16492 12260 16526
rect 11580 16440 12260 16492
rect 12940 17066 13620 17120
rect 12940 17032 12992 17066
rect 13026 17032 13082 17066
rect 13116 17032 13172 17066
rect 13206 17032 13262 17066
rect 13296 17032 13352 17066
rect 13386 17032 13442 17066
rect 13476 17032 13532 17066
rect 13566 17032 13620 17066
rect 12940 16976 13620 17032
rect 12940 16942 12992 16976
rect 13026 16942 13082 16976
rect 13116 16942 13172 16976
rect 13206 16942 13262 16976
rect 13296 16942 13352 16976
rect 13386 16942 13442 16976
rect 13476 16942 13532 16976
rect 13566 16942 13620 16976
rect 12940 16886 13620 16942
rect 12940 16852 12992 16886
rect 13026 16852 13082 16886
rect 13116 16852 13172 16886
rect 13206 16852 13262 16886
rect 13296 16852 13352 16886
rect 13386 16852 13442 16886
rect 13476 16852 13532 16886
rect 13566 16852 13620 16886
rect 12940 16796 13620 16852
rect 12940 16762 12992 16796
rect 13026 16762 13082 16796
rect 13116 16762 13172 16796
rect 13206 16762 13262 16796
rect 13296 16762 13352 16796
rect 13386 16762 13442 16796
rect 13476 16762 13532 16796
rect 13566 16762 13620 16796
rect 12940 16706 13620 16762
rect 12940 16672 12992 16706
rect 13026 16672 13082 16706
rect 13116 16672 13172 16706
rect 13206 16672 13262 16706
rect 13296 16672 13352 16706
rect 13386 16672 13442 16706
rect 13476 16672 13532 16706
rect 13566 16672 13620 16706
rect 12940 16616 13620 16672
rect 12940 16582 12992 16616
rect 13026 16582 13082 16616
rect 13116 16582 13172 16616
rect 13206 16582 13262 16616
rect 13296 16582 13352 16616
rect 13386 16582 13442 16616
rect 13476 16582 13532 16616
rect 13566 16582 13620 16616
rect 12940 16526 13620 16582
rect 12940 16492 12992 16526
rect 13026 16492 13082 16526
rect 13116 16492 13172 16526
rect 13206 16492 13262 16526
rect 13296 16492 13352 16526
rect 13386 16492 13442 16526
rect 13476 16492 13532 16526
rect 13566 16492 13620 16526
rect 12940 16440 13620 16492
rect 14300 17066 14980 17120
rect 14300 17032 14352 17066
rect 14386 17032 14442 17066
rect 14476 17032 14532 17066
rect 14566 17032 14622 17066
rect 14656 17032 14712 17066
rect 14746 17032 14802 17066
rect 14836 17032 14892 17066
rect 14926 17032 14980 17066
rect 14300 16976 14980 17032
rect 14300 16942 14352 16976
rect 14386 16942 14442 16976
rect 14476 16942 14532 16976
rect 14566 16942 14622 16976
rect 14656 16942 14712 16976
rect 14746 16942 14802 16976
rect 14836 16942 14892 16976
rect 14926 16942 14980 16976
rect 14300 16886 14980 16942
rect 14300 16852 14352 16886
rect 14386 16852 14442 16886
rect 14476 16852 14532 16886
rect 14566 16852 14622 16886
rect 14656 16852 14712 16886
rect 14746 16852 14802 16886
rect 14836 16852 14892 16886
rect 14926 16852 14980 16886
rect 14300 16796 14980 16852
rect 14300 16762 14352 16796
rect 14386 16762 14442 16796
rect 14476 16762 14532 16796
rect 14566 16762 14622 16796
rect 14656 16762 14712 16796
rect 14746 16762 14802 16796
rect 14836 16762 14892 16796
rect 14926 16762 14980 16796
rect 14300 16706 14980 16762
rect 14300 16672 14352 16706
rect 14386 16672 14442 16706
rect 14476 16672 14532 16706
rect 14566 16672 14622 16706
rect 14656 16672 14712 16706
rect 14746 16672 14802 16706
rect 14836 16672 14892 16706
rect 14926 16672 14980 16706
rect 14300 16616 14980 16672
rect 14300 16582 14352 16616
rect 14386 16582 14442 16616
rect 14476 16582 14532 16616
rect 14566 16582 14622 16616
rect 14656 16582 14712 16616
rect 14746 16582 14802 16616
rect 14836 16582 14892 16616
rect 14926 16582 14980 16616
rect 14300 16526 14980 16582
rect 14300 16492 14352 16526
rect 14386 16492 14442 16526
rect 14476 16492 14532 16526
rect 14566 16492 14622 16526
rect 14656 16492 14712 16526
rect 14746 16492 14802 16526
rect 14836 16492 14892 16526
rect 14926 16492 14980 16526
rect 14300 16440 14980 16492
rect 11580 15706 12260 15760
rect 11580 15672 11632 15706
rect 11666 15672 11722 15706
rect 11756 15672 11812 15706
rect 11846 15672 11902 15706
rect 11936 15672 11992 15706
rect 12026 15672 12082 15706
rect 12116 15672 12172 15706
rect 12206 15672 12260 15706
rect 11580 15616 12260 15672
rect 11580 15582 11632 15616
rect 11666 15582 11722 15616
rect 11756 15582 11812 15616
rect 11846 15582 11902 15616
rect 11936 15582 11992 15616
rect 12026 15582 12082 15616
rect 12116 15582 12172 15616
rect 12206 15582 12260 15616
rect 11580 15526 12260 15582
rect 11580 15492 11632 15526
rect 11666 15492 11722 15526
rect 11756 15492 11812 15526
rect 11846 15492 11902 15526
rect 11936 15492 11992 15526
rect 12026 15492 12082 15526
rect 12116 15492 12172 15526
rect 12206 15492 12260 15526
rect 11580 15436 12260 15492
rect 11580 15402 11632 15436
rect 11666 15402 11722 15436
rect 11756 15402 11812 15436
rect 11846 15402 11902 15436
rect 11936 15402 11992 15436
rect 12026 15402 12082 15436
rect 12116 15402 12172 15436
rect 12206 15402 12260 15436
rect 11580 15346 12260 15402
rect 11580 15312 11632 15346
rect 11666 15312 11722 15346
rect 11756 15312 11812 15346
rect 11846 15312 11902 15346
rect 11936 15312 11992 15346
rect 12026 15312 12082 15346
rect 12116 15312 12172 15346
rect 12206 15312 12260 15346
rect 11580 15256 12260 15312
rect 11580 15222 11632 15256
rect 11666 15222 11722 15256
rect 11756 15222 11812 15256
rect 11846 15222 11902 15256
rect 11936 15222 11992 15256
rect 12026 15222 12082 15256
rect 12116 15222 12172 15256
rect 12206 15222 12260 15256
rect 11580 15166 12260 15222
rect 11580 15132 11632 15166
rect 11666 15132 11722 15166
rect 11756 15132 11812 15166
rect 11846 15132 11902 15166
rect 11936 15132 11992 15166
rect 12026 15132 12082 15166
rect 12116 15132 12172 15166
rect 12206 15132 12260 15166
rect 11580 15080 12260 15132
rect 12940 15706 13620 15760
rect 12940 15672 12992 15706
rect 13026 15672 13082 15706
rect 13116 15672 13172 15706
rect 13206 15672 13262 15706
rect 13296 15672 13352 15706
rect 13386 15672 13442 15706
rect 13476 15672 13532 15706
rect 13566 15672 13620 15706
rect 12940 15616 13620 15672
rect 12940 15582 12992 15616
rect 13026 15582 13082 15616
rect 13116 15582 13172 15616
rect 13206 15582 13262 15616
rect 13296 15582 13352 15616
rect 13386 15582 13442 15616
rect 13476 15582 13532 15616
rect 13566 15582 13620 15616
rect 12940 15526 13620 15582
rect 12940 15492 12992 15526
rect 13026 15492 13082 15526
rect 13116 15492 13172 15526
rect 13206 15492 13262 15526
rect 13296 15492 13352 15526
rect 13386 15492 13442 15526
rect 13476 15492 13532 15526
rect 13566 15492 13620 15526
rect 12940 15436 13620 15492
rect 12940 15402 12992 15436
rect 13026 15402 13082 15436
rect 13116 15402 13172 15436
rect 13206 15402 13262 15436
rect 13296 15402 13352 15436
rect 13386 15402 13442 15436
rect 13476 15402 13532 15436
rect 13566 15402 13620 15436
rect 12940 15346 13620 15402
rect 12940 15312 12992 15346
rect 13026 15312 13082 15346
rect 13116 15312 13172 15346
rect 13206 15312 13262 15346
rect 13296 15312 13352 15346
rect 13386 15312 13442 15346
rect 13476 15312 13532 15346
rect 13566 15312 13620 15346
rect 12940 15256 13620 15312
rect 12940 15222 12992 15256
rect 13026 15222 13082 15256
rect 13116 15222 13172 15256
rect 13206 15222 13262 15256
rect 13296 15222 13352 15256
rect 13386 15222 13442 15256
rect 13476 15222 13532 15256
rect 13566 15222 13620 15256
rect 12940 15166 13620 15222
rect 12940 15132 12992 15166
rect 13026 15132 13082 15166
rect 13116 15132 13172 15166
rect 13206 15132 13262 15166
rect 13296 15132 13352 15166
rect 13386 15132 13442 15166
rect 13476 15132 13532 15166
rect 13566 15132 13620 15166
rect 12940 15080 13620 15132
rect 14300 15706 14980 15760
rect 14300 15672 14352 15706
rect 14386 15672 14442 15706
rect 14476 15672 14532 15706
rect 14566 15672 14622 15706
rect 14656 15672 14712 15706
rect 14746 15672 14802 15706
rect 14836 15672 14892 15706
rect 14926 15672 14980 15706
rect 14300 15616 14980 15672
rect 14300 15582 14352 15616
rect 14386 15582 14442 15616
rect 14476 15582 14532 15616
rect 14566 15582 14622 15616
rect 14656 15582 14712 15616
rect 14746 15582 14802 15616
rect 14836 15582 14892 15616
rect 14926 15582 14980 15616
rect 14300 15526 14980 15582
rect 14300 15492 14352 15526
rect 14386 15492 14442 15526
rect 14476 15492 14532 15526
rect 14566 15492 14622 15526
rect 14656 15492 14712 15526
rect 14746 15492 14802 15526
rect 14836 15492 14892 15526
rect 14926 15492 14980 15526
rect 14300 15436 14980 15492
rect 14300 15402 14352 15436
rect 14386 15402 14442 15436
rect 14476 15402 14532 15436
rect 14566 15402 14622 15436
rect 14656 15402 14712 15436
rect 14746 15402 14802 15436
rect 14836 15402 14892 15436
rect 14926 15402 14980 15436
rect 14300 15346 14980 15402
rect 14300 15312 14352 15346
rect 14386 15312 14442 15346
rect 14476 15312 14532 15346
rect 14566 15312 14622 15346
rect 14656 15312 14712 15346
rect 14746 15312 14802 15346
rect 14836 15312 14892 15346
rect 14926 15312 14980 15346
rect 14300 15256 14980 15312
rect 14300 15222 14352 15256
rect 14386 15222 14442 15256
rect 14476 15222 14532 15256
rect 14566 15222 14622 15256
rect 14656 15222 14712 15256
rect 14746 15222 14802 15256
rect 14836 15222 14892 15256
rect 14926 15222 14980 15256
rect 14300 15166 14980 15222
rect 14300 15132 14352 15166
rect 14386 15132 14442 15166
rect 14476 15132 14532 15166
rect 14566 15132 14622 15166
rect 14656 15132 14712 15166
rect 14746 15132 14802 15166
rect 14836 15132 14892 15166
rect 14926 15132 14980 15166
rect 14300 15080 14980 15132
rect 10520 11390 10600 11420
rect 10520 11350 10540 11390
rect 10580 11350 10600 11390
rect 10520 11290 10600 11350
rect 10520 11250 10540 11290
rect 10580 11250 10600 11290
rect 10520 11220 10600 11250
rect 10640 11390 10720 11420
rect 10640 11350 10660 11390
rect 10700 11350 10720 11390
rect 10640 11290 10720 11350
rect 10640 11250 10660 11290
rect 10700 11250 10720 11290
rect 10640 11220 10720 11250
rect 10760 11390 10840 11420
rect 10760 11350 10780 11390
rect 10820 11350 10840 11390
rect 10760 11290 10840 11350
rect 10760 11250 10780 11290
rect 10820 11250 10840 11290
rect 10760 11220 10840 11250
rect 10880 11390 10960 11420
rect 10880 11350 10900 11390
rect 10940 11350 10960 11390
rect 10880 11290 10960 11350
rect 10880 11250 10900 11290
rect 10940 11250 10960 11290
rect 10880 11220 10960 11250
rect 11000 11390 11080 11420
rect 11000 11350 11020 11390
rect 11060 11350 11080 11390
rect 11000 11290 11080 11350
rect 11000 11250 11020 11290
rect 11060 11250 11080 11290
rect 11000 11220 11080 11250
rect 11120 11390 11200 11420
rect 11120 11350 11140 11390
rect 11180 11350 11200 11390
rect 11120 11290 11200 11350
rect 11120 11250 11140 11290
rect 11180 11250 11200 11290
rect 11120 11220 11200 11250
rect 11240 11390 11320 11420
rect 11240 11350 11260 11390
rect 11300 11350 11320 11390
rect 11240 11290 11320 11350
rect 11240 11250 11260 11290
rect 11300 11250 11320 11290
rect 11240 11220 11320 11250
rect 11360 11390 11440 11420
rect 11360 11350 11380 11390
rect 11420 11350 11440 11390
rect 11360 11290 11440 11350
rect 11360 11250 11380 11290
rect 11420 11250 11440 11290
rect 11360 11220 11440 11250
rect 11480 11390 11560 11420
rect 11480 11350 11500 11390
rect 11540 11350 11560 11390
rect 11480 11290 11560 11350
rect 11480 11250 11500 11290
rect 11540 11250 11560 11290
rect 11480 11220 11560 11250
rect 11600 11390 11680 11420
rect 11600 11350 11620 11390
rect 11660 11350 11680 11390
rect 11600 11290 11680 11350
rect 11600 11250 11620 11290
rect 11660 11250 11680 11290
rect 11600 11220 11680 11250
rect 11720 11390 11800 11420
rect 11720 11350 11740 11390
rect 11780 11350 11800 11390
rect 11720 11290 11800 11350
rect 11720 11250 11740 11290
rect 11780 11250 11800 11290
rect 11720 11220 11800 11250
rect 11840 11390 11920 11420
rect 11840 11350 11860 11390
rect 11900 11350 11920 11390
rect 11840 11290 11920 11350
rect 11840 11250 11860 11290
rect 11900 11250 11920 11290
rect 11840 11220 11920 11250
rect 11960 11390 12040 11420
rect 11960 11350 11980 11390
rect 12020 11350 12040 11390
rect 11960 11290 12040 11350
rect 11960 11250 11980 11290
rect 12020 11250 12040 11290
rect 11960 11220 12040 11250
rect 12080 11390 12160 11420
rect 12080 11350 12100 11390
rect 12140 11350 12160 11390
rect 12080 11290 12160 11350
rect 12080 11250 12100 11290
rect 12140 11250 12160 11290
rect 12080 11220 12160 11250
rect 12200 11390 12280 11420
rect 12200 11350 12220 11390
rect 12260 11350 12280 11390
rect 12200 11290 12280 11350
rect 12200 11250 12220 11290
rect 12260 11250 12280 11290
rect 12200 11220 12280 11250
rect 12320 11390 12400 11420
rect 12320 11350 12340 11390
rect 12380 11350 12400 11390
rect 12320 11290 12400 11350
rect 12320 11250 12340 11290
rect 12380 11250 12400 11290
rect 12320 11220 12400 11250
rect 12440 11390 12520 11420
rect 12440 11350 12460 11390
rect 12500 11350 12520 11390
rect 12440 11290 12520 11350
rect 12440 11250 12460 11290
rect 12500 11250 12520 11290
rect 12440 11220 12520 11250
rect 12560 11390 12640 11420
rect 12560 11350 12580 11390
rect 12620 11350 12640 11390
rect 12560 11290 12640 11350
rect 12560 11250 12580 11290
rect 12620 11250 12640 11290
rect 12560 11220 12640 11250
rect 12680 11390 12760 11420
rect 12680 11350 12700 11390
rect 12740 11350 12760 11390
rect 12680 11290 12760 11350
rect 12680 11250 12700 11290
rect 12740 11250 12760 11290
rect 12680 11220 12760 11250
rect 12800 11390 12880 11420
rect 12800 11350 12820 11390
rect 12860 11350 12880 11390
rect 12800 11290 12880 11350
rect 12800 11250 12820 11290
rect 12860 11250 12880 11290
rect 12800 11220 12880 11250
rect 12920 11390 13000 11420
rect 12920 11350 12940 11390
rect 12980 11350 13000 11390
rect 12920 11290 13000 11350
rect 12920 11250 12940 11290
rect 12980 11250 13000 11290
rect 12920 11220 13000 11250
rect 13560 11390 13640 11420
rect 13560 11350 13580 11390
rect 13620 11350 13640 11390
rect 13560 11290 13640 11350
rect 13560 11250 13580 11290
rect 13620 11250 13640 11290
rect 13560 11220 13640 11250
rect 13680 11390 13760 11420
rect 13680 11350 13700 11390
rect 13740 11350 13760 11390
rect 13680 11290 13760 11350
rect 13680 11250 13700 11290
rect 13740 11250 13760 11290
rect 13680 11220 13760 11250
rect 13800 11390 13880 11420
rect 13800 11350 13820 11390
rect 13860 11350 13880 11390
rect 13800 11290 13880 11350
rect 13800 11250 13820 11290
rect 13860 11250 13880 11290
rect 13800 11220 13880 11250
rect 13920 11390 14000 11420
rect 13920 11350 13940 11390
rect 13980 11350 14000 11390
rect 13920 11290 14000 11350
rect 13920 11250 13940 11290
rect 13980 11250 14000 11290
rect 13920 11220 14000 11250
rect 14040 11390 14120 11420
rect 14040 11350 14060 11390
rect 14100 11350 14120 11390
rect 14040 11290 14120 11350
rect 14040 11250 14060 11290
rect 14100 11250 14120 11290
rect 14040 11220 14120 11250
rect 14160 11390 14240 11420
rect 14160 11350 14180 11390
rect 14220 11350 14240 11390
rect 14160 11290 14240 11350
rect 14160 11250 14180 11290
rect 14220 11250 14240 11290
rect 14160 11220 14240 11250
rect 14280 11390 14360 11420
rect 14280 11350 14300 11390
rect 14340 11350 14360 11390
rect 14280 11290 14360 11350
rect 14280 11250 14300 11290
rect 14340 11250 14360 11290
rect 14280 11220 14360 11250
rect 14400 11390 14480 11420
rect 14400 11350 14420 11390
rect 14460 11350 14480 11390
rect 14400 11290 14480 11350
rect 14400 11250 14420 11290
rect 14460 11250 14480 11290
rect 14400 11220 14480 11250
rect 14520 11390 14600 11420
rect 14520 11350 14540 11390
rect 14580 11350 14600 11390
rect 14520 11290 14600 11350
rect 14520 11250 14540 11290
rect 14580 11250 14600 11290
rect 14520 11220 14600 11250
rect 14640 11390 14720 11420
rect 14640 11350 14660 11390
rect 14700 11350 14720 11390
rect 14640 11290 14720 11350
rect 14640 11250 14660 11290
rect 14700 11250 14720 11290
rect 14640 11220 14720 11250
rect 14760 11390 14840 11420
rect 14760 11350 14780 11390
rect 14820 11350 14840 11390
rect 14760 11290 14840 11350
rect 14760 11250 14780 11290
rect 14820 11250 14840 11290
rect 14760 11220 14840 11250
rect 14880 11390 14960 11420
rect 14880 11350 14900 11390
rect 14940 11350 14960 11390
rect 14880 11290 14960 11350
rect 14880 11250 14900 11290
rect 14940 11250 14960 11290
rect 14880 11220 14960 11250
rect 15000 11390 15080 11420
rect 15000 11350 15020 11390
rect 15060 11350 15080 11390
rect 15000 11290 15080 11350
rect 15000 11250 15020 11290
rect 15060 11250 15080 11290
rect 15000 11220 15080 11250
rect 15120 11390 15200 11420
rect 15120 11350 15140 11390
rect 15180 11350 15200 11390
rect 15120 11290 15200 11350
rect 15120 11250 15140 11290
rect 15180 11250 15200 11290
rect 15120 11220 15200 11250
rect 15240 11390 15320 11420
rect 15240 11350 15260 11390
rect 15300 11350 15320 11390
rect 15240 11290 15320 11350
rect 15240 11250 15260 11290
rect 15300 11250 15320 11290
rect 15240 11220 15320 11250
rect 15360 11390 15440 11420
rect 15360 11350 15380 11390
rect 15420 11350 15440 11390
rect 15360 11290 15440 11350
rect 15360 11250 15380 11290
rect 15420 11250 15440 11290
rect 15360 11220 15440 11250
rect 15480 11390 15560 11420
rect 15480 11350 15500 11390
rect 15540 11350 15560 11390
rect 15480 11290 15560 11350
rect 15480 11250 15500 11290
rect 15540 11250 15560 11290
rect 15480 11220 15560 11250
rect 15600 11390 15680 11420
rect 15600 11350 15620 11390
rect 15660 11350 15680 11390
rect 15600 11290 15680 11350
rect 15600 11250 15620 11290
rect 15660 11250 15680 11290
rect 15600 11220 15680 11250
rect 15720 11390 15800 11420
rect 15720 11350 15740 11390
rect 15780 11350 15800 11390
rect 15720 11290 15800 11350
rect 15720 11250 15740 11290
rect 15780 11250 15800 11290
rect 15720 11220 15800 11250
rect 15840 11390 15920 11420
rect 15840 11350 15860 11390
rect 15900 11350 15920 11390
rect 15840 11290 15920 11350
rect 15840 11250 15860 11290
rect 15900 11250 15920 11290
rect 15840 11220 15920 11250
rect 15960 11390 16040 11420
rect 15960 11350 15980 11390
rect 16020 11350 16040 11390
rect 15960 11290 16040 11350
rect 15960 11250 15980 11290
rect 16020 11250 16040 11290
rect 15960 11220 16040 11250
rect 11620 10230 11700 10260
rect 11620 10190 11640 10230
rect 11680 10190 11700 10230
rect 11620 10130 11700 10190
rect 11620 10090 11640 10130
rect 11680 10090 11700 10130
rect 11620 10030 11700 10090
rect 11620 9990 11640 10030
rect 11680 9990 11700 10030
rect 11620 9930 11700 9990
rect 11620 9890 11640 9930
rect 11680 9890 11700 9930
rect 11620 9830 11700 9890
rect 11620 9790 11640 9830
rect 11680 9790 11700 9830
rect 11620 9730 11700 9790
rect 11620 9690 11640 9730
rect 11680 9690 11700 9730
rect 11620 9660 11700 9690
rect 11800 10230 11880 10260
rect 11800 10190 11820 10230
rect 11860 10190 11880 10230
rect 11800 10130 11880 10190
rect 11800 10090 11820 10130
rect 11860 10090 11880 10130
rect 11800 10030 11880 10090
rect 11800 9990 11820 10030
rect 11860 9990 11880 10030
rect 11800 9930 11880 9990
rect 11800 9890 11820 9930
rect 11860 9890 11880 9930
rect 11800 9830 11880 9890
rect 11800 9790 11820 9830
rect 11860 9790 11880 9830
rect 11800 9730 11880 9790
rect 11800 9690 11820 9730
rect 11860 9690 11880 9730
rect 11800 9660 11880 9690
rect 11980 10230 12060 10260
rect 11980 10190 12000 10230
rect 12040 10190 12060 10230
rect 11980 10130 12060 10190
rect 11980 10090 12000 10130
rect 12040 10090 12060 10130
rect 11980 10030 12060 10090
rect 11980 9990 12000 10030
rect 12040 9990 12060 10030
rect 11980 9930 12060 9990
rect 11980 9890 12000 9930
rect 12040 9890 12060 9930
rect 11980 9830 12060 9890
rect 11980 9790 12000 9830
rect 12040 9790 12060 9830
rect 11980 9730 12060 9790
rect 11980 9690 12000 9730
rect 12040 9690 12060 9730
rect 11980 9660 12060 9690
rect 12160 10230 12240 10260
rect 12160 10190 12180 10230
rect 12220 10190 12240 10230
rect 12160 10130 12240 10190
rect 12160 10090 12180 10130
rect 12220 10090 12240 10130
rect 12160 10030 12240 10090
rect 12160 9990 12180 10030
rect 12220 9990 12240 10030
rect 12160 9930 12240 9990
rect 12160 9890 12180 9930
rect 12220 9890 12240 9930
rect 12160 9830 12240 9890
rect 12160 9790 12180 9830
rect 12220 9790 12240 9830
rect 12160 9730 12240 9790
rect 12160 9690 12180 9730
rect 12220 9690 12240 9730
rect 12160 9660 12240 9690
rect 12340 10230 12420 10260
rect 12340 10190 12360 10230
rect 12400 10190 12420 10230
rect 12340 10130 12420 10190
rect 12340 10090 12360 10130
rect 12400 10090 12420 10130
rect 12340 10030 12420 10090
rect 12340 9990 12360 10030
rect 12400 9990 12420 10030
rect 12340 9930 12420 9990
rect 12340 9890 12360 9930
rect 12400 9890 12420 9930
rect 12340 9830 12420 9890
rect 12340 9790 12360 9830
rect 12400 9790 12420 9830
rect 12340 9730 12420 9790
rect 12340 9690 12360 9730
rect 12400 9690 12420 9730
rect 12340 9660 12420 9690
rect 12520 10230 12600 10260
rect 12520 10190 12540 10230
rect 12580 10190 12600 10230
rect 12520 10130 12600 10190
rect 12520 10090 12540 10130
rect 12580 10090 12600 10130
rect 12520 10030 12600 10090
rect 12520 9990 12540 10030
rect 12580 9990 12600 10030
rect 12520 9930 12600 9990
rect 12520 9890 12540 9930
rect 12580 9890 12600 9930
rect 12520 9830 12600 9890
rect 12520 9790 12540 9830
rect 12580 9790 12600 9830
rect 12520 9730 12600 9790
rect 12520 9690 12540 9730
rect 12580 9690 12600 9730
rect 12520 9660 12600 9690
rect 12700 10230 12780 10260
rect 12700 10190 12720 10230
rect 12760 10190 12780 10230
rect 12700 10130 12780 10190
rect 12700 10090 12720 10130
rect 12760 10090 12780 10130
rect 12700 10030 12780 10090
rect 12700 9990 12720 10030
rect 12760 9990 12780 10030
rect 12700 9930 12780 9990
rect 12700 9890 12720 9930
rect 12760 9890 12780 9930
rect 12700 9830 12780 9890
rect 12700 9790 12720 9830
rect 12760 9790 12780 9830
rect 12700 9730 12780 9790
rect 12700 9690 12720 9730
rect 12760 9690 12780 9730
rect 12700 9660 12780 9690
rect 12880 10230 12960 10260
rect 12880 10190 12900 10230
rect 12940 10190 12960 10230
rect 12880 10130 12960 10190
rect 12880 10090 12900 10130
rect 12940 10090 12960 10130
rect 12880 10030 12960 10090
rect 12880 9990 12900 10030
rect 12940 9990 12960 10030
rect 12880 9930 12960 9990
rect 12880 9890 12900 9930
rect 12940 9890 12960 9930
rect 12880 9830 12960 9890
rect 12880 9790 12900 9830
rect 12940 9790 12960 9830
rect 12880 9730 12960 9790
rect 12880 9690 12900 9730
rect 12940 9690 12960 9730
rect 12880 9660 12960 9690
rect 13060 10230 13140 10260
rect 13060 10190 13080 10230
rect 13120 10190 13140 10230
rect 13060 10130 13140 10190
rect 13060 10090 13080 10130
rect 13120 10090 13140 10130
rect 13060 10030 13140 10090
rect 13060 9990 13080 10030
rect 13120 9990 13140 10030
rect 13060 9930 13140 9990
rect 13060 9890 13080 9930
rect 13120 9890 13140 9930
rect 13060 9830 13140 9890
rect 13060 9790 13080 9830
rect 13120 9790 13140 9830
rect 13060 9730 13140 9790
rect 13060 9690 13080 9730
rect 13120 9690 13140 9730
rect 13060 9660 13140 9690
rect 13240 10230 13320 10260
rect 13240 10190 13260 10230
rect 13300 10190 13320 10230
rect 13240 10130 13320 10190
rect 13240 10090 13260 10130
rect 13300 10090 13320 10130
rect 13240 10030 13320 10090
rect 13240 9990 13260 10030
rect 13300 9990 13320 10030
rect 13240 9930 13320 9990
rect 13240 9890 13260 9930
rect 13300 9890 13320 9930
rect 13240 9830 13320 9890
rect 13240 9790 13260 9830
rect 13300 9790 13320 9830
rect 13240 9730 13320 9790
rect 13240 9690 13260 9730
rect 13300 9690 13320 9730
rect 13240 9660 13320 9690
rect 13420 10230 13500 10260
rect 13420 10190 13440 10230
rect 13480 10190 13500 10230
rect 13420 10130 13500 10190
rect 13420 10090 13440 10130
rect 13480 10090 13500 10130
rect 13420 10030 13500 10090
rect 13420 9990 13440 10030
rect 13480 9990 13500 10030
rect 13420 9930 13500 9990
rect 13420 9890 13440 9930
rect 13480 9890 13500 9930
rect 13420 9830 13500 9890
rect 13420 9790 13440 9830
rect 13480 9790 13500 9830
rect 13420 9730 13500 9790
rect 13420 9690 13440 9730
rect 13480 9690 13500 9730
rect 13420 9660 13500 9690
rect 13600 10230 13680 10260
rect 13600 10190 13620 10230
rect 13660 10190 13680 10230
rect 13600 10130 13680 10190
rect 13600 10090 13620 10130
rect 13660 10090 13680 10130
rect 13600 10030 13680 10090
rect 13600 9990 13620 10030
rect 13660 9990 13680 10030
rect 13600 9930 13680 9990
rect 13600 9890 13620 9930
rect 13660 9890 13680 9930
rect 13600 9830 13680 9890
rect 13600 9790 13620 9830
rect 13660 9790 13680 9830
rect 13600 9730 13680 9790
rect 13600 9690 13620 9730
rect 13660 9690 13680 9730
rect 13600 9660 13680 9690
rect 13780 10230 13860 10260
rect 13780 10190 13800 10230
rect 13840 10190 13860 10230
rect 13780 10130 13860 10190
rect 13780 10090 13800 10130
rect 13840 10090 13860 10130
rect 13780 10030 13860 10090
rect 13780 9990 13800 10030
rect 13840 9990 13860 10030
rect 13780 9930 13860 9990
rect 13780 9890 13800 9930
rect 13840 9890 13860 9930
rect 13780 9830 13860 9890
rect 13780 9790 13800 9830
rect 13840 9790 13860 9830
rect 13780 9730 13860 9790
rect 13780 9690 13800 9730
rect 13840 9690 13860 9730
rect 13780 9660 13860 9690
rect 13960 10230 14040 10260
rect 13960 10190 13980 10230
rect 14020 10190 14040 10230
rect 13960 10130 14040 10190
rect 13960 10090 13980 10130
rect 14020 10090 14040 10130
rect 13960 10030 14040 10090
rect 13960 9990 13980 10030
rect 14020 9990 14040 10030
rect 13960 9930 14040 9990
rect 13960 9890 13980 9930
rect 14020 9890 14040 9930
rect 13960 9830 14040 9890
rect 13960 9790 13980 9830
rect 14020 9790 14040 9830
rect 13960 9730 14040 9790
rect 13960 9690 13980 9730
rect 14020 9690 14040 9730
rect 13960 9660 14040 9690
rect 14140 10230 14220 10260
rect 14140 10190 14160 10230
rect 14200 10190 14220 10230
rect 14140 10130 14220 10190
rect 14140 10090 14160 10130
rect 14200 10090 14220 10130
rect 14140 10030 14220 10090
rect 14140 9990 14160 10030
rect 14200 9990 14220 10030
rect 14140 9930 14220 9990
rect 14140 9890 14160 9930
rect 14200 9890 14220 9930
rect 14140 9830 14220 9890
rect 14140 9790 14160 9830
rect 14200 9790 14220 9830
rect 14140 9730 14220 9790
rect 14140 9690 14160 9730
rect 14200 9690 14220 9730
rect 14140 9660 14220 9690
rect 14320 10230 14400 10260
rect 14320 10190 14340 10230
rect 14380 10190 14400 10230
rect 14320 10130 14400 10190
rect 14320 10090 14340 10130
rect 14380 10090 14400 10130
rect 14320 10030 14400 10090
rect 14320 9990 14340 10030
rect 14380 9990 14400 10030
rect 14320 9930 14400 9990
rect 14320 9890 14340 9930
rect 14380 9890 14400 9930
rect 14320 9830 14400 9890
rect 14320 9790 14340 9830
rect 14380 9790 14400 9830
rect 14320 9730 14400 9790
rect 14320 9690 14340 9730
rect 14380 9690 14400 9730
rect 14320 9660 14400 9690
rect 14500 10230 14580 10260
rect 14500 10190 14520 10230
rect 14560 10190 14580 10230
rect 14500 10130 14580 10190
rect 14500 10090 14520 10130
rect 14560 10090 14580 10130
rect 14500 10030 14580 10090
rect 14500 9990 14520 10030
rect 14560 9990 14580 10030
rect 14500 9930 14580 9990
rect 14500 9890 14520 9930
rect 14560 9890 14580 9930
rect 14500 9830 14580 9890
rect 14500 9790 14520 9830
rect 14560 9790 14580 9830
rect 14500 9730 14580 9790
rect 14500 9690 14520 9730
rect 14560 9690 14580 9730
rect 14500 9660 14580 9690
rect 14680 10230 14760 10260
rect 14680 10190 14700 10230
rect 14740 10190 14760 10230
rect 14680 10130 14760 10190
rect 14680 10090 14700 10130
rect 14740 10090 14760 10130
rect 14680 10030 14760 10090
rect 14680 9990 14700 10030
rect 14740 9990 14760 10030
rect 14680 9930 14760 9990
rect 14680 9890 14700 9930
rect 14740 9890 14760 9930
rect 14680 9830 14760 9890
rect 14680 9790 14700 9830
rect 14740 9790 14760 9830
rect 14680 9730 14760 9790
rect 14680 9690 14700 9730
rect 14740 9690 14760 9730
rect 14680 9660 14760 9690
rect 14860 10230 14940 10260
rect 14860 10190 14880 10230
rect 14920 10190 14940 10230
rect 14860 10130 14940 10190
rect 14860 10090 14880 10130
rect 14920 10090 14940 10130
rect 14860 10030 14940 10090
rect 14860 9990 14880 10030
rect 14920 9990 14940 10030
rect 14860 9930 14940 9990
rect 14860 9890 14880 9930
rect 14920 9890 14940 9930
rect 14860 9830 14940 9890
rect 15480 10030 15570 10060
rect 15480 9990 15510 10030
rect 15550 9990 15570 10030
rect 15480 9930 15570 9990
rect 15480 9890 15510 9930
rect 15550 9890 15570 9930
rect 15480 9860 15570 9890
rect 15600 10030 15680 10060
rect 15600 9990 15620 10030
rect 15660 9990 15680 10030
rect 15600 9930 15680 9990
rect 15600 9890 15620 9930
rect 15660 9890 15680 9930
rect 15600 9860 15680 9890
rect 15710 10030 15790 10060
rect 15710 9990 15730 10030
rect 15770 9990 15790 10030
rect 15710 9930 15790 9990
rect 15710 9890 15730 9930
rect 15770 9890 15790 9930
rect 15710 9860 15790 9890
rect 15820 10030 15900 10060
rect 15820 9990 15840 10030
rect 15880 9990 15900 10030
rect 15820 9930 15900 9990
rect 15820 9890 15840 9930
rect 15880 9890 15900 9930
rect 15820 9860 15900 9890
rect 15930 10030 16010 10060
rect 15930 9990 15950 10030
rect 15990 9990 16010 10030
rect 15930 9930 16010 9990
rect 15930 9890 15950 9930
rect 15990 9890 16010 9930
rect 15930 9860 16010 9890
rect 14860 9790 14880 9830
rect 14920 9790 14940 9830
rect 14860 9730 14940 9790
rect 14860 9690 14880 9730
rect 14920 9690 14940 9730
rect 14860 9660 14940 9690
rect 11630 9230 11710 9260
rect 11630 9190 11650 9230
rect 11690 9190 11710 9230
rect 11630 9130 11710 9190
rect 11630 9090 11650 9130
rect 11690 9090 11710 9130
rect 11630 9060 11710 9090
rect 11740 9230 11820 9260
rect 11740 9190 11760 9230
rect 11800 9190 11820 9230
rect 11740 9130 11820 9190
rect 11740 9090 11760 9130
rect 11800 9090 11820 9130
rect 11740 9060 11820 9090
rect 11850 9230 11930 9260
rect 11850 9190 11870 9230
rect 11910 9190 11930 9230
rect 11850 9130 11930 9190
rect 11850 9090 11870 9130
rect 11910 9090 11930 9130
rect 11850 9060 11930 9090
rect 11960 9230 12040 9260
rect 11960 9190 11980 9230
rect 12020 9190 12040 9230
rect 11960 9130 12040 9190
rect 11960 9090 11980 9130
rect 12020 9090 12040 9130
rect 11960 9060 12040 9090
rect 12070 9230 12150 9260
rect 12070 9190 12090 9230
rect 12130 9190 12150 9230
rect 12070 9130 12150 9190
rect 12070 9090 12090 9130
rect 12130 9090 12150 9130
rect 12070 9060 12150 9090
rect 12180 9230 12260 9260
rect 12180 9190 12200 9230
rect 12240 9190 12260 9230
rect 12180 9130 12260 9190
rect 12180 9090 12200 9130
rect 12240 9090 12260 9130
rect 12180 9060 12260 9090
rect 12290 9230 12370 9260
rect 12290 9190 12310 9230
rect 12350 9190 12370 9230
rect 12290 9130 12370 9190
rect 12290 9090 12310 9130
rect 12350 9090 12370 9130
rect 12290 9060 12370 9090
rect 12400 9230 12480 9260
rect 12400 9190 12420 9230
rect 12460 9190 12480 9230
rect 12400 9130 12480 9190
rect 12400 9090 12420 9130
rect 12460 9090 12480 9130
rect 12400 9060 12480 9090
rect 12510 9230 12590 9260
rect 12510 9190 12530 9230
rect 12570 9190 12590 9230
rect 12510 9130 12590 9190
rect 12510 9090 12530 9130
rect 12570 9090 12590 9130
rect 12510 9060 12590 9090
rect 12620 9230 12700 9260
rect 12620 9190 12640 9230
rect 12680 9190 12700 9230
rect 12620 9130 12700 9190
rect 12620 9090 12640 9130
rect 12680 9090 12700 9130
rect 12620 9060 12700 9090
rect 12730 9230 12810 9260
rect 12730 9190 12750 9230
rect 12790 9190 12810 9230
rect 12730 9130 12810 9190
rect 12730 9090 12750 9130
rect 12790 9090 12810 9130
rect 12730 9060 12810 9090
rect 12840 9230 12920 9260
rect 12840 9190 12860 9230
rect 12900 9190 12920 9230
rect 12840 9130 12920 9190
rect 12840 9090 12860 9130
rect 12900 9090 12920 9130
rect 12840 9060 12920 9090
rect 12950 9230 13030 9260
rect 12950 9190 12970 9230
rect 13010 9190 13030 9230
rect 12950 9130 13030 9190
rect 12950 9090 12970 9130
rect 13010 9090 13030 9130
rect 12950 9060 13030 9090
rect 13530 9230 13610 9260
rect 13530 9190 13550 9230
rect 13590 9190 13610 9230
rect 13530 9130 13610 9190
rect 13530 9090 13550 9130
rect 13590 9090 13610 9130
rect 13530 9060 13610 9090
rect 13640 9230 13720 9260
rect 13640 9190 13660 9230
rect 13700 9190 13720 9230
rect 13640 9130 13720 9190
rect 13640 9090 13660 9130
rect 13700 9090 13720 9130
rect 13640 9060 13720 9090
rect 13750 9230 13830 9260
rect 13750 9190 13770 9230
rect 13810 9190 13830 9230
rect 13750 9130 13830 9190
rect 13750 9090 13770 9130
rect 13810 9090 13830 9130
rect 13750 9060 13830 9090
rect 13860 9230 13940 9260
rect 13860 9190 13880 9230
rect 13920 9190 13940 9230
rect 13860 9130 13940 9190
rect 13860 9090 13880 9130
rect 13920 9090 13940 9130
rect 13860 9060 13940 9090
rect 13970 9230 14050 9260
rect 13970 9190 13990 9230
rect 14030 9190 14050 9230
rect 13970 9130 14050 9190
rect 13970 9090 13990 9130
rect 14030 9090 14050 9130
rect 13970 9060 14050 9090
rect 14080 9230 14160 9260
rect 14080 9190 14100 9230
rect 14140 9190 14160 9230
rect 14080 9130 14160 9190
rect 14080 9090 14100 9130
rect 14140 9090 14160 9130
rect 14080 9060 14160 9090
rect 14190 9230 14270 9260
rect 14190 9190 14210 9230
rect 14250 9190 14270 9230
rect 14190 9130 14270 9190
rect 14190 9090 14210 9130
rect 14250 9090 14270 9130
rect 14190 9060 14270 9090
rect 14300 9230 14380 9260
rect 14300 9190 14320 9230
rect 14360 9190 14380 9230
rect 14300 9130 14380 9190
rect 14300 9090 14320 9130
rect 14360 9090 14380 9130
rect 14300 9060 14380 9090
rect 14410 9230 14490 9260
rect 14410 9190 14430 9230
rect 14470 9190 14490 9230
rect 14410 9130 14490 9190
rect 14410 9090 14430 9130
rect 14470 9090 14490 9130
rect 14410 9060 14490 9090
rect 14520 9230 14600 9260
rect 14520 9190 14540 9230
rect 14580 9190 14600 9230
rect 14520 9130 14600 9190
rect 14520 9090 14540 9130
rect 14580 9090 14600 9130
rect 14520 9060 14600 9090
rect 14630 9230 14710 9260
rect 14630 9190 14650 9230
rect 14690 9190 14710 9230
rect 14630 9130 14710 9190
rect 14630 9090 14650 9130
rect 14690 9090 14710 9130
rect 14630 9060 14710 9090
rect 14740 9230 14820 9260
rect 14740 9190 14760 9230
rect 14800 9190 14820 9230
rect 14740 9130 14820 9190
rect 14740 9090 14760 9130
rect 14800 9090 14820 9130
rect 14740 9060 14820 9090
rect 14850 9230 14930 9260
rect 14850 9190 14870 9230
rect 14910 9190 14930 9230
rect 14850 9130 14930 9190
rect 14850 9090 14870 9130
rect 14910 9090 14930 9130
rect 14850 9060 14930 9090
<< ndiffc >>
rect 11180 13810 11220 13850
rect 11180 13710 11220 13750
rect 13260 13810 13300 13850
rect 13260 13710 13300 13750
rect 15340 13810 15380 13850
rect 15340 13710 15380 13750
rect 10760 13200 10800 13240
rect 10760 13100 10800 13140
rect 10760 13000 10800 13040
rect 10760 12900 10800 12940
rect 10760 12800 10800 12840
rect 11840 13200 11880 13240
rect 12000 13200 12040 13240
rect 11840 13100 11880 13140
rect 12000 13100 12040 13140
rect 11840 13000 11880 13040
rect 12000 13000 12040 13040
rect 11840 12900 11880 12940
rect 12000 12900 12040 12940
rect 11840 12800 11880 12840
rect 12000 12800 12040 12840
rect 13080 13200 13120 13240
rect 13080 13100 13120 13140
rect 13080 13000 13120 13040
rect 13080 12900 13120 12940
rect 13080 12800 13120 12840
rect 13440 13200 13480 13240
rect 13440 13100 13480 13140
rect 13440 13000 13480 13040
rect 13440 12900 13480 12940
rect 13440 12800 13480 12840
rect 14520 13200 14560 13240
rect 14680 13200 14720 13240
rect 14520 13100 14560 13140
rect 14680 13100 14720 13140
rect 14520 13000 14560 13040
rect 14680 13000 14720 13040
rect 14520 12900 14560 12940
rect 14680 12900 14720 12940
rect 14520 12800 14560 12840
rect 14680 12800 14720 12840
rect 15760 13200 15800 13240
rect 15760 13100 15800 13140
rect 15760 13000 15800 13040
rect 15760 12900 15800 12940
rect 15760 12800 15800 12840
rect 11380 12190 11420 12230
rect 11500 12190 11540 12230
rect 11620 12190 11660 12230
rect 11740 12190 11780 12230
rect 11860 12190 11900 12230
rect 11980 12190 12020 12230
rect 12100 12190 12140 12230
rect 12220 12190 12260 12230
rect 12340 12190 12380 12230
rect 12460 12190 12500 12230
rect 12580 12190 12620 12230
rect 13940 12190 13980 12230
rect 14060 12190 14100 12230
rect 14180 12190 14220 12230
rect 14300 12190 14340 12230
rect 14420 12190 14460 12230
rect 14540 12190 14580 12230
rect 14660 12190 14700 12230
rect 14780 12190 14820 12230
rect 14900 12190 14940 12230
rect 15020 12190 15060 12230
rect 15140 12190 15180 12230
<< pdiffc >>
rect 11632 18392 11666 18426
rect 11722 18392 11756 18426
rect 11812 18392 11846 18426
rect 11902 18392 11936 18426
rect 11992 18392 12026 18426
rect 12082 18392 12116 18426
rect 12172 18392 12206 18426
rect 11632 18302 11666 18336
rect 11722 18302 11756 18336
rect 11812 18302 11846 18336
rect 11902 18302 11936 18336
rect 11992 18302 12026 18336
rect 12082 18302 12116 18336
rect 12172 18302 12206 18336
rect 11632 18212 11666 18246
rect 11722 18212 11756 18246
rect 11812 18212 11846 18246
rect 11902 18212 11936 18246
rect 11992 18212 12026 18246
rect 12082 18212 12116 18246
rect 12172 18212 12206 18246
rect 11632 18122 11666 18156
rect 11722 18122 11756 18156
rect 11812 18122 11846 18156
rect 11902 18122 11936 18156
rect 11992 18122 12026 18156
rect 12082 18122 12116 18156
rect 12172 18122 12206 18156
rect 11632 18032 11666 18066
rect 11722 18032 11756 18066
rect 11812 18032 11846 18066
rect 11902 18032 11936 18066
rect 11992 18032 12026 18066
rect 12082 18032 12116 18066
rect 12172 18032 12206 18066
rect 11632 17942 11666 17976
rect 11722 17942 11756 17976
rect 11812 17942 11846 17976
rect 11902 17942 11936 17976
rect 11992 17942 12026 17976
rect 12082 17942 12116 17976
rect 12172 17942 12206 17976
rect 11632 17852 11666 17886
rect 11722 17852 11756 17886
rect 11812 17852 11846 17886
rect 11902 17852 11936 17886
rect 11992 17852 12026 17886
rect 12082 17852 12116 17886
rect 12172 17852 12206 17886
rect 12992 18392 13026 18426
rect 13082 18392 13116 18426
rect 13172 18392 13206 18426
rect 13262 18392 13296 18426
rect 13352 18392 13386 18426
rect 13442 18392 13476 18426
rect 13532 18392 13566 18426
rect 12992 18302 13026 18336
rect 13082 18302 13116 18336
rect 13172 18302 13206 18336
rect 13262 18302 13296 18336
rect 13352 18302 13386 18336
rect 13442 18302 13476 18336
rect 13532 18302 13566 18336
rect 12992 18212 13026 18246
rect 13082 18212 13116 18246
rect 13172 18212 13206 18246
rect 13262 18212 13296 18246
rect 13352 18212 13386 18246
rect 13442 18212 13476 18246
rect 13532 18212 13566 18246
rect 12992 18122 13026 18156
rect 13082 18122 13116 18156
rect 13172 18122 13206 18156
rect 13262 18122 13296 18156
rect 13352 18122 13386 18156
rect 13442 18122 13476 18156
rect 13532 18122 13566 18156
rect 12992 18032 13026 18066
rect 13082 18032 13116 18066
rect 13172 18032 13206 18066
rect 13262 18032 13296 18066
rect 13352 18032 13386 18066
rect 13442 18032 13476 18066
rect 13532 18032 13566 18066
rect 12992 17942 13026 17976
rect 13082 17942 13116 17976
rect 13172 17942 13206 17976
rect 13262 17942 13296 17976
rect 13352 17942 13386 17976
rect 13442 17942 13476 17976
rect 13532 17942 13566 17976
rect 12992 17852 13026 17886
rect 13082 17852 13116 17886
rect 13172 17852 13206 17886
rect 13262 17852 13296 17886
rect 13352 17852 13386 17886
rect 13442 17852 13476 17886
rect 13532 17852 13566 17886
rect 14352 18392 14386 18426
rect 14442 18392 14476 18426
rect 14532 18392 14566 18426
rect 14622 18392 14656 18426
rect 14712 18392 14746 18426
rect 14802 18392 14836 18426
rect 14892 18392 14926 18426
rect 14352 18302 14386 18336
rect 14442 18302 14476 18336
rect 14532 18302 14566 18336
rect 14622 18302 14656 18336
rect 14712 18302 14746 18336
rect 14802 18302 14836 18336
rect 14892 18302 14926 18336
rect 14352 18212 14386 18246
rect 14442 18212 14476 18246
rect 14532 18212 14566 18246
rect 14622 18212 14656 18246
rect 14712 18212 14746 18246
rect 14802 18212 14836 18246
rect 14892 18212 14926 18246
rect 14352 18122 14386 18156
rect 14442 18122 14476 18156
rect 14532 18122 14566 18156
rect 14622 18122 14656 18156
rect 14712 18122 14746 18156
rect 14802 18122 14836 18156
rect 14892 18122 14926 18156
rect 14352 18032 14386 18066
rect 14442 18032 14476 18066
rect 14532 18032 14566 18066
rect 14622 18032 14656 18066
rect 14712 18032 14746 18066
rect 14802 18032 14836 18066
rect 14892 18032 14926 18066
rect 14352 17942 14386 17976
rect 14442 17942 14476 17976
rect 14532 17942 14566 17976
rect 14622 17942 14656 17976
rect 14712 17942 14746 17976
rect 14802 17942 14836 17976
rect 14892 17942 14926 17976
rect 14352 17852 14386 17886
rect 14442 17852 14476 17886
rect 14532 17852 14566 17886
rect 14622 17852 14656 17886
rect 14712 17852 14746 17886
rect 14802 17852 14836 17886
rect 14892 17852 14926 17886
rect 11632 17032 11666 17066
rect 11722 17032 11756 17066
rect 11812 17032 11846 17066
rect 11902 17032 11936 17066
rect 11992 17032 12026 17066
rect 12082 17032 12116 17066
rect 12172 17032 12206 17066
rect 11632 16942 11666 16976
rect 11722 16942 11756 16976
rect 11812 16942 11846 16976
rect 11902 16942 11936 16976
rect 11992 16942 12026 16976
rect 12082 16942 12116 16976
rect 12172 16942 12206 16976
rect 11632 16852 11666 16886
rect 11722 16852 11756 16886
rect 11812 16852 11846 16886
rect 11902 16852 11936 16886
rect 11992 16852 12026 16886
rect 12082 16852 12116 16886
rect 12172 16852 12206 16886
rect 11632 16762 11666 16796
rect 11722 16762 11756 16796
rect 11812 16762 11846 16796
rect 11902 16762 11936 16796
rect 11992 16762 12026 16796
rect 12082 16762 12116 16796
rect 12172 16762 12206 16796
rect 11632 16672 11666 16706
rect 11722 16672 11756 16706
rect 11812 16672 11846 16706
rect 11902 16672 11936 16706
rect 11992 16672 12026 16706
rect 12082 16672 12116 16706
rect 12172 16672 12206 16706
rect 11632 16582 11666 16616
rect 11722 16582 11756 16616
rect 11812 16582 11846 16616
rect 11902 16582 11936 16616
rect 11992 16582 12026 16616
rect 12082 16582 12116 16616
rect 12172 16582 12206 16616
rect 11632 16492 11666 16526
rect 11722 16492 11756 16526
rect 11812 16492 11846 16526
rect 11902 16492 11936 16526
rect 11992 16492 12026 16526
rect 12082 16492 12116 16526
rect 12172 16492 12206 16526
rect 12992 17032 13026 17066
rect 13082 17032 13116 17066
rect 13172 17032 13206 17066
rect 13262 17032 13296 17066
rect 13352 17032 13386 17066
rect 13442 17032 13476 17066
rect 13532 17032 13566 17066
rect 12992 16942 13026 16976
rect 13082 16942 13116 16976
rect 13172 16942 13206 16976
rect 13262 16942 13296 16976
rect 13352 16942 13386 16976
rect 13442 16942 13476 16976
rect 13532 16942 13566 16976
rect 12992 16852 13026 16886
rect 13082 16852 13116 16886
rect 13172 16852 13206 16886
rect 13262 16852 13296 16886
rect 13352 16852 13386 16886
rect 13442 16852 13476 16886
rect 13532 16852 13566 16886
rect 12992 16762 13026 16796
rect 13082 16762 13116 16796
rect 13172 16762 13206 16796
rect 13262 16762 13296 16796
rect 13352 16762 13386 16796
rect 13442 16762 13476 16796
rect 13532 16762 13566 16796
rect 12992 16672 13026 16706
rect 13082 16672 13116 16706
rect 13172 16672 13206 16706
rect 13262 16672 13296 16706
rect 13352 16672 13386 16706
rect 13442 16672 13476 16706
rect 13532 16672 13566 16706
rect 12992 16582 13026 16616
rect 13082 16582 13116 16616
rect 13172 16582 13206 16616
rect 13262 16582 13296 16616
rect 13352 16582 13386 16616
rect 13442 16582 13476 16616
rect 13532 16582 13566 16616
rect 12992 16492 13026 16526
rect 13082 16492 13116 16526
rect 13172 16492 13206 16526
rect 13262 16492 13296 16526
rect 13352 16492 13386 16526
rect 13442 16492 13476 16526
rect 13532 16492 13566 16526
rect 14352 17032 14386 17066
rect 14442 17032 14476 17066
rect 14532 17032 14566 17066
rect 14622 17032 14656 17066
rect 14712 17032 14746 17066
rect 14802 17032 14836 17066
rect 14892 17032 14926 17066
rect 14352 16942 14386 16976
rect 14442 16942 14476 16976
rect 14532 16942 14566 16976
rect 14622 16942 14656 16976
rect 14712 16942 14746 16976
rect 14802 16942 14836 16976
rect 14892 16942 14926 16976
rect 14352 16852 14386 16886
rect 14442 16852 14476 16886
rect 14532 16852 14566 16886
rect 14622 16852 14656 16886
rect 14712 16852 14746 16886
rect 14802 16852 14836 16886
rect 14892 16852 14926 16886
rect 14352 16762 14386 16796
rect 14442 16762 14476 16796
rect 14532 16762 14566 16796
rect 14622 16762 14656 16796
rect 14712 16762 14746 16796
rect 14802 16762 14836 16796
rect 14892 16762 14926 16796
rect 14352 16672 14386 16706
rect 14442 16672 14476 16706
rect 14532 16672 14566 16706
rect 14622 16672 14656 16706
rect 14712 16672 14746 16706
rect 14802 16672 14836 16706
rect 14892 16672 14926 16706
rect 14352 16582 14386 16616
rect 14442 16582 14476 16616
rect 14532 16582 14566 16616
rect 14622 16582 14656 16616
rect 14712 16582 14746 16616
rect 14802 16582 14836 16616
rect 14892 16582 14926 16616
rect 14352 16492 14386 16526
rect 14442 16492 14476 16526
rect 14532 16492 14566 16526
rect 14622 16492 14656 16526
rect 14712 16492 14746 16526
rect 14802 16492 14836 16526
rect 14892 16492 14926 16526
rect 11632 15672 11666 15706
rect 11722 15672 11756 15706
rect 11812 15672 11846 15706
rect 11902 15672 11936 15706
rect 11992 15672 12026 15706
rect 12082 15672 12116 15706
rect 12172 15672 12206 15706
rect 11632 15582 11666 15616
rect 11722 15582 11756 15616
rect 11812 15582 11846 15616
rect 11902 15582 11936 15616
rect 11992 15582 12026 15616
rect 12082 15582 12116 15616
rect 12172 15582 12206 15616
rect 11632 15492 11666 15526
rect 11722 15492 11756 15526
rect 11812 15492 11846 15526
rect 11902 15492 11936 15526
rect 11992 15492 12026 15526
rect 12082 15492 12116 15526
rect 12172 15492 12206 15526
rect 11632 15402 11666 15436
rect 11722 15402 11756 15436
rect 11812 15402 11846 15436
rect 11902 15402 11936 15436
rect 11992 15402 12026 15436
rect 12082 15402 12116 15436
rect 12172 15402 12206 15436
rect 11632 15312 11666 15346
rect 11722 15312 11756 15346
rect 11812 15312 11846 15346
rect 11902 15312 11936 15346
rect 11992 15312 12026 15346
rect 12082 15312 12116 15346
rect 12172 15312 12206 15346
rect 11632 15222 11666 15256
rect 11722 15222 11756 15256
rect 11812 15222 11846 15256
rect 11902 15222 11936 15256
rect 11992 15222 12026 15256
rect 12082 15222 12116 15256
rect 12172 15222 12206 15256
rect 11632 15132 11666 15166
rect 11722 15132 11756 15166
rect 11812 15132 11846 15166
rect 11902 15132 11936 15166
rect 11992 15132 12026 15166
rect 12082 15132 12116 15166
rect 12172 15132 12206 15166
rect 12992 15672 13026 15706
rect 13082 15672 13116 15706
rect 13172 15672 13206 15706
rect 13262 15672 13296 15706
rect 13352 15672 13386 15706
rect 13442 15672 13476 15706
rect 13532 15672 13566 15706
rect 12992 15582 13026 15616
rect 13082 15582 13116 15616
rect 13172 15582 13206 15616
rect 13262 15582 13296 15616
rect 13352 15582 13386 15616
rect 13442 15582 13476 15616
rect 13532 15582 13566 15616
rect 12992 15492 13026 15526
rect 13082 15492 13116 15526
rect 13172 15492 13206 15526
rect 13262 15492 13296 15526
rect 13352 15492 13386 15526
rect 13442 15492 13476 15526
rect 13532 15492 13566 15526
rect 12992 15402 13026 15436
rect 13082 15402 13116 15436
rect 13172 15402 13206 15436
rect 13262 15402 13296 15436
rect 13352 15402 13386 15436
rect 13442 15402 13476 15436
rect 13532 15402 13566 15436
rect 12992 15312 13026 15346
rect 13082 15312 13116 15346
rect 13172 15312 13206 15346
rect 13262 15312 13296 15346
rect 13352 15312 13386 15346
rect 13442 15312 13476 15346
rect 13532 15312 13566 15346
rect 12992 15222 13026 15256
rect 13082 15222 13116 15256
rect 13172 15222 13206 15256
rect 13262 15222 13296 15256
rect 13352 15222 13386 15256
rect 13442 15222 13476 15256
rect 13532 15222 13566 15256
rect 12992 15132 13026 15166
rect 13082 15132 13116 15166
rect 13172 15132 13206 15166
rect 13262 15132 13296 15166
rect 13352 15132 13386 15166
rect 13442 15132 13476 15166
rect 13532 15132 13566 15166
rect 14352 15672 14386 15706
rect 14442 15672 14476 15706
rect 14532 15672 14566 15706
rect 14622 15672 14656 15706
rect 14712 15672 14746 15706
rect 14802 15672 14836 15706
rect 14892 15672 14926 15706
rect 14352 15582 14386 15616
rect 14442 15582 14476 15616
rect 14532 15582 14566 15616
rect 14622 15582 14656 15616
rect 14712 15582 14746 15616
rect 14802 15582 14836 15616
rect 14892 15582 14926 15616
rect 14352 15492 14386 15526
rect 14442 15492 14476 15526
rect 14532 15492 14566 15526
rect 14622 15492 14656 15526
rect 14712 15492 14746 15526
rect 14802 15492 14836 15526
rect 14892 15492 14926 15526
rect 14352 15402 14386 15436
rect 14442 15402 14476 15436
rect 14532 15402 14566 15436
rect 14622 15402 14656 15436
rect 14712 15402 14746 15436
rect 14802 15402 14836 15436
rect 14892 15402 14926 15436
rect 14352 15312 14386 15346
rect 14442 15312 14476 15346
rect 14532 15312 14566 15346
rect 14622 15312 14656 15346
rect 14712 15312 14746 15346
rect 14802 15312 14836 15346
rect 14892 15312 14926 15346
rect 14352 15222 14386 15256
rect 14442 15222 14476 15256
rect 14532 15222 14566 15256
rect 14622 15222 14656 15256
rect 14712 15222 14746 15256
rect 14802 15222 14836 15256
rect 14892 15222 14926 15256
rect 14352 15132 14386 15166
rect 14442 15132 14476 15166
rect 14532 15132 14566 15166
rect 14622 15132 14656 15166
rect 14712 15132 14746 15166
rect 14802 15132 14836 15166
rect 14892 15132 14926 15166
rect 10540 11350 10580 11390
rect 10540 11250 10580 11290
rect 10660 11350 10700 11390
rect 10660 11250 10700 11290
rect 10780 11350 10820 11390
rect 10780 11250 10820 11290
rect 10900 11350 10940 11390
rect 10900 11250 10940 11290
rect 11020 11350 11060 11390
rect 11020 11250 11060 11290
rect 11140 11350 11180 11390
rect 11140 11250 11180 11290
rect 11260 11350 11300 11390
rect 11260 11250 11300 11290
rect 11380 11350 11420 11390
rect 11380 11250 11420 11290
rect 11500 11350 11540 11390
rect 11500 11250 11540 11290
rect 11620 11350 11660 11390
rect 11620 11250 11660 11290
rect 11740 11350 11780 11390
rect 11740 11250 11780 11290
rect 11860 11350 11900 11390
rect 11860 11250 11900 11290
rect 11980 11350 12020 11390
rect 11980 11250 12020 11290
rect 12100 11350 12140 11390
rect 12100 11250 12140 11290
rect 12220 11350 12260 11390
rect 12220 11250 12260 11290
rect 12340 11350 12380 11390
rect 12340 11250 12380 11290
rect 12460 11350 12500 11390
rect 12460 11250 12500 11290
rect 12580 11350 12620 11390
rect 12580 11250 12620 11290
rect 12700 11350 12740 11390
rect 12700 11250 12740 11290
rect 12820 11350 12860 11390
rect 12820 11250 12860 11290
rect 12940 11350 12980 11390
rect 12940 11250 12980 11290
rect 13580 11350 13620 11390
rect 13580 11250 13620 11290
rect 13700 11350 13740 11390
rect 13700 11250 13740 11290
rect 13820 11350 13860 11390
rect 13820 11250 13860 11290
rect 13940 11350 13980 11390
rect 13940 11250 13980 11290
rect 14060 11350 14100 11390
rect 14060 11250 14100 11290
rect 14180 11350 14220 11390
rect 14180 11250 14220 11290
rect 14300 11350 14340 11390
rect 14300 11250 14340 11290
rect 14420 11350 14460 11390
rect 14420 11250 14460 11290
rect 14540 11350 14580 11390
rect 14540 11250 14580 11290
rect 14660 11350 14700 11390
rect 14660 11250 14700 11290
rect 14780 11350 14820 11390
rect 14780 11250 14820 11290
rect 14900 11350 14940 11390
rect 14900 11250 14940 11290
rect 15020 11350 15060 11390
rect 15020 11250 15060 11290
rect 15140 11350 15180 11390
rect 15140 11250 15180 11290
rect 15260 11350 15300 11390
rect 15260 11250 15300 11290
rect 15380 11350 15420 11390
rect 15380 11250 15420 11290
rect 15500 11350 15540 11390
rect 15500 11250 15540 11290
rect 15620 11350 15660 11390
rect 15620 11250 15660 11290
rect 15740 11350 15780 11390
rect 15740 11250 15780 11290
rect 15860 11350 15900 11390
rect 15860 11250 15900 11290
rect 15980 11350 16020 11390
rect 15980 11250 16020 11290
rect 11640 10190 11680 10230
rect 11640 10090 11680 10130
rect 11640 9990 11680 10030
rect 11640 9890 11680 9930
rect 11640 9790 11680 9830
rect 11640 9690 11680 9730
rect 11820 10190 11860 10230
rect 11820 10090 11860 10130
rect 11820 9990 11860 10030
rect 11820 9890 11860 9930
rect 11820 9790 11860 9830
rect 11820 9690 11860 9730
rect 12000 10190 12040 10230
rect 12000 10090 12040 10130
rect 12000 9990 12040 10030
rect 12000 9890 12040 9930
rect 12000 9790 12040 9830
rect 12000 9690 12040 9730
rect 12180 10190 12220 10230
rect 12180 10090 12220 10130
rect 12180 9990 12220 10030
rect 12180 9890 12220 9930
rect 12180 9790 12220 9830
rect 12180 9690 12220 9730
rect 12360 10190 12400 10230
rect 12360 10090 12400 10130
rect 12360 9990 12400 10030
rect 12360 9890 12400 9930
rect 12360 9790 12400 9830
rect 12360 9690 12400 9730
rect 12540 10190 12580 10230
rect 12540 10090 12580 10130
rect 12540 9990 12580 10030
rect 12540 9890 12580 9930
rect 12540 9790 12580 9830
rect 12540 9690 12580 9730
rect 12720 10190 12760 10230
rect 12720 10090 12760 10130
rect 12720 9990 12760 10030
rect 12720 9890 12760 9930
rect 12720 9790 12760 9830
rect 12720 9690 12760 9730
rect 12900 10190 12940 10230
rect 12900 10090 12940 10130
rect 12900 9990 12940 10030
rect 12900 9890 12940 9930
rect 12900 9790 12940 9830
rect 12900 9690 12940 9730
rect 13080 10190 13120 10230
rect 13080 10090 13120 10130
rect 13080 9990 13120 10030
rect 13080 9890 13120 9930
rect 13080 9790 13120 9830
rect 13080 9690 13120 9730
rect 13260 10190 13300 10230
rect 13260 10090 13300 10130
rect 13260 9990 13300 10030
rect 13260 9890 13300 9930
rect 13260 9790 13300 9830
rect 13260 9690 13300 9730
rect 13440 10190 13480 10230
rect 13440 10090 13480 10130
rect 13440 9990 13480 10030
rect 13440 9890 13480 9930
rect 13440 9790 13480 9830
rect 13440 9690 13480 9730
rect 13620 10190 13660 10230
rect 13620 10090 13660 10130
rect 13620 9990 13660 10030
rect 13620 9890 13660 9930
rect 13620 9790 13660 9830
rect 13620 9690 13660 9730
rect 13800 10190 13840 10230
rect 13800 10090 13840 10130
rect 13800 9990 13840 10030
rect 13800 9890 13840 9930
rect 13800 9790 13840 9830
rect 13800 9690 13840 9730
rect 13980 10190 14020 10230
rect 13980 10090 14020 10130
rect 13980 9990 14020 10030
rect 13980 9890 14020 9930
rect 13980 9790 14020 9830
rect 13980 9690 14020 9730
rect 14160 10190 14200 10230
rect 14160 10090 14200 10130
rect 14160 9990 14200 10030
rect 14160 9890 14200 9930
rect 14160 9790 14200 9830
rect 14160 9690 14200 9730
rect 14340 10190 14380 10230
rect 14340 10090 14380 10130
rect 14340 9990 14380 10030
rect 14340 9890 14380 9930
rect 14340 9790 14380 9830
rect 14340 9690 14380 9730
rect 14520 10190 14560 10230
rect 14520 10090 14560 10130
rect 14520 9990 14560 10030
rect 14520 9890 14560 9930
rect 14520 9790 14560 9830
rect 14520 9690 14560 9730
rect 14700 10190 14740 10230
rect 14700 10090 14740 10130
rect 14700 9990 14740 10030
rect 14700 9890 14740 9930
rect 14700 9790 14740 9830
rect 14700 9690 14740 9730
rect 14880 10190 14920 10230
rect 14880 10090 14920 10130
rect 14880 9990 14920 10030
rect 14880 9890 14920 9930
rect 15510 9990 15550 10030
rect 15510 9890 15550 9930
rect 15620 9990 15660 10030
rect 15620 9890 15660 9930
rect 15730 9990 15770 10030
rect 15730 9890 15770 9930
rect 15840 9990 15880 10030
rect 15840 9890 15880 9930
rect 15950 9990 15990 10030
rect 15950 9890 15990 9930
rect 14880 9790 14920 9830
rect 14880 9690 14920 9730
rect 11650 9190 11690 9230
rect 11650 9090 11690 9130
rect 11760 9190 11800 9230
rect 11760 9090 11800 9130
rect 11870 9190 11910 9230
rect 11870 9090 11910 9130
rect 11980 9190 12020 9230
rect 11980 9090 12020 9130
rect 12090 9190 12130 9230
rect 12090 9090 12130 9130
rect 12200 9190 12240 9230
rect 12200 9090 12240 9130
rect 12310 9190 12350 9230
rect 12310 9090 12350 9130
rect 12420 9190 12460 9230
rect 12420 9090 12460 9130
rect 12530 9190 12570 9230
rect 12530 9090 12570 9130
rect 12640 9190 12680 9230
rect 12640 9090 12680 9130
rect 12750 9190 12790 9230
rect 12750 9090 12790 9130
rect 12860 9190 12900 9230
rect 12860 9090 12900 9130
rect 12970 9190 13010 9230
rect 12970 9090 13010 9130
rect 13550 9190 13590 9230
rect 13550 9090 13590 9130
rect 13660 9190 13700 9230
rect 13660 9090 13700 9130
rect 13770 9190 13810 9230
rect 13770 9090 13810 9130
rect 13880 9190 13920 9230
rect 13880 9090 13920 9130
rect 13990 9190 14030 9230
rect 13990 9090 14030 9130
rect 14100 9190 14140 9230
rect 14100 9090 14140 9130
rect 14210 9190 14250 9230
rect 14210 9090 14250 9130
rect 14320 9190 14360 9230
rect 14320 9090 14360 9130
rect 14430 9190 14470 9230
rect 14430 9090 14470 9130
rect 14540 9190 14580 9230
rect 14540 9090 14580 9130
rect 14650 9190 14690 9230
rect 14650 9090 14690 9130
rect 14760 9190 14800 9230
rect 14760 9090 14800 9130
rect 14870 9190 14910 9230
rect 14870 9090 14910 9130
<< psubdiff >>
rect 13230 19070 13330 19100
rect 13230 19030 13260 19070
rect 13300 19030 13330 19070
rect 13230 18990 13330 19030
rect 13230 18950 13260 18990
rect 13300 18950 13330 18990
rect 13230 18910 13330 18950
rect 13230 18870 13260 18910
rect 13300 18870 13330 18910
rect 13230 18840 13330 18870
rect 11276 18752 12564 18784
rect 11276 18718 11410 18752
rect 11444 18718 11500 18752
rect 11534 18718 11590 18752
rect 11624 18718 11680 18752
rect 11714 18718 11770 18752
rect 11804 18718 11860 18752
rect 11894 18718 11950 18752
rect 11984 18718 12040 18752
rect 12074 18718 12130 18752
rect 12164 18718 12220 18752
rect 12254 18718 12310 18752
rect 12344 18718 12400 18752
rect 12434 18718 12564 18752
rect 11276 18683 12564 18718
rect 11276 18668 11377 18683
rect 11276 18634 11309 18668
rect 11343 18634 11377 18668
rect 11276 18578 11377 18634
rect 12463 18668 12564 18683
rect 12463 18634 12496 18668
rect 12530 18634 12564 18668
rect 11276 18544 11309 18578
rect 11343 18544 11377 18578
rect 11276 18488 11377 18544
rect 11276 18454 11309 18488
rect 11343 18454 11377 18488
rect 11276 18398 11377 18454
rect 11276 18364 11309 18398
rect 11343 18364 11377 18398
rect 11276 18308 11377 18364
rect 11276 18274 11309 18308
rect 11343 18274 11377 18308
rect 11276 18218 11377 18274
rect 11276 18184 11309 18218
rect 11343 18184 11377 18218
rect 11276 18128 11377 18184
rect 11276 18094 11309 18128
rect 11343 18094 11377 18128
rect 11276 18038 11377 18094
rect 11276 18004 11309 18038
rect 11343 18004 11377 18038
rect 11276 17948 11377 18004
rect 11276 17914 11309 17948
rect 11343 17914 11377 17948
rect 11276 17858 11377 17914
rect 11276 17824 11309 17858
rect 11343 17824 11377 17858
rect 11276 17768 11377 17824
rect 11276 17734 11309 17768
rect 11343 17734 11377 17768
rect 11276 17678 11377 17734
rect 11276 17644 11309 17678
rect 11343 17644 11377 17678
rect 12463 18578 12564 18634
rect 12463 18544 12496 18578
rect 12530 18544 12564 18578
rect 12463 18488 12564 18544
rect 12463 18454 12496 18488
rect 12530 18454 12564 18488
rect 12463 18398 12564 18454
rect 12463 18364 12496 18398
rect 12530 18364 12564 18398
rect 12463 18308 12564 18364
rect 12463 18274 12496 18308
rect 12530 18274 12564 18308
rect 12463 18218 12564 18274
rect 12463 18184 12496 18218
rect 12530 18184 12564 18218
rect 12463 18128 12564 18184
rect 12463 18094 12496 18128
rect 12530 18094 12564 18128
rect 12463 18038 12564 18094
rect 12463 18004 12496 18038
rect 12530 18004 12564 18038
rect 12463 17948 12564 18004
rect 12463 17914 12496 17948
rect 12530 17914 12564 17948
rect 12463 17858 12564 17914
rect 12463 17824 12496 17858
rect 12530 17824 12564 17858
rect 12463 17768 12564 17824
rect 12463 17734 12496 17768
rect 12530 17734 12564 17768
rect 12463 17678 12564 17734
rect 11276 17597 11377 17644
rect 12463 17644 12496 17678
rect 12530 17644 12564 17678
rect 12463 17597 12564 17644
rect 11276 17588 12564 17597
rect 11276 17554 11309 17588
rect 11343 17565 12496 17588
rect 11343 17554 11410 17565
rect 11276 17531 11410 17554
rect 11444 17531 11500 17565
rect 11534 17531 11590 17565
rect 11624 17531 11680 17565
rect 11714 17531 11770 17565
rect 11804 17531 11860 17565
rect 11894 17531 11950 17565
rect 11984 17531 12040 17565
rect 12074 17531 12130 17565
rect 12164 17531 12220 17565
rect 12254 17531 12310 17565
rect 12344 17531 12400 17565
rect 12434 17554 12496 17565
rect 12530 17554 12564 17588
rect 12434 17531 12564 17554
rect 11276 17496 12564 17531
rect 12636 18752 13924 18784
rect 12636 18718 12770 18752
rect 12804 18718 12860 18752
rect 12894 18718 12950 18752
rect 12984 18718 13040 18752
rect 13074 18718 13130 18752
rect 13164 18718 13220 18752
rect 13254 18718 13310 18752
rect 13344 18718 13400 18752
rect 13434 18718 13490 18752
rect 13524 18718 13580 18752
rect 13614 18718 13670 18752
rect 13704 18718 13760 18752
rect 13794 18718 13924 18752
rect 12636 18683 13924 18718
rect 12636 18668 12737 18683
rect 12636 18634 12669 18668
rect 12703 18634 12737 18668
rect 12636 18578 12737 18634
rect 13823 18668 13924 18683
rect 13823 18634 13856 18668
rect 13890 18634 13924 18668
rect 12636 18544 12669 18578
rect 12703 18544 12737 18578
rect 12636 18488 12737 18544
rect 12636 18454 12669 18488
rect 12703 18454 12737 18488
rect 12636 18398 12737 18454
rect 12636 18364 12669 18398
rect 12703 18364 12737 18398
rect 12636 18308 12737 18364
rect 12636 18274 12669 18308
rect 12703 18274 12737 18308
rect 12636 18218 12737 18274
rect 12636 18184 12669 18218
rect 12703 18184 12737 18218
rect 12636 18128 12737 18184
rect 12636 18094 12669 18128
rect 12703 18094 12737 18128
rect 12636 18038 12737 18094
rect 12636 18004 12669 18038
rect 12703 18004 12737 18038
rect 12636 17948 12737 18004
rect 12636 17914 12669 17948
rect 12703 17914 12737 17948
rect 12636 17858 12737 17914
rect 12636 17824 12669 17858
rect 12703 17824 12737 17858
rect 12636 17768 12737 17824
rect 12636 17734 12669 17768
rect 12703 17734 12737 17768
rect 12636 17678 12737 17734
rect 12636 17644 12669 17678
rect 12703 17644 12737 17678
rect 13823 18578 13924 18634
rect 13823 18544 13856 18578
rect 13890 18544 13924 18578
rect 13823 18488 13924 18544
rect 13823 18454 13856 18488
rect 13890 18454 13924 18488
rect 13823 18398 13924 18454
rect 13823 18364 13856 18398
rect 13890 18364 13924 18398
rect 13823 18308 13924 18364
rect 13823 18274 13856 18308
rect 13890 18274 13924 18308
rect 13823 18218 13924 18274
rect 13823 18184 13856 18218
rect 13890 18184 13924 18218
rect 13823 18128 13924 18184
rect 13823 18094 13856 18128
rect 13890 18094 13924 18128
rect 13823 18038 13924 18094
rect 13823 18004 13856 18038
rect 13890 18004 13924 18038
rect 13823 17948 13924 18004
rect 13823 17914 13856 17948
rect 13890 17914 13924 17948
rect 13823 17858 13924 17914
rect 13823 17824 13856 17858
rect 13890 17824 13924 17858
rect 13823 17768 13924 17824
rect 13823 17734 13856 17768
rect 13890 17734 13924 17768
rect 13823 17678 13924 17734
rect 12636 17597 12737 17644
rect 13823 17644 13856 17678
rect 13890 17644 13924 17678
rect 13823 17597 13924 17644
rect 12636 17588 13924 17597
rect 12636 17554 12669 17588
rect 12703 17565 13856 17588
rect 12703 17554 12770 17565
rect 12636 17531 12770 17554
rect 12804 17531 12860 17565
rect 12894 17531 12950 17565
rect 12984 17531 13040 17565
rect 13074 17531 13130 17565
rect 13164 17531 13220 17565
rect 13254 17531 13310 17565
rect 13344 17531 13400 17565
rect 13434 17531 13490 17565
rect 13524 17531 13580 17565
rect 13614 17531 13670 17565
rect 13704 17531 13760 17565
rect 13794 17554 13856 17565
rect 13890 17554 13924 17588
rect 13794 17531 13924 17554
rect 12636 17496 13924 17531
rect 13996 18752 15284 18784
rect 13996 18718 14130 18752
rect 14164 18718 14220 18752
rect 14254 18718 14310 18752
rect 14344 18718 14400 18752
rect 14434 18718 14490 18752
rect 14524 18718 14580 18752
rect 14614 18718 14670 18752
rect 14704 18718 14760 18752
rect 14794 18718 14850 18752
rect 14884 18718 14940 18752
rect 14974 18718 15030 18752
rect 15064 18718 15120 18752
rect 15154 18718 15284 18752
rect 13996 18683 15284 18718
rect 13996 18668 14097 18683
rect 13996 18634 14029 18668
rect 14063 18634 14097 18668
rect 13996 18578 14097 18634
rect 15183 18668 15284 18683
rect 15183 18634 15216 18668
rect 15250 18634 15284 18668
rect 13996 18544 14029 18578
rect 14063 18544 14097 18578
rect 13996 18488 14097 18544
rect 13996 18454 14029 18488
rect 14063 18454 14097 18488
rect 13996 18398 14097 18454
rect 13996 18364 14029 18398
rect 14063 18364 14097 18398
rect 13996 18308 14097 18364
rect 13996 18274 14029 18308
rect 14063 18274 14097 18308
rect 13996 18218 14097 18274
rect 13996 18184 14029 18218
rect 14063 18184 14097 18218
rect 13996 18128 14097 18184
rect 13996 18094 14029 18128
rect 14063 18094 14097 18128
rect 13996 18038 14097 18094
rect 13996 18004 14029 18038
rect 14063 18004 14097 18038
rect 13996 17948 14097 18004
rect 13996 17914 14029 17948
rect 14063 17914 14097 17948
rect 13996 17858 14097 17914
rect 13996 17824 14029 17858
rect 14063 17824 14097 17858
rect 13996 17768 14097 17824
rect 13996 17734 14029 17768
rect 14063 17734 14097 17768
rect 13996 17678 14097 17734
rect 13996 17644 14029 17678
rect 14063 17644 14097 17678
rect 15183 18578 15284 18634
rect 15183 18544 15216 18578
rect 15250 18544 15284 18578
rect 15183 18488 15284 18544
rect 15183 18454 15216 18488
rect 15250 18454 15284 18488
rect 15183 18398 15284 18454
rect 15183 18364 15216 18398
rect 15250 18364 15284 18398
rect 15183 18308 15284 18364
rect 15183 18274 15216 18308
rect 15250 18274 15284 18308
rect 15183 18218 15284 18274
rect 15183 18184 15216 18218
rect 15250 18184 15284 18218
rect 15183 18128 15284 18184
rect 15183 18094 15216 18128
rect 15250 18094 15284 18128
rect 15183 18038 15284 18094
rect 15183 18004 15216 18038
rect 15250 18004 15284 18038
rect 15183 17948 15284 18004
rect 15183 17914 15216 17948
rect 15250 17914 15284 17948
rect 15183 17858 15284 17914
rect 15183 17824 15216 17858
rect 15250 17824 15284 17858
rect 15183 17768 15284 17824
rect 15183 17734 15216 17768
rect 15250 17734 15284 17768
rect 15183 17678 15284 17734
rect 13996 17597 14097 17644
rect 15183 17644 15216 17678
rect 15250 17644 15284 17678
rect 15183 17597 15284 17644
rect 13996 17588 15284 17597
rect 13996 17554 14029 17588
rect 14063 17565 15216 17588
rect 14063 17554 14130 17565
rect 13996 17531 14130 17554
rect 14164 17531 14220 17565
rect 14254 17531 14310 17565
rect 14344 17531 14400 17565
rect 14434 17531 14490 17565
rect 14524 17531 14580 17565
rect 14614 17531 14670 17565
rect 14704 17531 14760 17565
rect 14794 17531 14850 17565
rect 14884 17531 14940 17565
rect 14974 17531 15030 17565
rect 15064 17531 15120 17565
rect 15154 17554 15216 17565
rect 15250 17554 15284 17588
rect 15154 17531 15284 17554
rect 13996 17496 15284 17531
rect 11276 17392 12564 17424
rect 11276 17358 11410 17392
rect 11444 17358 11500 17392
rect 11534 17358 11590 17392
rect 11624 17358 11680 17392
rect 11714 17358 11770 17392
rect 11804 17358 11860 17392
rect 11894 17358 11950 17392
rect 11984 17358 12040 17392
rect 12074 17358 12130 17392
rect 12164 17358 12220 17392
rect 12254 17358 12310 17392
rect 12344 17358 12400 17392
rect 12434 17358 12564 17392
rect 11276 17323 12564 17358
rect 11276 17308 11377 17323
rect 11276 17274 11309 17308
rect 11343 17274 11377 17308
rect 11276 17218 11377 17274
rect 12463 17308 12564 17323
rect 12463 17274 12496 17308
rect 12530 17274 12564 17308
rect 11276 17184 11309 17218
rect 11343 17184 11377 17218
rect 11276 17128 11377 17184
rect 11276 17094 11309 17128
rect 11343 17094 11377 17128
rect 11276 17038 11377 17094
rect 11276 17004 11309 17038
rect 11343 17004 11377 17038
rect 11276 16948 11377 17004
rect 11276 16914 11309 16948
rect 11343 16914 11377 16948
rect 11276 16858 11377 16914
rect 11276 16824 11309 16858
rect 11343 16824 11377 16858
rect 11276 16768 11377 16824
rect 11276 16734 11309 16768
rect 11343 16734 11377 16768
rect 11276 16678 11377 16734
rect 11276 16644 11309 16678
rect 11343 16644 11377 16678
rect 11276 16588 11377 16644
rect 11276 16554 11309 16588
rect 11343 16554 11377 16588
rect 11276 16498 11377 16554
rect 11276 16464 11309 16498
rect 11343 16464 11377 16498
rect 11276 16408 11377 16464
rect 11276 16374 11309 16408
rect 11343 16374 11377 16408
rect 11276 16318 11377 16374
rect 11276 16284 11309 16318
rect 11343 16284 11377 16318
rect 12463 17218 12564 17274
rect 12463 17184 12496 17218
rect 12530 17184 12564 17218
rect 12463 17128 12564 17184
rect 12463 17094 12496 17128
rect 12530 17094 12564 17128
rect 12463 17038 12564 17094
rect 12463 17004 12496 17038
rect 12530 17004 12564 17038
rect 12463 16948 12564 17004
rect 12463 16914 12496 16948
rect 12530 16914 12564 16948
rect 12463 16858 12564 16914
rect 12463 16824 12496 16858
rect 12530 16824 12564 16858
rect 12463 16768 12564 16824
rect 12463 16734 12496 16768
rect 12530 16734 12564 16768
rect 12463 16678 12564 16734
rect 12463 16644 12496 16678
rect 12530 16644 12564 16678
rect 12463 16588 12564 16644
rect 12463 16554 12496 16588
rect 12530 16554 12564 16588
rect 12463 16498 12564 16554
rect 12463 16464 12496 16498
rect 12530 16464 12564 16498
rect 12463 16408 12564 16464
rect 12463 16374 12496 16408
rect 12530 16374 12564 16408
rect 12463 16318 12564 16374
rect 11276 16237 11377 16284
rect 12463 16284 12496 16318
rect 12530 16284 12564 16318
rect 12463 16237 12564 16284
rect 11276 16228 12564 16237
rect 11276 16194 11309 16228
rect 11343 16205 12496 16228
rect 11343 16194 11410 16205
rect 11276 16171 11410 16194
rect 11444 16171 11500 16205
rect 11534 16171 11590 16205
rect 11624 16171 11680 16205
rect 11714 16171 11770 16205
rect 11804 16171 11860 16205
rect 11894 16171 11950 16205
rect 11984 16171 12040 16205
rect 12074 16171 12130 16205
rect 12164 16171 12220 16205
rect 12254 16171 12310 16205
rect 12344 16171 12400 16205
rect 12434 16194 12496 16205
rect 12530 16194 12564 16228
rect 12434 16171 12564 16194
rect 11276 16136 12564 16171
rect 12636 17392 13924 17424
rect 12636 17358 12770 17392
rect 12804 17358 12860 17392
rect 12894 17358 12950 17392
rect 12984 17358 13040 17392
rect 13074 17358 13130 17392
rect 13164 17358 13220 17392
rect 13254 17358 13310 17392
rect 13344 17358 13400 17392
rect 13434 17358 13490 17392
rect 13524 17358 13580 17392
rect 13614 17358 13670 17392
rect 13704 17358 13760 17392
rect 13794 17358 13924 17392
rect 12636 17323 13924 17358
rect 12636 17308 12737 17323
rect 12636 17274 12669 17308
rect 12703 17274 12737 17308
rect 12636 17218 12737 17274
rect 13823 17308 13924 17323
rect 13823 17274 13856 17308
rect 13890 17274 13924 17308
rect 12636 17184 12669 17218
rect 12703 17184 12737 17218
rect 12636 17128 12737 17184
rect 12636 17094 12669 17128
rect 12703 17094 12737 17128
rect 12636 17038 12737 17094
rect 12636 17004 12669 17038
rect 12703 17004 12737 17038
rect 12636 16948 12737 17004
rect 12636 16914 12669 16948
rect 12703 16914 12737 16948
rect 12636 16858 12737 16914
rect 12636 16824 12669 16858
rect 12703 16824 12737 16858
rect 12636 16768 12737 16824
rect 12636 16734 12669 16768
rect 12703 16734 12737 16768
rect 12636 16678 12737 16734
rect 12636 16644 12669 16678
rect 12703 16644 12737 16678
rect 12636 16588 12737 16644
rect 12636 16554 12669 16588
rect 12703 16554 12737 16588
rect 12636 16498 12737 16554
rect 12636 16464 12669 16498
rect 12703 16464 12737 16498
rect 12636 16408 12737 16464
rect 12636 16374 12669 16408
rect 12703 16374 12737 16408
rect 12636 16318 12737 16374
rect 12636 16284 12669 16318
rect 12703 16284 12737 16318
rect 13823 17218 13924 17274
rect 13823 17184 13856 17218
rect 13890 17184 13924 17218
rect 13823 17128 13924 17184
rect 13823 17094 13856 17128
rect 13890 17094 13924 17128
rect 13823 17038 13924 17094
rect 13823 17004 13856 17038
rect 13890 17004 13924 17038
rect 13823 16948 13924 17004
rect 13823 16914 13856 16948
rect 13890 16914 13924 16948
rect 13823 16858 13924 16914
rect 13823 16824 13856 16858
rect 13890 16824 13924 16858
rect 13823 16768 13924 16824
rect 13823 16734 13856 16768
rect 13890 16734 13924 16768
rect 13823 16678 13924 16734
rect 13823 16644 13856 16678
rect 13890 16644 13924 16678
rect 13823 16588 13924 16644
rect 13823 16554 13856 16588
rect 13890 16554 13924 16588
rect 13823 16498 13924 16554
rect 13823 16464 13856 16498
rect 13890 16464 13924 16498
rect 13823 16408 13924 16464
rect 13823 16374 13856 16408
rect 13890 16374 13924 16408
rect 13823 16318 13924 16374
rect 12636 16237 12737 16284
rect 13823 16284 13856 16318
rect 13890 16284 13924 16318
rect 13823 16237 13924 16284
rect 12636 16228 13924 16237
rect 12636 16194 12669 16228
rect 12703 16205 13856 16228
rect 12703 16194 12770 16205
rect 12636 16171 12770 16194
rect 12804 16171 12860 16205
rect 12894 16171 12950 16205
rect 12984 16171 13040 16205
rect 13074 16171 13130 16205
rect 13164 16171 13220 16205
rect 13254 16171 13310 16205
rect 13344 16171 13400 16205
rect 13434 16171 13490 16205
rect 13524 16171 13580 16205
rect 13614 16171 13670 16205
rect 13704 16171 13760 16205
rect 13794 16194 13856 16205
rect 13890 16194 13924 16228
rect 13794 16171 13924 16194
rect 12636 16136 13924 16171
rect 13996 17392 15284 17424
rect 13996 17358 14130 17392
rect 14164 17358 14220 17392
rect 14254 17358 14310 17392
rect 14344 17358 14400 17392
rect 14434 17358 14490 17392
rect 14524 17358 14580 17392
rect 14614 17358 14670 17392
rect 14704 17358 14760 17392
rect 14794 17358 14850 17392
rect 14884 17358 14940 17392
rect 14974 17358 15030 17392
rect 15064 17358 15120 17392
rect 15154 17358 15284 17392
rect 13996 17323 15284 17358
rect 13996 17308 14097 17323
rect 13996 17274 14029 17308
rect 14063 17274 14097 17308
rect 13996 17218 14097 17274
rect 15183 17308 15284 17323
rect 15183 17274 15216 17308
rect 15250 17274 15284 17308
rect 13996 17184 14029 17218
rect 14063 17184 14097 17218
rect 13996 17128 14097 17184
rect 13996 17094 14029 17128
rect 14063 17094 14097 17128
rect 13996 17038 14097 17094
rect 13996 17004 14029 17038
rect 14063 17004 14097 17038
rect 13996 16948 14097 17004
rect 13996 16914 14029 16948
rect 14063 16914 14097 16948
rect 13996 16858 14097 16914
rect 13996 16824 14029 16858
rect 14063 16824 14097 16858
rect 13996 16768 14097 16824
rect 13996 16734 14029 16768
rect 14063 16734 14097 16768
rect 13996 16678 14097 16734
rect 13996 16644 14029 16678
rect 14063 16644 14097 16678
rect 13996 16588 14097 16644
rect 13996 16554 14029 16588
rect 14063 16554 14097 16588
rect 13996 16498 14097 16554
rect 13996 16464 14029 16498
rect 14063 16464 14097 16498
rect 13996 16408 14097 16464
rect 13996 16374 14029 16408
rect 14063 16374 14097 16408
rect 13996 16318 14097 16374
rect 13996 16284 14029 16318
rect 14063 16284 14097 16318
rect 15183 17218 15284 17274
rect 15183 17184 15216 17218
rect 15250 17184 15284 17218
rect 15183 17128 15284 17184
rect 15183 17094 15216 17128
rect 15250 17094 15284 17128
rect 15183 17038 15284 17094
rect 15183 17004 15216 17038
rect 15250 17004 15284 17038
rect 15183 16948 15284 17004
rect 15183 16914 15216 16948
rect 15250 16914 15284 16948
rect 15183 16858 15284 16914
rect 15183 16824 15216 16858
rect 15250 16824 15284 16858
rect 15183 16768 15284 16824
rect 15183 16734 15216 16768
rect 15250 16734 15284 16768
rect 15183 16678 15284 16734
rect 15183 16644 15216 16678
rect 15250 16644 15284 16678
rect 15183 16588 15284 16644
rect 15183 16554 15216 16588
rect 15250 16554 15284 16588
rect 15183 16498 15284 16554
rect 15183 16464 15216 16498
rect 15250 16464 15284 16498
rect 15183 16408 15284 16464
rect 15183 16374 15216 16408
rect 15250 16374 15284 16408
rect 15183 16318 15284 16374
rect 13996 16237 14097 16284
rect 15183 16284 15216 16318
rect 15250 16284 15284 16318
rect 15183 16237 15284 16284
rect 13996 16228 15284 16237
rect 13996 16194 14029 16228
rect 14063 16205 15216 16228
rect 14063 16194 14130 16205
rect 13996 16171 14130 16194
rect 14164 16171 14220 16205
rect 14254 16171 14310 16205
rect 14344 16171 14400 16205
rect 14434 16171 14490 16205
rect 14524 16171 14580 16205
rect 14614 16171 14670 16205
rect 14704 16171 14760 16205
rect 14794 16171 14850 16205
rect 14884 16171 14940 16205
rect 14974 16171 15030 16205
rect 15064 16171 15120 16205
rect 15154 16194 15216 16205
rect 15250 16194 15284 16228
rect 15154 16171 15284 16194
rect 13996 16136 15284 16171
rect 11276 16032 12564 16064
rect 11276 15998 11410 16032
rect 11444 15998 11500 16032
rect 11534 15998 11590 16032
rect 11624 15998 11680 16032
rect 11714 15998 11770 16032
rect 11804 15998 11860 16032
rect 11894 15998 11950 16032
rect 11984 15998 12040 16032
rect 12074 15998 12130 16032
rect 12164 15998 12220 16032
rect 12254 15998 12310 16032
rect 12344 15998 12400 16032
rect 12434 15998 12564 16032
rect 11276 15963 12564 15998
rect 11276 15948 11377 15963
rect 11276 15914 11309 15948
rect 11343 15914 11377 15948
rect 11276 15858 11377 15914
rect 12463 15948 12564 15963
rect 12463 15914 12496 15948
rect 12530 15914 12564 15948
rect 11276 15824 11309 15858
rect 11343 15824 11377 15858
rect 11276 15768 11377 15824
rect 11276 15734 11309 15768
rect 11343 15734 11377 15768
rect 11276 15678 11377 15734
rect 11276 15644 11309 15678
rect 11343 15644 11377 15678
rect 11276 15588 11377 15644
rect 11276 15554 11309 15588
rect 11343 15554 11377 15588
rect 11276 15498 11377 15554
rect 11276 15464 11309 15498
rect 11343 15464 11377 15498
rect 11276 15408 11377 15464
rect 11276 15374 11309 15408
rect 11343 15374 11377 15408
rect 11276 15318 11377 15374
rect 11276 15284 11309 15318
rect 11343 15284 11377 15318
rect 11276 15228 11377 15284
rect 11276 15194 11309 15228
rect 11343 15194 11377 15228
rect 11276 15138 11377 15194
rect 11276 15104 11309 15138
rect 11343 15104 11377 15138
rect 11276 15048 11377 15104
rect 11276 15014 11309 15048
rect 11343 15014 11377 15048
rect 11276 14958 11377 15014
rect 11276 14924 11309 14958
rect 11343 14924 11377 14958
rect 12463 15858 12564 15914
rect 12463 15824 12496 15858
rect 12530 15824 12564 15858
rect 12463 15768 12564 15824
rect 12463 15734 12496 15768
rect 12530 15734 12564 15768
rect 12463 15678 12564 15734
rect 12463 15644 12496 15678
rect 12530 15644 12564 15678
rect 12463 15588 12564 15644
rect 12463 15554 12496 15588
rect 12530 15554 12564 15588
rect 12463 15498 12564 15554
rect 12463 15464 12496 15498
rect 12530 15464 12564 15498
rect 12463 15408 12564 15464
rect 12463 15374 12496 15408
rect 12530 15374 12564 15408
rect 12463 15318 12564 15374
rect 12463 15284 12496 15318
rect 12530 15284 12564 15318
rect 12463 15228 12564 15284
rect 12463 15194 12496 15228
rect 12530 15194 12564 15228
rect 12463 15138 12564 15194
rect 12463 15104 12496 15138
rect 12530 15104 12564 15138
rect 12463 15048 12564 15104
rect 12463 15014 12496 15048
rect 12530 15014 12564 15048
rect 12463 14958 12564 15014
rect 11276 14877 11377 14924
rect 12463 14924 12496 14958
rect 12530 14924 12564 14958
rect 12463 14877 12564 14924
rect 11276 14868 12564 14877
rect 11276 14834 11309 14868
rect 11343 14845 12496 14868
rect 11343 14834 11410 14845
rect 11276 14811 11410 14834
rect 11444 14811 11500 14845
rect 11534 14811 11590 14845
rect 11624 14811 11680 14845
rect 11714 14811 11770 14845
rect 11804 14811 11860 14845
rect 11894 14811 11950 14845
rect 11984 14811 12040 14845
rect 12074 14811 12130 14845
rect 12164 14811 12220 14845
rect 12254 14811 12310 14845
rect 12344 14811 12400 14845
rect 12434 14834 12496 14845
rect 12530 14834 12564 14868
rect 12434 14811 12564 14834
rect 11276 14776 12564 14811
rect 12636 16032 13924 16064
rect 12636 15998 12770 16032
rect 12804 15998 12860 16032
rect 12894 15998 12950 16032
rect 12984 15998 13040 16032
rect 13074 15998 13130 16032
rect 13164 15998 13220 16032
rect 13254 15998 13310 16032
rect 13344 15998 13400 16032
rect 13434 15998 13490 16032
rect 13524 15998 13580 16032
rect 13614 15998 13670 16032
rect 13704 15998 13760 16032
rect 13794 15998 13924 16032
rect 12636 15963 13924 15998
rect 12636 15948 12737 15963
rect 12636 15914 12669 15948
rect 12703 15914 12737 15948
rect 12636 15858 12737 15914
rect 13823 15948 13924 15963
rect 13823 15914 13856 15948
rect 13890 15914 13924 15948
rect 12636 15824 12669 15858
rect 12703 15824 12737 15858
rect 12636 15768 12737 15824
rect 12636 15734 12669 15768
rect 12703 15734 12737 15768
rect 12636 15678 12737 15734
rect 12636 15644 12669 15678
rect 12703 15644 12737 15678
rect 12636 15588 12737 15644
rect 12636 15554 12669 15588
rect 12703 15554 12737 15588
rect 12636 15498 12737 15554
rect 12636 15464 12669 15498
rect 12703 15464 12737 15498
rect 12636 15408 12737 15464
rect 12636 15374 12669 15408
rect 12703 15374 12737 15408
rect 12636 15318 12737 15374
rect 12636 15284 12669 15318
rect 12703 15284 12737 15318
rect 12636 15228 12737 15284
rect 12636 15194 12669 15228
rect 12703 15194 12737 15228
rect 12636 15138 12737 15194
rect 12636 15104 12669 15138
rect 12703 15104 12737 15138
rect 12636 15048 12737 15104
rect 12636 15014 12669 15048
rect 12703 15014 12737 15048
rect 12636 14958 12737 15014
rect 12636 14924 12669 14958
rect 12703 14924 12737 14958
rect 13823 15858 13924 15914
rect 13823 15824 13856 15858
rect 13890 15824 13924 15858
rect 13823 15768 13924 15824
rect 13823 15734 13856 15768
rect 13890 15734 13924 15768
rect 13823 15678 13924 15734
rect 13823 15644 13856 15678
rect 13890 15644 13924 15678
rect 13823 15588 13924 15644
rect 13823 15554 13856 15588
rect 13890 15554 13924 15588
rect 13823 15498 13924 15554
rect 13823 15464 13856 15498
rect 13890 15464 13924 15498
rect 13823 15408 13924 15464
rect 13823 15374 13856 15408
rect 13890 15374 13924 15408
rect 13823 15318 13924 15374
rect 13823 15284 13856 15318
rect 13890 15284 13924 15318
rect 13823 15228 13924 15284
rect 13823 15194 13856 15228
rect 13890 15194 13924 15228
rect 13823 15138 13924 15194
rect 13823 15104 13856 15138
rect 13890 15104 13924 15138
rect 13823 15048 13924 15104
rect 13823 15014 13856 15048
rect 13890 15014 13924 15048
rect 13823 14958 13924 15014
rect 12636 14877 12737 14924
rect 13823 14924 13856 14958
rect 13890 14924 13924 14958
rect 13823 14877 13924 14924
rect 12636 14868 13924 14877
rect 12636 14834 12669 14868
rect 12703 14845 13856 14868
rect 12703 14834 12770 14845
rect 12636 14811 12770 14834
rect 12804 14811 12860 14845
rect 12894 14811 12950 14845
rect 12984 14811 13040 14845
rect 13074 14811 13130 14845
rect 13164 14811 13220 14845
rect 13254 14811 13310 14845
rect 13344 14811 13400 14845
rect 13434 14811 13490 14845
rect 13524 14811 13580 14845
rect 13614 14811 13670 14845
rect 13704 14811 13760 14845
rect 13794 14834 13856 14845
rect 13890 14834 13924 14868
rect 13794 14811 13924 14834
rect 12636 14776 13924 14811
rect 13996 16032 15284 16064
rect 13996 15998 14130 16032
rect 14164 15998 14220 16032
rect 14254 15998 14310 16032
rect 14344 15998 14400 16032
rect 14434 15998 14490 16032
rect 14524 15998 14580 16032
rect 14614 15998 14670 16032
rect 14704 15998 14760 16032
rect 14794 15998 14850 16032
rect 14884 15998 14940 16032
rect 14974 15998 15030 16032
rect 15064 15998 15120 16032
rect 15154 15998 15284 16032
rect 13996 15963 15284 15998
rect 13996 15948 14097 15963
rect 13996 15914 14029 15948
rect 14063 15914 14097 15948
rect 13996 15858 14097 15914
rect 15183 15948 15284 15963
rect 15183 15914 15216 15948
rect 15250 15914 15284 15948
rect 13996 15824 14029 15858
rect 14063 15824 14097 15858
rect 13996 15768 14097 15824
rect 13996 15734 14029 15768
rect 14063 15734 14097 15768
rect 13996 15678 14097 15734
rect 13996 15644 14029 15678
rect 14063 15644 14097 15678
rect 13996 15588 14097 15644
rect 13996 15554 14029 15588
rect 14063 15554 14097 15588
rect 13996 15498 14097 15554
rect 13996 15464 14029 15498
rect 14063 15464 14097 15498
rect 13996 15408 14097 15464
rect 13996 15374 14029 15408
rect 14063 15374 14097 15408
rect 13996 15318 14097 15374
rect 13996 15284 14029 15318
rect 14063 15284 14097 15318
rect 13996 15228 14097 15284
rect 13996 15194 14029 15228
rect 14063 15194 14097 15228
rect 13996 15138 14097 15194
rect 13996 15104 14029 15138
rect 14063 15104 14097 15138
rect 13996 15048 14097 15104
rect 13996 15014 14029 15048
rect 14063 15014 14097 15048
rect 13996 14958 14097 15014
rect 13996 14924 14029 14958
rect 14063 14924 14097 14958
rect 15183 15858 15284 15914
rect 15183 15824 15216 15858
rect 15250 15824 15284 15858
rect 15183 15768 15284 15824
rect 15183 15734 15216 15768
rect 15250 15734 15284 15768
rect 15183 15678 15284 15734
rect 15183 15644 15216 15678
rect 15250 15644 15284 15678
rect 15183 15588 15284 15644
rect 15183 15554 15216 15588
rect 15250 15554 15284 15588
rect 15183 15498 15284 15554
rect 15183 15464 15216 15498
rect 15250 15464 15284 15498
rect 15183 15408 15284 15464
rect 15183 15374 15216 15408
rect 15250 15374 15284 15408
rect 15183 15318 15284 15374
rect 15183 15284 15216 15318
rect 15250 15284 15284 15318
rect 15183 15228 15284 15284
rect 15183 15194 15216 15228
rect 15250 15194 15284 15228
rect 15183 15138 15284 15194
rect 15183 15104 15216 15138
rect 15250 15104 15284 15138
rect 15183 15048 15284 15104
rect 15183 15014 15216 15048
rect 15250 15014 15284 15048
rect 15183 14958 15284 15014
rect 13996 14877 14097 14924
rect 15183 14924 15216 14958
rect 15250 14924 15284 14958
rect 15183 14877 15284 14924
rect 13996 14868 15284 14877
rect 13996 14834 14029 14868
rect 14063 14845 15216 14868
rect 14063 14834 14130 14845
rect 13996 14811 14130 14834
rect 14164 14811 14220 14845
rect 14254 14811 14310 14845
rect 14344 14811 14400 14845
rect 14434 14811 14490 14845
rect 14524 14811 14580 14845
rect 14614 14811 14670 14845
rect 14704 14811 14760 14845
rect 14794 14811 14850 14845
rect 14884 14811 14940 14845
rect 14974 14811 15030 14845
rect 15064 14811 15120 14845
rect 15154 14834 15216 14845
rect 15250 14834 15284 14868
rect 15154 14811 15284 14834
rect 13996 14776 15284 14811
rect 15400 13850 15480 13880
rect 15400 13810 15420 13850
rect 15460 13810 15480 13850
rect 15400 13750 15480 13810
rect 15400 13710 15420 13750
rect 15460 13710 15480 13750
rect 15400 13680 15480 13710
rect 11900 13240 11980 13270
rect 11900 13200 11920 13240
rect 11960 13200 11980 13240
rect 11900 13140 11980 13200
rect 11900 13100 11920 13140
rect 11960 13100 11980 13140
rect 11900 13040 11980 13100
rect 11900 13000 11920 13040
rect 11960 13000 11980 13040
rect 11900 12940 11980 13000
rect 11900 12900 11920 12940
rect 11960 12900 11980 12940
rect 11900 12840 11980 12900
rect 11900 12800 11920 12840
rect 11960 12800 11980 12840
rect 11900 12770 11980 12800
rect 14580 13240 14660 13270
rect 14580 13200 14600 13240
rect 14640 13200 14660 13240
rect 14580 13140 14660 13200
rect 14580 13100 14600 13140
rect 14640 13100 14660 13140
rect 14580 13040 14660 13100
rect 14580 13000 14600 13040
rect 14640 13000 14660 13040
rect 14580 12940 14660 13000
rect 14580 12900 14600 12940
rect 14640 12900 14660 12940
rect 14580 12840 14660 12900
rect 14580 12800 14600 12840
rect 14640 12800 14660 12840
rect 14580 12770 14660 12800
rect 12800 12320 12880 12350
rect 12800 12280 12820 12320
rect 12860 12280 12880 12320
rect 12800 12240 12880 12280
rect 12800 12200 12820 12240
rect 12860 12200 12880 12240
rect 12800 12160 12880 12200
rect 12800 12120 12820 12160
rect 12860 12120 12880 12160
rect 12800 12090 12880 12120
rect 13680 12320 13760 12350
rect 13680 12280 13700 12320
rect 13740 12280 13760 12320
rect 13680 12240 13760 12280
rect 13680 12200 13700 12240
rect 13740 12200 13760 12240
rect 13680 12160 13760 12200
rect 13680 12120 13700 12160
rect 13740 12120 13760 12160
rect 13680 12090 13760 12120
<< nsubdiff >>
rect 8603 18555 8699 18589
rect 8959 18555 9055 18589
rect 8603 18493 8637 18555
rect 9021 18493 9055 18555
rect 8603 16527 8637 16589
rect 9021 16527 9055 16589
rect 8603 16493 8699 16527
rect 8959 16493 9055 16527
rect 9383 18561 9479 18595
rect 9739 18561 9835 18595
rect 9383 18499 9417 18561
rect 9801 18499 9835 18561
rect 9383 14957 9417 15019
rect 10163 18563 10259 18597
rect 10851 18563 10947 18597
rect 10163 18501 10197 18563
rect 10913 18501 10947 18563
rect 10163 16181 10197 16243
rect 11439 18602 12401 18621
rect 11439 18568 11550 18602
rect 11584 18568 11640 18602
rect 11674 18568 11730 18602
rect 11764 18568 11820 18602
rect 11854 18568 11910 18602
rect 11944 18568 12000 18602
rect 12034 18568 12090 18602
rect 12124 18568 12180 18602
rect 12214 18568 12270 18602
rect 12304 18568 12401 18602
rect 11439 18549 12401 18568
rect 11439 18508 11511 18549
rect 11439 18474 11458 18508
rect 11492 18474 11511 18508
rect 12329 18489 12401 18549
rect 11439 18418 11511 18474
rect 11439 18384 11458 18418
rect 11492 18384 11511 18418
rect 11439 18328 11511 18384
rect 11439 18294 11458 18328
rect 11492 18294 11511 18328
rect 11439 18238 11511 18294
rect 11439 18204 11458 18238
rect 11492 18204 11511 18238
rect 11439 18148 11511 18204
rect 11439 18114 11458 18148
rect 11492 18114 11511 18148
rect 11439 18058 11511 18114
rect 11439 18024 11458 18058
rect 11492 18024 11511 18058
rect 11439 17968 11511 18024
rect 11439 17934 11458 17968
rect 11492 17934 11511 17968
rect 11439 17878 11511 17934
rect 11439 17844 11458 17878
rect 11492 17844 11511 17878
rect 11439 17788 11511 17844
rect 12329 18455 12348 18489
rect 12382 18455 12401 18489
rect 12329 18399 12401 18455
rect 12329 18365 12348 18399
rect 12382 18365 12401 18399
rect 12329 18309 12401 18365
rect 12329 18275 12348 18309
rect 12382 18275 12401 18309
rect 12329 18219 12401 18275
rect 12329 18185 12348 18219
rect 12382 18185 12401 18219
rect 12329 18129 12401 18185
rect 12329 18095 12348 18129
rect 12382 18095 12401 18129
rect 12329 18039 12401 18095
rect 12329 18005 12348 18039
rect 12382 18005 12401 18039
rect 12329 17949 12401 18005
rect 12329 17915 12348 17949
rect 12382 17915 12401 17949
rect 12329 17859 12401 17915
rect 12329 17825 12348 17859
rect 12382 17825 12401 17859
rect 11439 17754 11458 17788
rect 11492 17754 11511 17788
rect 11439 17731 11511 17754
rect 12329 17769 12401 17825
rect 12329 17735 12348 17769
rect 12382 17735 12401 17769
rect 12329 17731 12401 17735
rect 11439 17712 12401 17731
rect 11439 17678 11516 17712
rect 11550 17678 11606 17712
rect 11640 17678 11696 17712
rect 11730 17678 11786 17712
rect 11820 17678 11876 17712
rect 11910 17678 11966 17712
rect 12000 17678 12056 17712
rect 12090 17678 12146 17712
rect 12180 17678 12236 17712
rect 12270 17678 12401 17712
rect 11439 17659 12401 17678
rect 12799 18602 13761 18621
rect 12799 18568 12910 18602
rect 12944 18568 13000 18602
rect 13034 18568 13090 18602
rect 13124 18568 13180 18602
rect 13214 18568 13270 18602
rect 13304 18568 13360 18602
rect 13394 18568 13450 18602
rect 13484 18568 13540 18602
rect 13574 18568 13630 18602
rect 13664 18568 13761 18602
rect 12799 18549 13761 18568
rect 12799 18508 12871 18549
rect 12799 18474 12818 18508
rect 12852 18474 12871 18508
rect 13689 18489 13761 18549
rect 12799 18418 12871 18474
rect 12799 18384 12818 18418
rect 12852 18384 12871 18418
rect 12799 18328 12871 18384
rect 12799 18294 12818 18328
rect 12852 18294 12871 18328
rect 12799 18238 12871 18294
rect 12799 18204 12818 18238
rect 12852 18204 12871 18238
rect 12799 18148 12871 18204
rect 12799 18114 12818 18148
rect 12852 18114 12871 18148
rect 12799 18058 12871 18114
rect 12799 18024 12818 18058
rect 12852 18024 12871 18058
rect 12799 17968 12871 18024
rect 12799 17934 12818 17968
rect 12852 17934 12871 17968
rect 12799 17878 12871 17934
rect 12799 17844 12818 17878
rect 12852 17844 12871 17878
rect 12799 17788 12871 17844
rect 13689 18455 13708 18489
rect 13742 18455 13761 18489
rect 13689 18399 13761 18455
rect 13689 18365 13708 18399
rect 13742 18365 13761 18399
rect 13689 18309 13761 18365
rect 13689 18275 13708 18309
rect 13742 18275 13761 18309
rect 13689 18219 13761 18275
rect 13689 18185 13708 18219
rect 13742 18185 13761 18219
rect 13689 18129 13761 18185
rect 13689 18095 13708 18129
rect 13742 18095 13761 18129
rect 13689 18039 13761 18095
rect 13689 18005 13708 18039
rect 13742 18005 13761 18039
rect 13689 17949 13761 18005
rect 13689 17915 13708 17949
rect 13742 17915 13761 17949
rect 13689 17859 13761 17915
rect 13689 17825 13708 17859
rect 13742 17825 13761 17859
rect 12799 17754 12818 17788
rect 12852 17754 12871 17788
rect 12799 17731 12871 17754
rect 13689 17769 13761 17825
rect 13689 17735 13708 17769
rect 13742 17735 13761 17769
rect 13689 17731 13761 17735
rect 12799 17712 13761 17731
rect 12799 17678 12876 17712
rect 12910 17678 12966 17712
rect 13000 17678 13056 17712
rect 13090 17678 13146 17712
rect 13180 17678 13236 17712
rect 13270 17678 13326 17712
rect 13360 17678 13416 17712
rect 13450 17678 13506 17712
rect 13540 17678 13596 17712
rect 13630 17678 13761 17712
rect 12799 17659 13761 17678
rect 14159 18602 15121 18621
rect 14159 18568 14270 18602
rect 14304 18568 14360 18602
rect 14394 18568 14450 18602
rect 14484 18568 14540 18602
rect 14574 18568 14630 18602
rect 14664 18568 14720 18602
rect 14754 18568 14810 18602
rect 14844 18568 14900 18602
rect 14934 18568 14990 18602
rect 15024 18568 15121 18602
rect 14159 18549 15121 18568
rect 14159 18508 14231 18549
rect 14159 18474 14178 18508
rect 14212 18474 14231 18508
rect 15049 18489 15121 18549
rect 14159 18418 14231 18474
rect 14159 18384 14178 18418
rect 14212 18384 14231 18418
rect 14159 18328 14231 18384
rect 14159 18294 14178 18328
rect 14212 18294 14231 18328
rect 14159 18238 14231 18294
rect 14159 18204 14178 18238
rect 14212 18204 14231 18238
rect 14159 18148 14231 18204
rect 14159 18114 14178 18148
rect 14212 18114 14231 18148
rect 14159 18058 14231 18114
rect 14159 18024 14178 18058
rect 14212 18024 14231 18058
rect 14159 17968 14231 18024
rect 14159 17934 14178 17968
rect 14212 17934 14231 17968
rect 14159 17878 14231 17934
rect 14159 17844 14178 17878
rect 14212 17844 14231 17878
rect 14159 17788 14231 17844
rect 15049 18455 15068 18489
rect 15102 18455 15121 18489
rect 15049 18399 15121 18455
rect 15049 18365 15068 18399
rect 15102 18365 15121 18399
rect 15049 18309 15121 18365
rect 15049 18275 15068 18309
rect 15102 18275 15121 18309
rect 15049 18219 15121 18275
rect 15049 18185 15068 18219
rect 15102 18185 15121 18219
rect 15049 18129 15121 18185
rect 15049 18095 15068 18129
rect 15102 18095 15121 18129
rect 15049 18039 15121 18095
rect 15049 18005 15068 18039
rect 15102 18005 15121 18039
rect 15049 17949 15121 18005
rect 15049 17915 15068 17949
rect 15102 17915 15121 17949
rect 15049 17859 15121 17915
rect 15049 17825 15068 17859
rect 15102 17825 15121 17859
rect 14159 17754 14178 17788
rect 14212 17754 14231 17788
rect 14159 17731 14231 17754
rect 15049 17769 15121 17825
rect 15049 17735 15068 17769
rect 15102 17735 15121 17769
rect 15049 17731 15121 17735
rect 14159 17712 15121 17731
rect 14159 17678 14236 17712
rect 14270 17678 14326 17712
rect 14360 17678 14416 17712
rect 14450 17678 14506 17712
rect 14540 17678 14596 17712
rect 14630 17678 14686 17712
rect 14720 17678 14776 17712
rect 14810 17678 14866 17712
rect 14900 17678 14956 17712
rect 14990 17678 15121 17712
rect 14159 17659 15121 17678
rect 15483 18563 15579 18597
rect 16171 18563 16267 18597
rect 15483 18501 15517 18563
rect 10913 16181 10947 16243
rect 10163 16147 10259 16181
rect 10851 16147 10947 16181
rect 11439 17242 12401 17261
rect 11439 17208 11550 17242
rect 11584 17208 11640 17242
rect 11674 17208 11730 17242
rect 11764 17208 11820 17242
rect 11854 17208 11910 17242
rect 11944 17208 12000 17242
rect 12034 17208 12090 17242
rect 12124 17208 12180 17242
rect 12214 17208 12270 17242
rect 12304 17208 12401 17242
rect 11439 17189 12401 17208
rect 11439 17148 11511 17189
rect 11439 17114 11458 17148
rect 11492 17114 11511 17148
rect 12329 17129 12401 17189
rect 11439 17058 11511 17114
rect 11439 17024 11458 17058
rect 11492 17024 11511 17058
rect 11439 16968 11511 17024
rect 11439 16934 11458 16968
rect 11492 16934 11511 16968
rect 11439 16878 11511 16934
rect 11439 16844 11458 16878
rect 11492 16844 11511 16878
rect 11439 16788 11511 16844
rect 11439 16754 11458 16788
rect 11492 16754 11511 16788
rect 11439 16698 11511 16754
rect 11439 16664 11458 16698
rect 11492 16664 11511 16698
rect 11439 16608 11511 16664
rect 11439 16574 11458 16608
rect 11492 16574 11511 16608
rect 11439 16518 11511 16574
rect 11439 16484 11458 16518
rect 11492 16484 11511 16518
rect 11439 16428 11511 16484
rect 12329 17095 12348 17129
rect 12382 17095 12401 17129
rect 12329 17039 12401 17095
rect 12329 17005 12348 17039
rect 12382 17005 12401 17039
rect 12329 16949 12401 17005
rect 12329 16915 12348 16949
rect 12382 16915 12401 16949
rect 12329 16859 12401 16915
rect 12329 16825 12348 16859
rect 12382 16825 12401 16859
rect 12329 16769 12401 16825
rect 12329 16735 12348 16769
rect 12382 16735 12401 16769
rect 12329 16679 12401 16735
rect 12329 16645 12348 16679
rect 12382 16645 12401 16679
rect 12329 16589 12401 16645
rect 12329 16555 12348 16589
rect 12382 16555 12401 16589
rect 12329 16499 12401 16555
rect 12329 16465 12348 16499
rect 12382 16465 12401 16499
rect 11439 16394 11458 16428
rect 11492 16394 11511 16428
rect 11439 16371 11511 16394
rect 12329 16409 12401 16465
rect 12329 16375 12348 16409
rect 12382 16375 12401 16409
rect 12329 16371 12401 16375
rect 11439 16352 12401 16371
rect 11439 16318 11516 16352
rect 11550 16318 11606 16352
rect 11640 16318 11696 16352
rect 11730 16318 11786 16352
rect 11820 16318 11876 16352
rect 11910 16318 11966 16352
rect 12000 16318 12056 16352
rect 12090 16318 12146 16352
rect 12180 16318 12236 16352
rect 12270 16318 12401 16352
rect 11439 16299 12401 16318
rect 12799 17242 13761 17261
rect 12799 17208 12910 17242
rect 12944 17208 13000 17242
rect 13034 17208 13090 17242
rect 13124 17208 13180 17242
rect 13214 17208 13270 17242
rect 13304 17208 13360 17242
rect 13394 17208 13450 17242
rect 13484 17208 13540 17242
rect 13574 17208 13630 17242
rect 13664 17208 13761 17242
rect 12799 17189 13761 17208
rect 12799 17148 12871 17189
rect 12799 17114 12818 17148
rect 12852 17114 12871 17148
rect 13689 17129 13761 17189
rect 12799 17058 12871 17114
rect 12799 17024 12818 17058
rect 12852 17024 12871 17058
rect 12799 16968 12871 17024
rect 12799 16934 12818 16968
rect 12852 16934 12871 16968
rect 12799 16878 12871 16934
rect 12799 16844 12818 16878
rect 12852 16844 12871 16878
rect 12799 16788 12871 16844
rect 12799 16754 12818 16788
rect 12852 16754 12871 16788
rect 12799 16698 12871 16754
rect 12799 16664 12818 16698
rect 12852 16664 12871 16698
rect 12799 16608 12871 16664
rect 12799 16574 12818 16608
rect 12852 16574 12871 16608
rect 12799 16518 12871 16574
rect 12799 16484 12818 16518
rect 12852 16484 12871 16518
rect 12799 16428 12871 16484
rect 13689 17095 13708 17129
rect 13742 17095 13761 17129
rect 13689 17039 13761 17095
rect 13689 17005 13708 17039
rect 13742 17005 13761 17039
rect 13689 16949 13761 17005
rect 13689 16915 13708 16949
rect 13742 16915 13761 16949
rect 13689 16859 13761 16915
rect 13689 16825 13708 16859
rect 13742 16825 13761 16859
rect 13689 16769 13761 16825
rect 13689 16735 13708 16769
rect 13742 16735 13761 16769
rect 13689 16679 13761 16735
rect 13689 16645 13708 16679
rect 13742 16645 13761 16679
rect 13689 16589 13761 16645
rect 13689 16555 13708 16589
rect 13742 16555 13761 16589
rect 13689 16499 13761 16555
rect 13689 16465 13708 16499
rect 13742 16465 13761 16499
rect 12799 16394 12818 16428
rect 12852 16394 12871 16428
rect 12799 16371 12871 16394
rect 13689 16409 13761 16465
rect 13689 16375 13708 16409
rect 13742 16375 13761 16409
rect 13689 16371 13761 16375
rect 12799 16352 13761 16371
rect 12799 16318 12876 16352
rect 12910 16318 12966 16352
rect 13000 16318 13056 16352
rect 13090 16318 13146 16352
rect 13180 16318 13236 16352
rect 13270 16318 13326 16352
rect 13360 16318 13416 16352
rect 13450 16318 13506 16352
rect 13540 16318 13596 16352
rect 13630 16318 13761 16352
rect 12799 16299 13761 16318
rect 14159 17242 15121 17261
rect 14159 17208 14270 17242
rect 14304 17208 14360 17242
rect 14394 17208 14450 17242
rect 14484 17208 14540 17242
rect 14574 17208 14630 17242
rect 14664 17208 14720 17242
rect 14754 17208 14810 17242
rect 14844 17208 14900 17242
rect 14934 17208 14990 17242
rect 15024 17208 15121 17242
rect 14159 17189 15121 17208
rect 14159 17148 14231 17189
rect 14159 17114 14178 17148
rect 14212 17114 14231 17148
rect 15049 17129 15121 17189
rect 14159 17058 14231 17114
rect 14159 17024 14178 17058
rect 14212 17024 14231 17058
rect 14159 16968 14231 17024
rect 14159 16934 14178 16968
rect 14212 16934 14231 16968
rect 14159 16878 14231 16934
rect 14159 16844 14178 16878
rect 14212 16844 14231 16878
rect 14159 16788 14231 16844
rect 14159 16754 14178 16788
rect 14212 16754 14231 16788
rect 14159 16698 14231 16754
rect 14159 16664 14178 16698
rect 14212 16664 14231 16698
rect 14159 16608 14231 16664
rect 14159 16574 14178 16608
rect 14212 16574 14231 16608
rect 14159 16518 14231 16574
rect 14159 16484 14178 16518
rect 14212 16484 14231 16518
rect 14159 16428 14231 16484
rect 15049 17095 15068 17129
rect 15102 17095 15121 17129
rect 15049 17039 15121 17095
rect 15049 17005 15068 17039
rect 15102 17005 15121 17039
rect 15049 16949 15121 17005
rect 15049 16915 15068 16949
rect 15102 16915 15121 16949
rect 15049 16859 15121 16915
rect 15049 16825 15068 16859
rect 15102 16825 15121 16859
rect 15049 16769 15121 16825
rect 15049 16735 15068 16769
rect 15102 16735 15121 16769
rect 15049 16679 15121 16735
rect 15049 16645 15068 16679
rect 15102 16645 15121 16679
rect 15049 16589 15121 16645
rect 15049 16555 15068 16589
rect 15102 16555 15121 16589
rect 15049 16499 15121 16555
rect 15049 16465 15068 16499
rect 15102 16465 15121 16499
rect 14159 16394 14178 16428
rect 14212 16394 14231 16428
rect 14159 16371 14231 16394
rect 15049 16409 15121 16465
rect 15049 16375 15068 16409
rect 15102 16375 15121 16409
rect 15049 16371 15121 16375
rect 14159 16352 15121 16371
rect 14159 16318 14236 16352
rect 14270 16318 14326 16352
rect 14360 16318 14416 16352
rect 14450 16318 14506 16352
rect 14540 16318 14596 16352
rect 14630 16318 14686 16352
rect 14720 16318 14776 16352
rect 14810 16318 14866 16352
rect 14900 16318 14956 16352
rect 14990 16318 15121 16352
rect 14159 16299 15121 16318
rect 16233 18501 16267 18563
rect 15483 16181 15517 16243
rect 16233 16181 16267 16243
rect 15483 16147 15579 16181
rect 16171 16147 16267 16181
rect 16593 18561 16689 18595
rect 16949 18561 17045 18595
rect 16593 18499 16627 18561
rect 9801 14957 9835 15019
rect 9383 14923 9479 14957
rect 9739 14923 9835 14957
rect 11439 15882 12401 15901
rect 11439 15848 11550 15882
rect 11584 15848 11640 15882
rect 11674 15848 11730 15882
rect 11764 15848 11820 15882
rect 11854 15848 11910 15882
rect 11944 15848 12000 15882
rect 12034 15848 12090 15882
rect 12124 15848 12180 15882
rect 12214 15848 12270 15882
rect 12304 15848 12401 15882
rect 11439 15829 12401 15848
rect 11439 15788 11511 15829
rect 11439 15754 11458 15788
rect 11492 15754 11511 15788
rect 12329 15769 12401 15829
rect 11439 15698 11511 15754
rect 11439 15664 11458 15698
rect 11492 15664 11511 15698
rect 11439 15608 11511 15664
rect 11439 15574 11458 15608
rect 11492 15574 11511 15608
rect 11439 15518 11511 15574
rect 11439 15484 11458 15518
rect 11492 15484 11511 15518
rect 11439 15428 11511 15484
rect 11439 15394 11458 15428
rect 11492 15394 11511 15428
rect 11439 15338 11511 15394
rect 11439 15304 11458 15338
rect 11492 15304 11511 15338
rect 11439 15248 11511 15304
rect 11439 15214 11458 15248
rect 11492 15214 11511 15248
rect 11439 15158 11511 15214
rect 11439 15124 11458 15158
rect 11492 15124 11511 15158
rect 11439 15068 11511 15124
rect 12329 15735 12348 15769
rect 12382 15735 12401 15769
rect 12329 15679 12401 15735
rect 12329 15645 12348 15679
rect 12382 15645 12401 15679
rect 12329 15589 12401 15645
rect 12329 15555 12348 15589
rect 12382 15555 12401 15589
rect 12329 15499 12401 15555
rect 12329 15465 12348 15499
rect 12382 15465 12401 15499
rect 12329 15409 12401 15465
rect 12329 15375 12348 15409
rect 12382 15375 12401 15409
rect 12329 15319 12401 15375
rect 12329 15285 12348 15319
rect 12382 15285 12401 15319
rect 12329 15229 12401 15285
rect 12329 15195 12348 15229
rect 12382 15195 12401 15229
rect 12329 15139 12401 15195
rect 12329 15105 12348 15139
rect 12382 15105 12401 15139
rect 11439 15034 11458 15068
rect 11492 15034 11511 15068
rect 11439 15011 11511 15034
rect 12329 15049 12401 15105
rect 12329 15015 12348 15049
rect 12382 15015 12401 15049
rect 12329 15011 12401 15015
rect 11439 14992 12401 15011
rect 11439 14958 11516 14992
rect 11550 14958 11606 14992
rect 11640 14958 11696 14992
rect 11730 14958 11786 14992
rect 11820 14958 11876 14992
rect 11910 14958 11966 14992
rect 12000 14958 12056 14992
rect 12090 14958 12146 14992
rect 12180 14958 12236 14992
rect 12270 14958 12401 14992
rect 11439 14939 12401 14958
rect 12799 15882 13761 15901
rect 12799 15848 12910 15882
rect 12944 15848 13000 15882
rect 13034 15848 13090 15882
rect 13124 15848 13180 15882
rect 13214 15848 13270 15882
rect 13304 15848 13360 15882
rect 13394 15848 13450 15882
rect 13484 15848 13540 15882
rect 13574 15848 13630 15882
rect 13664 15848 13761 15882
rect 12799 15829 13761 15848
rect 12799 15788 12871 15829
rect 12799 15754 12818 15788
rect 12852 15754 12871 15788
rect 13689 15769 13761 15829
rect 12799 15698 12871 15754
rect 12799 15664 12818 15698
rect 12852 15664 12871 15698
rect 12799 15608 12871 15664
rect 12799 15574 12818 15608
rect 12852 15574 12871 15608
rect 12799 15518 12871 15574
rect 12799 15484 12818 15518
rect 12852 15484 12871 15518
rect 12799 15428 12871 15484
rect 12799 15394 12818 15428
rect 12852 15394 12871 15428
rect 12799 15338 12871 15394
rect 12799 15304 12818 15338
rect 12852 15304 12871 15338
rect 12799 15248 12871 15304
rect 12799 15214 12818 15248
rect 12852 15214 12871 15248
rect 12799 15158 12871 15214
rect 12799 15124 12818 15158
rect 12852 15124 12871 15158
rect 12799 15068 12871 15124
rect 13689 15735 13708 15769
rect 13742 15735 13761 15769
rect 13689 15679 13761 15735
rect 13689 15645 13708 15679
rect 13742 15645 13761 15679
rect 13689 15589 13761 15645
rect 13689 15555 13708 15589
rect 13742 15555 13761 15589
rect 13689 15499 13761 15555
rect 13689 15465 13708 15499
rect 13742 15465 13761 15499
rect 13689 15409 13761 15465
rect 13689 15375 13708 15409
rect 13742 15375 13761 15409
rect 13689 15319 13761 15375
rect 13689 15285 13708 15319
rect 13742 15285 13761 15319
rect 13689 15229 13761 15285
rect 13689 15195 13708 15229
rect 13742 15195 13761 15229
rect 13689 15139 13761 15195
rect 13689 15105 13708 15139
rect 13742 15105 13761 15139
rect 12799 15034 12818 15068
rect 12852 15034 12871 15068
rect 12799 15011 12871 15034
rect 13689 15049 13761 15105
rect 13689 15015 13708 15049
rect 13742 15015 13761 15049
rect 13689 15011 13761 15015
rect 12799 14992 13761 15011
rect 12799 14958 12876 14992
rect 12910 14958 12966 14992
rect 13000 14958 13056 14992
rect 13090 14958 13146 14992
rect 13180 14958 13236 14992
rect 13270 14958 13326 14992
rect 13360 14958 13416 14992
rect 13450 14958 13506 14992
rect 13540 14958 13596 14992
rect 13630 14958 13761 14992
rect 12799 14939 13761 14958
rect 14159 15882 15121 15901
rect 14159 15848 14270 15882
rect 14304 15848 14360 15882
rect 14394 15848 14450 15882
rect 14484 15848 14540 15882
rect 14574 15848 14630 15882
rect 14664 15848 14720 15882
rect 14754 15848 14810 15882
rect 14844 15848 14900 15882
rect 14934 15848 14990 15882
rect 15024 15848 15121 15882
rect 14159 15829 15121 15848
rect 14159 15788 14231 15829
rect 14159 15754 14178 15788
rect 14212 15754 14231 15788
rect 15049 15769 15121 15829
rect 14159 15698 14231 15754
rect 14159 15664 14178 15698
rect 14212 15664 14231 15698
rect 14159 15608 14231 15664
rect 14159 15574 14178 15608
rect 14212 15574 14231 15608
rect 14159 15518 14231 15574
rect 14159 15484 14178 15518
rect 14212 15484 14231 15518
rect 14159 15428 14231 15484
rect 14159 15394 14178 15428
rect 14212 15394 14231 15428
rect 14159 15338 14231 15394
rect 14159 15304 14178 15338
rect 14212 15304 14231 15338
rect 14159 15248 14231 15304
rect 14159 15214 14178 15248
rect 14212 15214 14231 15248
rect 14159 15158 14231 15214
rect 14159 15124 14178 15158
rect 14212 15124 14231 15158
rect 14159 15068 14231 15124
rect 15049 15735 15068 15769
rect 15102 15735 15121 15769
rect 15049 15679 15121 15735
rect 15049 15645 15068 15679
rect 15102 15645 15121 15679
rect 15049 15589 15121 15645
rect 15049 15555 15068 15589
rect 15102 15555 15121 15589
rect 15049 15499 15121 15555
rect 15049 15465 15068 15499
rect 15102 15465 15121 15499
rect 15049 15409 15121 15465
rect 15049 15375 15068 15409
rect 15102 15375 15121 15409
rect 15049 15319 15121 15375
rect 15049 15285 15068 15319
rect 15102 15285 15121 15319
rect 15049 15229 15121 15285
rect 15049 15195 15068 15229
rect 15102 15195 15121 15229
rect 15049 15139 15121 15195
rect 15049 15105 15068 15139
rect 15102 15105 15121 15139
rect 14159 15034 14178 15068
rect 14212 15034 14231 15068
rect 14159 15011 14231 15034
rect 15049 15049 15121 15105
rect 15049 15015 15068 15049
rect 15102 15015 15121 15049
rect 15049 15011 15121 15015
rect 14159 14992 15121 15011
rect 14159 14958 14236 14992
rect 14270 14958 14326 14992
rect 14360 14958 14416 14992
rect 14450 14958 14506 14992
rect 14540 14958 14596 14992
rect 14630 14958 14686 14992
rect 14720 14958 14776 14992
rect 14810 14958 14866 14992
rect 14900 14958 14956 14992
rect 14990 14958 15121 14992
rect 14159 14939 15121 14958
rect 17011 18499 17045 18561
rect 16593 15847 16627 15909
rect 17383 18555 17479 18589
rect 17739 18555 17835 18589
rect 17383 18493 17417 18555
rect 17801 18493 17835 18555
rect 17383 16527 17417 16589
rect 17801 16527 17835 16589
rect 17383 16493 17479 16527
rect 17739 16493 17835 16527
rect 17011 15847 17045 15909
rect 16593 15813 16689 15847
rect 16949 15813 17045 15847
rect 11403 14571 11499 14605
rect 15057 14571 15153 14605
rect 11403 14509 11437 14571
rect 15119 14509 15153 14571
rect 11403 14187 11437 14249
rect 15119 14187 15153 14249
rect 11403 14153 11499 14187
rect 15057 14153 15153 14187
rect 10440 11390 10520 11420
rect 10440 11350 10460 11390
rect 10500 11350 10520 11390
rect 10440 11290 10520 11350
rect 10440 11250 10460 11290
rect 10500 11250 10520 11290
rect 10440 11220 10520 11250
rect 13000 11390 13080 11420
rect 13000 11350 13020 11390
rect 13060 11350 13080 11390
rect 13000 11290 13080 11350
rect 13000 11250 13020 11290
rect 13060 11250 13080 11290
rect 13000 11220 13080 11250
rect 13480 11390 13560 11420
rect 13480 11350 13500 11390
rect 13540 11350 13560 11390
rect 13480 11290 13560 11350
rect 13480 11250 13500 11290
rect 13540 11250 13560 11290
rect 13480 11220 13560 11250
rect 16040 11390 16120 11420
rect 16040 11350 16060 11390
rect 16100 11350 16120 11390
rect 16040 11290 16120 11350
rect 16040 11250 16060 11290
rect 16100 11250 16120 11290
rect 16040 11220 16120 11250
rect 11540 10230 11620 10260
rect 11540 10190 11560 10230
rect 11600 10190 11620 10230
rect 11540 10130 11620 10190
rect 11540 10090 11560 10130
rect 11600 10090 11620 10130
rect 11540 10030 11620 10090
rect 11540 9990 11560 10030
rect 11600 9990 11620 10030
rect 11540 9930 11620 9990
rect 11540 9890 11560 9930
rect 11600 9890 11620 9930
rect 11540 9830 11620 9890
rect 11540 9790 11560 9830
rect 11600 9790 11620 9830
rect 11540 9730 11620 9790
rect 11540 9690 11560 9730
rect 11600 9690 11620 9730
rect 11540 9660 11620 9690
rect 14940 10230 15020 10260
rect 14940 10190 14960 10230
rect 15000 10190 15020 10230
rect 14940 10130 15020 10190
rect 14940 10090 14960 10130
rect 15000 10090 15020 10130
rect 14940 10030 15020 10090
rect 14940 9990 14960 10030
rect 15000 9990 15020 10030
rect 14940 9930 15020 9990
rect 14940 9890 14960 9930
rect 15000 9890 15020 9930
rect 14940 9830 15020 9890
rect 15400 10030 15480 10060
rect 15400 9990 15420 10030
rect 15460 9990 15480 10030
rect 15400 9930 15480 9990
rect 15400 9890 15420 9930
rect 15460 9890 15480 9930
rect 15400 9860 15480 9890
rect 16010 10030 16090 10060
rect 16010 9990 16030 10030
rect 16070 9990 16090 10030
rect 16010 9930 16090 9990
rect 16010 9890 16030 9930
rect 16070 9890 16090 9930
rect 16010 9860 16090 9890
rect 14940 9790 14960 9830
rect 15000 9790 15020 9830
rect 14940 9730 15020 9790
rect 14940 9690 14960 9730
rect 15000 9690 15020 9730
rect 14940 9660 15020 9690
rect 11550 9230 11630 9260
rect 11550 9190 11570 9230
rect 11610 9190 11630 9230
rect 11550 9130 11630 9190
rect 11550 9090 11570 9130
rect 11610 9090 11630 9130
rect 11550 9060 11630 9090
rect 13030 9230 13110 9260
rect 13030 9190 13050 9230
rect 13090 9190 13110 9230
rect 13030 9130 13110 9190
rect 13030 9090 13050 9130
rect 13090 9090 13110 9130
rect 13030 9060 13110 9090
rect 13450 9230 13530 9260
rect 13450 9190 13470 9230
rect 13510 9190 13530 9230
rect 13450 9130 13530 9190
rect 13450 9090 13470 9130
rect 13510 9090 13530 9130
rect 13450 9060 13530 9090
rect 14930 9230 15010 9260
rect 14930 9190 14950 9230
rect 14990 9190 15010 9230
rect 14930 9130 15010 9190
rect 14930 9090 14950 9130
rect 14990 9090 15010 9130
rect 14930 9060 15010 9090
<< psubdiffcont >>
rect 13260 19030 13300 19070
rect 13260 18950 13300 18990
rect 13260 18870 13300 18910
rect 11410 18718 11444 18752
rect 11500 18718 11534 18752
rect 11590 18718 11624 18752
rect 11680 18718 11714 18752
rect 11770 18718 11804 18752
rect 11860 18718 11894 18752
rect 11950 18718 11984 18752
rect 12040 18718 12074 18752
rect 12130 18718 12164 18752
rect 12220 18718 12254 18752
rect 12310 18718 12344 18752
rect 12400 18718 12434 18752
rect 11309 18634 11343 18668
rect 12496 18634 12530 18668
rect 11309 18544 11343 18578
rect 11309 18454 11343 18488
rect 11309 18364 11343 18398
rect 11309 18274 11343 18308
rect 11309 18184 11343 18218
rect 11309 18094 11343 18128
rect 11309 18004 11343 18038
rect 11309 17914 11343 17948
rect 11309 17824 11343 17858
rect 11309 17734 11343 17768
rect 11309 17644 11343 17678
rect 12496 18544 12530 18578
rect 12496 18454 12530 18488
rect 12496 18364 12530 18398
rect 12496 18274 12530 18308
rect 12496 18184 12530 18218
rect 12496 18094 12530 18128
rect 12496 18004 12530 18038
rect 12496 17914 12530 17948
rect 12496 17824 12530 17858
rect 12496 17734 12530 17768
rect 12496 17644 12530 17678
rect 11309 17554 11343 17588
rect 11410 17531 11444 17565
rect 11500 17531 11534 17565
rect 11590 17531 11624 17565
rect 11680 17531 11714 17565
rect 11770 17531 11804 17565
rect 11860 17531 11894 17565
rect 11950 17531 11984 17565
rect 12040 17531 12074 17565
rect 12130 17531 12164 17565
rect 12220 17531 12254 17565
rect 12310 17531 12344 17565
rect 12400 17531 12434 17565
rect 12496 17554 12530 17588
rect 12770 18718 12804 18752
rect 12860 18718 12894 18752
rect 12950 18718 12984 18752
rect 13040 18718 13074 18752
rect 13130 18718 13164 18752
rect 13220 18718 13254 18752
rect 13310 18718 13344 18752
rect 13400 18718 13434 18752
rect 13490 18718 13524 18752
rect 13580 18718 13614 18752
rect 13670 18718 13704 18752
rect 13760 18718 13794 18752
rect 12669 18634 12703 18668
rect 13856 18634 13890 18668
rect 12669 18544 12703 18578
rect 12669 18454 12703 18488
rect 12669 18364 12703 18398
rect 12669 18274 12703 18308
rect 12669 18184 12703 18218
rect 12669 18094 12703 18128
rect 12669 18004 12703 18038
rect 12669 17914 12703 17948
rect 12669 17824 12703 17858
rect 12669 17734 12703 17768
rect 12669 17644 12703 17678
rect 13856 18544 13890 18578
rect 13856 18454 13890 18488
rect 13856 18364 13890 18398
rect 13856 18274 13890 18308
rect 13856 18184 13890 18218
rect 13856 18094 13890 18128
rect 13856 18004 13890 18038
rect 13856 17914 13890 17948
rect 13856 17824 13890 17858
rect 13856 17734 13890 17768
rect 13856 17644 13890 17678
rect 12669 17554 12703 17588
rect 12770 17531 12804 17565
rect 12860 17531 12894 17565
rect 12950 17531 12984 17565
rect 13040 17531 13074 17565
rect 13130 17531 13164 17565
rect 13220 17531 13254 17565
rect 13310 17531 13344 17565
rect 13400 17531 13434 17565
rect 13490 17531 13524 17565
rect 13580 17531 13614 17565
rect 13670 17531 13704 17565
rect 13760 17531 13794 17565
rect 13856 17554 13890 17588
rect 14130 18718 14164 18752
rect 14220 18718 14254 18752
rect 14310 18718 14344 18752
rect 14400 18718 14434 18752
rect 14490 18718 14524 18752
rect 14580 18718 14614 18752
rect 14670 18718 14704 18752
rect 14760 18718 14794 18752
rect 14850 18718 14884 18752
rect 14940 18718 14974 18752
rect 15030 18718 15064 18752
rect 15120 18718 15154 18752
rect 14029 18634 14063 18668
rect 15216 18634 15250 18668
rect 14029 18544 14063 18578
rect 14029 18454 14063 18488
rect 14029 18364 14063 18398
rect 14029 18274 14063 18308
rect 14029 18184 14063 18218
rect 14029 18094 14063 18128
rect 14029 18004 14063 18038
rect 14029 17914 14063 17948
rect 14029 17824 14063 17858
rect 14029 17734 14063 17768
rect 14029 17644 14063 17678
rect 15216 18544 15250 18578
rect 15216 18454 15250 18488
rect 15216 18364 15250 18398
rect 15216 18274 15250 18308
rect 15216 18184 15250 18218
rect 15216 18094 15250 18128
rect 15216 18004 15250 18038
rect 15216 17914 15250 17948
rect 15216 17824 15250 17858
rect 15216 17734 15250 17768
rect 15216 17644 15250 17678
rect 14029 17554 14063 17588
rect 14130 17531 14164 17565
rect 14220 17531 14254 17565
rect 14310 17531 14344 17565
rect 14400 17531 14434 17565
rect 14490 17531 14524 17565
rect 14580 17531 14614 17565
rect 14670 17531 14704 17565
rect 14760 17531 14794 17565
rect 14850 17531 14884 17565
rect 14940 17531 14974 17565
rect 15030 17531 15064 17565
rect 15120 17531 15154 17565
rect 15216 17554 15250 17588
rect 11410 17358 11444 17392
rect 11500 17358 11534 17392
rect 11590 17358 11624 17392
rect 11680 17358 11714 17392
rect 11770 17358 11804 17392
rect 11860 17358 11894 17392
rect 11950 17358 11984 17392
rect 12040 17358 12074 17392
rect 12130 17358 12164 17392
rect 12220 17358 12254 17392
rect 12310 17358 12344 17392
rect 12400 17358 12434 17392
rect 11309 17274 11343 17308
rect 12496 17274 12530 17308
rect 11309 17184 11343 17218
rect 11309 17094 11343 17128
rect 11309 17004 11343 17038
rect 11309 16914 11343 16948
rect 11309 16824 11343 16858
rect 11309 16734 11343 16768
rect 11309 16644 11343 16678
rect 11309 16554 11343 16588
rect 11309 16464 11343 16498
rect 11309 16374 11343 16408
rect 11309 16284 11343 16318
rect 12496 17184 12530 17218
rect 12496 17094 12530 17128
rect 12496 17004 12530 17038
rect 12496 16914 12530 16948
rect 12496 16824 12530 16858
rect 12496 16734 12530 16768
rect 12496 16644 12530 16678
rect 12496 16554 12530 16588
rect 12496 16464 12530 16498
rect 12496 16374 12530 16408
rect 12496 16284 12530 16318
rect 11309 16194 11343 16228
rect 11410 16171 11444 16205
rect 11500 16171 11534 16205
rect 11590 16171 11624 16205
rect 11680 16171 11714 16205
rect 11770 16171 11804 16205
rect 11860 16171 11894 16205
rect 11950 16171 11984 16205
rect 12040 16171 12074 16205
rect 12130 16171 12164 16205
rect 12220 16171 12254 16205
rect 12310 16171 12344 16205
rect 12400 16171 12434 16205
rect 12496 16194 12530 16228
rect 12770 17358 12804 17392
rect 12860 17358 12894 17392
rect 12950 17358 12984 17392
rect 13040 17358 13074 17392
rect 13130 17358 13164 17392
rect 13220 17358 13254 17392
rect 13310 17358 13344 17392
rect 13400 17358 13434 17392
rect 13490 17358 13524 17392
rect 13580 17358 13614 17392
rect 13670 17358 13704 17392
rect 13760 17358 13794 17392
rect 12669 17274 12703 17308
rect 13856 17274 13890 17308
rect 12669 17184 12703 17218
rect 12669 17094 12703 17128
rect 12669 17004 12703 17038
rect 12669 16914 12703 16948
rect 12669 16824 12703 16858
rect 12669 16734 12703 16768
rect 12669 16644 12703 16678
rect 12669 16554 12703 16588
rect 12669 16464 12703 16498
rect 12669 16374 12703 16408
rect 12669 16284 12703 16318
rect 13856 17184 13890 17218
rect 13856 17094 13890 17128
rect 13856 17004 13890 17038
rect 13856 16914 13890 16948
rect 13856 16824 13890 16858
rect 13856 16734 13890 16768
rect 13856 16644 13890 16678
rect 13856 16554 13890 16588
rect 13856 16464 13890 16498
rect 13856 16374 13890 16408
rect 13856 16284 13890 16318
rect 12669 16194 12703 16228
rect 12770 16171 12804 16205
rect 12860 16171 12894 16205
rect 12950 16171 12984 16205
rect 13040 16171 13074 16205
rect 13130 16171 13164 16205
rect 13220 16171 13254 16205
rect 13310 16171 13344 16205
rect 13400 16171 13434 16205
rect 13490 16171 13524 16205
rect 13580 16171 13614 16205
rect 13670 16171 13704 16205
rect 13760 16171 13794 16205
rect 13856 16194 13890 16228
rect 14130 17358 14164 17392
rect 14220 17358 14254 17392
rect 14310 17358 14344 17392
rect 14400 17358 14434 17392
rect 14490 17358 14524 17392
rect 14580 17358 14614 17392
rect 14670 17358 14704 17392
rect 14760 17358 14794 17392
rect 14850 17358 14884 17392
rect 14940 17358 14974 17392
rect 15030 17358 15064 17392
rect 15120 17358 15154 17392
rect 14029 17274 14063 17308
rect 15216 17274 15250 17308
rect 14029 17184 14063 17218
rect 14029 17094 14063 17128
rect 14029 17004 14063 17038
rect 14029 16914 14063 16948
rect 14029 16824 14063 16858
rect 14029 16734 14063 16768
rect 14029 16644 14063 16678
rect 14029 16554 14063 16588
rect 14029 16464 14063 16498
rect 14029 16374 14063 16408
rect 14029 16284 14063 16318
rect 15216 17184 15250 17218
rect 15216 17094 15250 17128
rect 15216 17004 15250 17038
rect 15216 16914 15250 16948
rect 15216 16824 15250 16858
rect 15216 16734 15250 16768
rect 15216 16644 15250 16678
rect 15216 16554 15250 16588
rect 15216 16464 15250 16498
rect 15216 16374 15250 16408
rect 15216 16284 15250 16318
rect 14029 16194 14063 16228
rect 14130 16171 14164 16205
rect 14220 16171 14254 16205
rect 14310 16171 14344 16205
rect 14400 16171 14434 16205
rect 14490 16171 14524 16205
rect 14580 16171 14614 16205
rect 14670 16171 14704 16205
rect 14760 16171 14794 16205
rect 14850 16171 14884 16205
rect 14940 16171 14974 16205
rect 15030 16171 15064 16205
rect 15120 16171 15154 16205
rect 15216 16194 15250 16228
rect 11410 15998 11444 16032
rect 11500 15998 11534 16032
rect 11590 15998 11624 16032
rect 11680 15998 11714 16032
rect 11770 15998 11804 16032
rect 11860 15998 11894 16032
rect 11950 15998 11984 16032
rect 12040 15998 12074 16032
rect 12130 15998 12164 16032
rect 12220 15998 12254 16032
rect 12310 15998 12344 16032
rect 12400 15998 12434 16032
rect 11309 15914 11343 15948
rect 12496 15914 12530 15948
rect 11309 15824 11343 15858
rect 11309 15734 11343 15768
rect 11309 15644 11343 15678
rect 11309 15554 11343 15588
rect 11309 15464 11343 15498
rect 11309 15374 11343 15408
rect 11309 15284 11343 15318
rect 11309 15194 11343 15228
rect 11309 15104 11343 15138
rect 11309 15014 11343 15048
rect 11309 14924 11343 14958
rect 12496 15824 12530 15858
rect 12496 15734 12530 15768
rect 12496 15644 12530 15678
rect 12496 15554 12530 15588
rect 12496 15464 12530 15498
rect 12496 15374 12530 15408
rect 12496 15284 12530 15318
rect 12496 15194 12530 15228
rect 12496 15104 12530 15138
rect 12496 15014 12530 15048
rect 12496 14924 12530 14958
rect 11309 14834 11343 14868
rect 11410 14811 11444 14845
rect 11500 14811 11534 14845
rect 11590 14811 11624 14845
rect 11680 14811 11714 14845
rect 11770 14811 11804 14845
rect 11860 14811 11894 14845
rect 11950 14811 11984 14845
rect 12040 14811 12074 14845
rect 12130 14811 12164 14845
rect 12220 14811 12254 14845
rect 12310 14811 12344 14845
rect 12400 14811 12434 14845
rect 12496 14834 12530 14868
rect 12770 15998 12804 16032
rect 12860 15998 12894 16032
rect 12950 15998 12984 16032
rect 13040 15998 13074 16032
rect 13130 15998 13164 16032
rect 13220 15998 13254 16032
rect 13310 15998 13344 16032
rect 13400 15998 13434 16032
rect 13490 15998 13524 16032
rect 13580 15998 13614 16032
rect 13670 15998 13704 16032
rect 13760 15998 13794 16032
rect 12669 15914 12703 15948
rect 13856 15914 13890 15948
rect 12669 15824 12703 15858
rect 12669 15734 12703 15768
rect 12669 15644 12703 15678
rect 12669 15554 12703 15588
rect 12669 15464 12703 15498
rect 12669 15374 12703 15408
rect 12669 15284 12703 15318
rect 12669 15194 12703 15228
rect 12669 15104 12703 15138
rect 12669 15014 12703 15048
rect 12669 14924 12703 14958
rect 13856 15824 13890 15858
rect 13856 15734 13890 15768
rect 13856 15644 13890 15678
rect 13856 15554 13890 15588
rect 13856 15464 13890 15498
rect 13856 15374 13890 15408
rect 13856 15284 13890 15318
rect 13856 15194 13890 15228
rect 13856 15104 13890 15138
rect 13856 15014 13890 15048
rect 13856 14924 13890 14958
rect 12669 14834 12703 14868
rect 12770 14811 12804 14845
rect 12860 14811 12894 14845
rect 12950 14811 12984 14845
rect 13040 14811 13074 14845
rect 13130 14811 13164 14845
rect 13220 14811 13254 14845
rect 13310 14811 13344 14845
rect 13400 14811 13434 14845
rect 13490 14811 13524 14845
rect 13580 14811 13614 14845
rect 13670 14811 13704 14845
rect 13760 14811 13794 14845
rect 13856 14834 13890 14868
rect 14130 15998 14164 16032
rect 14220 15998 14254 16032
rect 14310 15998 14344 16032
rect 14400 15998 14434 16032
rect 14490 15998 14524 16032
rect 14580 15998 14614 16032
rect 14670 15998 14704 16032
rect 14760 15998 14794 16032
rect 14850 15998 14884 16032
rect 14940 15998 14974 16032
rect 15030 15998 15064 16032
rect 15120 15998 15154 16032
rect 14029 15914 14063 15948
rect 15216 15914 15250 15948
rect 14029 15824 14063 15858
rect 14029 15734 14063 15768
rect 14029 15644 14063 15678
rect 14029 15554 14063 15588
rect 14029 15464 14063 15498
rect 14029 15374 14063 15408
rect 14029 15284 14063 15318
rect 14029 15194 14063 15228
rect 14029 15104 14063 15138
rect 14029 15014 14063 15048
rect 14029 14924 14063 14958
rect 15216 15824 15250 15858
rect 15216 15734 15250 15768
rect 15216 15644 15250 15678
rect 15216 15554 15250 15588
rect 15216 15464 15250 15498
rect 15216 15374 15250 15408
rect 15216 15284 15250 15318
rect 15216 15194 15250 15228
rect 15216 15104 15250 15138
rect 15216 15014 15250 15048
rect 15216 14924 15250 14958
rect 14029 14834 14063 14868
rect 14130 14811 14164 14845
rect 14220 14811 14254 14845
rect 14310 14811 14344 14845
rect 14400 14811 14434 14845
rect 14490 14811 14524 14845
rect 14580 14811 14614 14845
rect 14670 14811 14704 14845
rect 14760 14811 14794 14845
rect 14850 14811 14884 14845
rect 14940 14811 14974 14845
rect 15030 14811 15064 14845
rect 15120 14811 15154 14845
rect 15216 14834 15250 14868
rect 15420 13810 15460 13850
rect 15420 13710 15460 13750
rect 11920 13200 11960 13240
rect 11920 13100 11960 13140
rect 11920 13000 11960 13040
rect 11920 12900 11960 12940
rect 11920 12800 11960 12840
rect 14600 13200 14640 13240
rect 14600 13100 14640 13140
rect 14600 13000 14640 13040
rect 14600 12900 14640 12940
rect 14600 12800 14640 12840
rect 12820 12280 12860 12320
rect 12820 12200 12860 12240
rect 12820 12120 12860 12160
rect 13700 12280 13740 12320
rect 13700 12200 13740 12240
rect 13700 12120 13740 12160
<< nsubdiffcont >>
rect 8699 18555 8959 18589
rect 8603 16589 8637 18493
rect 9021 16589 9055 18493
rect 8699 16493 8959 16527
rect 9479 18561 9739 18595
rect 9383 15019 9417 18499
rect 9801 15019 9835 18499
rect 10259 18563 10851 18597
rect 10163 16243 10197 18501
rect 10913 16243 10947 18501
rect 11550 18568 11584 18602
rect 11640 18568 11674 18602
rect 11730 18568 11764 18602
rect 11820 18568 11854 18602
rect 11910 18568 11944 18602
rect 12000 18568 12034 18602
rect 12090 18568 12124 18602
rect 12180 18568 12214 18602
rect 12270 18568 12304 18602
rect 11458 18474 11492 18508
rect 11458 18384 11492 18418
rect 11458 18294 11492 18328
rect 11458 18204 11492 18238
rect 11458 18114 11492 18148
rect 11458 18024 11492 18058
rect 11458 17934 11492 17968
rect 11458 17844 11492 17878
rect 12348 18455 12382 18489
rect 12348 18365 12382 18399
rect 12348 18275 12382 18309
rect 12348 18185 12382 18219
rect 12348 18095 12382 18129
rect 12348 18005 12382 18039
rect 12348 17915 12382 17949
rect 12348 17825 12382 17859
rect 11458 17754 11492 17788
rect 12348 17735 12382 17769
rect 11516 17678 11550 17712
rect 11606 17678 11640 17712
rect 11696 17678 11730 17712
rect 11786 17678 11820 17712
rect 11876 17678 11910 17712
rect 11966 17678 12000 17712
rect 12056 17678 12090 17712
rect 12146 17678 12180 17712
rect 12236 17678 12270 17712
rect 12910 18568 12944 18602
rect 13000 18568 13034 18602
rect 13090 18568 13124 18602
rect 13180 18568 13214 18602
rect 13270 18568 13304 18602
rect 13360 18568 13394 18602
rect 13450 18568 13484 18602
rect 13540 18568 13574 18602
rect 13630 18568 13664 18602
rect 12818 18474 12852 18508
rect 12818 18384 12852 18418
rect 12818 18294 12852 18328
rect 12818 18204 12852 18238
rect 12818 18114 12852 18148
rect 12818 18024 12852 18058
rect 12818 17934 12852 17968
rect 12818 17844 12852 17878
rect 13708 18455 13742 18489
rect 13708 18365 13742 18399
rect 13708 18275 13742 18309
rect 13708 18185 13742 18219
rect 13708 18095 13742 18129
rect 13708 18005 13742 18039
rect 13708 17915 13742 17949
rect 13708 17825 13742 17859
rect 12818 17754 12852 17788
rect 13708 17735 13742 17769
rect 12876 17678 12910 17712
rect 12966 17678 13000 17712
rect 13056 17678 13090 17712
rect 13146 17678 13180 17712
rect 13236 17678 13270 17712
rect 13326 17678 13360 17712
rect 13416 17678 13450 17712
rect 13506 17678 13540 17712
rect 13596 17678 13630 17712
rect 14270 18568 14304 18602
rect 14360 18568 14394 18602
rect 14450 18568 14484 18602
rect 14540 18568 14574 18602
rect 14630 18568 14664 18602
rect 14720 18568 14754 18602
rect 14810 18568 14844 18602
rect 14900 18568 14934 18602
rect 14990 18568 15024 18602
rect 14178 18474 14212 18508
rect 14178 18384 14212 18418
rect 14178 18294 14212 18328
rect 14178 18204 14212 18238
rect 14178 18114 14212 18148
rect 14178 18024 14212 18058
rect 14178 17934 14212 17968
rect 14178 17844 14212 17878
rect 15068 18455 15102 18489
rect 15068 18365 15102 18399
rect 15068 18275 15102 18309
rect 15068 18185 15102 18219
rect 15068 18095 15102 18129
rect 15068 18005 15102 18039
rect 15068 17915 15102 17949
rect 15068 17825 15102 17859
rect 14178 17754 14212 17788
rect 15068 17735 15102 17769
rect 14236 17678 14270 17712
rect 14326 17678 14360 17712
rect 14416 17678 14450 17712
rect 14506 17678 14540 17712
rect 14596 17678 14630 17712
rect 14686 17678 14720 17712
rect 14776 17678 14810 17712
rect 14866 17678 14900 17712
rect 14956 17678 14990 17712
rect 15579 18563 16171 18597
rect 10259 16147 10851 16181
rect 11550 17208 11584 17242
rect 11640 17208 11674 17242
rect 11730 17208 11764 17242
rect 11820 17208 11854 17242
rect 11910 17208 11944 17242
rect 12000 17208 12034 17242
rect 12090 17208 12124 17242
rect 12180 17208 12214 17242
rect 12270 17208 12304 17242
rect 11458 17114 11492 17148
rect 11458 17024 11492 17058
rect 11458 16934 11492 16968
rect 11458 16844 11492 16878
rect 11458 16754 11492 16788
rect 11458 16664 11492 16698
rect 11458 16574 11492 16608
rect 11458 16484 11492 16518
rect 12348 17095 12382 17129
rect 12348 17005 12382 17039
rect 12348 16915 12382 16949
rect 12348 16825 12382 16859
rect 12348 16735 12382 16769
rect 12348 16645 12382 16679
rect 12348 16555 12382 16589
rect 12348 16465 12382 16499
rect 11458 16394 11492 16428
rect 12348 16375 12382 16409
rect 11516 16318 11550 16352
rect 11606 16318 11640 16352
rect 11696 16318 11730 16352
rect 11786 16318 11820 16352
rect 11876 16318 11910 16352
rect 11966 16318 12000 16352
rect 12056 16318 12090 16352
rect 12146 16318 12180 16352
rect 12236 16318 12270 16352
rect 12910 17208 12944 17242
rect 13000 17208 13034 17242
rect 13090 17208 13124 17242
rect 13180 17208 13214 17242
rect 13270 17208 13304 17242
rect 13360 17208 13394 17242
rect 13450 17208 13484 17242
rect 13540 17208 13574 17242
rect 13630 17208 13664 17242
rect 12818 17114 12852 17148
rect 12818 17024 12852 17058
rect 12818 16934 12852 16968
rect 12818 16844 12852 16878
rect 12818 16754 12852 16788
rect 12818 16664 12852 16698
rect 12818 16574 12852 16608
rect 12818 16484 12852 16518
rect 13708 17095 13742 17129
rect 13708 17005 13742 17039
rect 13708 16915 13742 16949
rect 13708 16825 13742 16859
rect 13708 16735 13742 16769
rect 13708 16645 13742 16679
rect 13708 16555 13742 16589
rect 13708 16465 13742 16499
rect 12818 16394 12852 16428
rect 13708 16375 13742 16409
rect 12876 16318 12910 16352
rect 12966 16318 13000 16352
rect 13056 16318 13090 16352
rect 13146 16318 13180 16352
rect 13236 16318 13270 16352
rect 13326 16318 13360 16352
rect 13416 16318 13450 16352
rect 13506 16318 13540 16352
rect 13596 16318 13630 16352
rect 14270 17208 14304 17242
rect 14360 17208 14394 17242
rect 14450 17208 14484 17242
rect 14540 17208 14574 17242
rect 14630 17208 14664 17242
rect 14720 17208 14754 17242
rect 14810 17208 14844 17242
rect 14900 17208 14934 17242
rect 14990 17208 15024 17242
rect 14178 17114 14212 17148
rect 14178 17024 14212 17058
rect 14178 16934 14212 16968
rect 14178 16844 14212 16878
rect 14178 16754 14212 16788
rect 14178 16664 14212 16698
rect 14178 16574 14212 16608
rect 14178 16484 14212 16518
rect 15068 17095 15102 17129
rect 15068 17005 15102 17039
rect 15068 16915 15102 16949
rect 15068 16825 15102 16859
rect 15068 16735 15102 16769
rect 15068 16645 15102 16679
rect 15068 16555 15102 16589
rect 15068 16465 15102 16499
rect 14178 16394 14212 16428
rect 15068 16375 15102 16409
rect 14236 16318 14270 16352
rect 14326 16318 14360 16352
rect 14416 16318 14450 16352
rect 14506 16318 14540 16352
rect 14596 16318 14630 16352
rect 14686 16318 14720 16352
rect 14776 16318 14810 16352
rect 14866 16318 14900 16352
rect 14956 16318 14990 16352
rect 15483 16243 15517 18501
rect 16233 16243 16267 18501
rect 15579 16147 16171 16181
rect 16689 18561 16949 18595
rect 9479 14923 9739 14957
rect 11550 15848 11584 15882
rect 11640 15848 11674 15882
rect 11730 15848 11764 15882
rect 11820 15848 11854 15882
rect 11910 15848 11944 15882
rect 12000 15848 12034 15882
rect 12090 15848 12124 15882
rect 12180 15848 12214 15882
rect 12270 15848 12304 15882
rect 11458 15754 11492 15788
rect 11458 15664 11492 15698
rect 11458 15574 11492 15608
rect 11458 15484 11492 15518
rect 11458 15394 11492 15428
rect 11458 15304 11492 15338
rect 11458 15214 11492 15248
rect 11458 15124 11492 15158
rect 12348 15735 12382 15769
rect 12348 15645 12382 15679
rect 12348 15555 12382 15589
rect 12348 15465 12382 15499
rect 12348 15375 12382 15409
rect 12348 15285 12382 15319
rect 12348 15195 12382 15229
rect 12348 15105 12382 15139
rect 11458 15034 11492 15068
rect 12348 15015 12382 15049
rect 11516 14958 11550 14992
rect 11606 14958 11640 14992
rect 11696 14958 11730 14992
rect 11786 14958 11820 14992
rect 11876 14958 11910 14992
rect 11966 14958 12000 14992
rect 12056 14958 12090 14992
rect 12146 14958 12180 14992
rect 12236 14958 12270 14992
rect 12910 15848 12944 15882
rect 13000 15848 13034 15882
rect 13090 15848 13124 15882
rect 13180 15848 13214 15882
rect 13270 15848 13304 15882
rect 13360 15848 13394 15882
rect 13450 15848 13484 15882
rect 13540 15848 13574 15882
rect 13630 15848 13664 15882
rect 12818 15754 12852 15788
rect 12818 15664 12852 15698
rect 12818 15574 12852 15608
rect 12818 15484 12852 15518
rect 12818 15394 12852 15428
rect 12818 15304 12852 15338
rect 12818 15214 12852 15248
rect 12818 15124 12852 15158
rect 13708 15735 13742 15769
rect 13708 15645 13742 15679
rect 13708 15555 13742 15589
rect 13708 15465 13742 15499
rect 13708 15375 13742 15409
rect 13708 15285 13742 15319
rect 13708 15195 13742 15229
rect 13708 15105 13742 15139
rect 12818 15034 12852 15068
rect 13708 15015 13742 15049
rect 12876 14958 12910 14992
rect 12966 14958 13000 14992
rect 13056 14958 13090 14992
rect 13146 14958 13180 14992
rect 13236 14958 13270 14992
rect 13326 14958 13360 14992
rect 13416 14958 13450 14992
rect 13506 14958 13540 14992
rect 13596 14958 13630 14992
rect 14270 15848 14304 15882
rect 14360 15848 14394 15882
rect 14450 15848 14484 15882
rect 14540 15848 14574 15882
rect 14630 15848 14664 15882
rect 14720 15848 14754 15882
rect 14810 15848 14844 15882
rect 14900 15848 14934 15882
rect 14990 15848 15024 15882
rect 14178 15754 14212 15788
rect 14178 15664 14212 15698
rect 14178 15574 14212 15608
rect 14178 15484 14212 15518
rect 14178 15394 14212 15428
rect 14178 15304 14212 15338
rect 14178 15214 14212 15248
rect 14178 15124 14212 15158
rect 15068 15735 15102 15769
rect 15068 15645 15102 15679
rect 15068 15555 15102 15589
rect 15068 15465 15102 15499
rect 15068 15375 15102 15409
rect 15068 15285 15102 15319
rect 15068 15195 15102 15229
rect 15068 15105 15102 15139
rect 14178 15034 14212 15068
rect 15068 15015 15102 15049
rect 14236 14958 14270 14992
rect 14326 14958 14360 14992
rect 14416 14958 14450 14992
rect 14506 14958 14540 14992
rect 14596 14958 14630 14992
rect 14686 14958 14720 14992
rect 14776 14958 14810 14992
rect 14866 14958 14900 14992
rect 14956 14958 14990 14992
rect 16593 15909 16627 18499
rect 17011 15909 17045 18499
rect 17479 18555 17739 18589
rect 17383 16589 17417 18493
rect 17801 16589 17835 18493
rect 17479 16493 17739 16527
rect 16689 15813 16949 15847
rect 11499 14571 15057 14605
rect 11403 14249 11437 14509
rect 15119 14249 15153 14509
rect 11499 14153 15057 14187
rect 10460 11350 10500 11390
rect 10460 11250 10500 11290
rect 13020 11350 13060 11390
rect 13020 11250 13060 11290
rect 13500 11350 13540 11390
rect 13500 11250 13540 11290
rect 16060 11350 16100 11390
rect 16060 11250 16100 11290
rect 11560 10190 11600 10230
rect 11560 10090 11600 10130
rect 11560 9990 11600 10030
rect 11560 9890 11600 9930
rect 11560 9790 11600 9830
rect 11560 9690 11600 9730
rect 14960 10190 15000 10230
rect 14960 10090 15000 10130
rect 14960 9990 15000 10030
rect 14960 9890 15000 9930
rect 15420 9990 15460 10030
rect 15420 9890 15460 9930
rect 16030 9990 16070 10030
rect 16030 9890 16070 9930
rect 14960 9790 15000 9830
rect 14960 9690 15000 9730
rect 11570 9190 11610 9230
rect 11570 9090 11610 9130
rect 13050 9190 13090 9230
rect 13050 9090 13090 9130
rect 13470 9190 13510 9230
rect 13470 9090 13510 9130
rect 14950 9190 14990 9230
rect 14950 9090 14990 9130
<< poly >>
rect 11240 13880 13240 13910
rect 13320 13880 15320 13910
rect 11240 13650 13240 13680
rect 13320 13650 15320 13680
rect 11320 13630 11400 13650
rect 11320 13590 11340 13630
rect 11380 13590 11400 13630
rect 11320 13570 11400 13590
rect 11480 13630 11560 13650
rect 11480 13590 11500 13630
rect 11540 13590 11560 13630
rect 11480 13570 11560 13590
rect 11640 13630 11720 13650
rect 11640 13590 11660 13630
rect 11700 13590 11720 13630
rect 11640 13570 11720 13590
rect 11800 13630 11880 13650
rect 11800 13590 11820 13630
rect 11860 13590 11880 13630
rect 11800 13570 11880 13590
rect 11960 13630 12040 13650
rect 11960 13590 11980 13630
rect 12020 13590 12040 13630
rect 11960 13570 12040 13590
rect 12120 13630 12200 13650
rect 12120 13590 12140 13630
rect 12180 13590 12200 13630
rect 12120 13570 12200 13590
rect 12280 13630 12360 13650
rect 12280 13590 12300 13630
rect 12340 13590 12360 13630
rect 12280 13570 12360 13590
rect 12440 13630 12520 13650
rect 12440 13590 12460 13630
rect 12500 13590 12520 13630
rect 12440 13570 12520 13590
rect 12600 13630 12680 13650
rect 12600 13590 12620 13630
rect 12660 13590 12680 13630
rect 12600 13570 12680 13590
rect 12760 13630 12840 13650
rect 12760 13590 12780 13630
rect 12820 13590 12840 13630
rect 12760 13570 12840 13590
rect 12920 13630 13000 13650
rect 12920 13590 12940 13630
rect 12980 13590 13000 13630
rect 12920 13570 13000 13590
rect 13080 13630 13160 13650
rect 13080 13590 13100 13630
rect 13140 13590 13160 13630
rect 13080 13570 13160 13590
rect 13400 13630 13480 13650
rect 13400 13590 13420 13630
rect 13460 13590 13480 13630
rect 13400 13570 13480 13590
rect 13560 13630 13640 13650
rect 13560 13590 13580 13630
rect 13620 13590 13640 13630
rect 13560 13570 13640 13590
rect 13720 13630 13800 13650
rect 13720 13590 13740 13630
rect 13780 13590 13800 13630
rect 13720 13570 13800 13590
rect 13880 13630 13960 13650
rect 13880 13590 13900 13630
rect 13940 13590 13960 13630
rect 13880 13570 13960 13590
rect 14040 13630 14120 13650
rect 14040 13590 14060 13630
rect 14100 13590 14120 13630
rect 14040 13570 14120 13590
rect 14200 13630 14280 13650
rect 14200 13590 14220 13630
rect 14260 13590 14280 13630
rect 14200 13570 14280 13590
rect 14360 13630 14440 13650
rect 14360 13590 14380 13630
rect 14420 13590 14440 13630
rect 14360 13570 14440 13590
rect 14520 13630 14600 13650
rect 14520 13590 14540 13630
rect 14580 13590 14600 13630
rect 14520 13570 14600 13590
rect 14680 13630 14760 13650
rect 14680 13590 14700 13630
rect 14740 13590 14760 13630
rect 14680 13570 14760 13590
rect 14840 13630 14920 13650
rect 14840 13590 14860 13630
rect 14900 13590 14920 13630
rect 14840 13570 14920 13590
rect 15000 13630 15080 13650
rect 15000 13590 15020 13630
rect 15060 13590 15080 13630
rect 15000 13570 15080 13590
rect 15160 13630 15240 13650
rect 15160 13590 15180 13630
rect 15220 13590 15240 13630
rect 15160 13570 15240 13590
rect 10820 13270 11820 13300
rect 12060 13270 13060 13300
rect 13500 13270 14500 13300
rect 14740 13270 15740 13300
rect 10820 12740 11820 12770
rect 12060 12740 13060 12770
rect 13500 12740 14500 12770
rect 14740 12740 15740 12770
rect 10920 12720 11000 12740
rect 10920 12680 10940 12720
rect 10980 12680 11000 12720
rect 10920 12660 11000 12680
rect 11160 12720 11240 12740
rect 11160 12680 11180 12720
rect 11220 12680 11240 12720
rect 11160 12660 11240 12680
rect 11400 12720 11480 12740
rect 11400 12680 11420 12720
rect 11460 12680 11480 12720
rect 11400 12660 11480 12680
rect 11640 12720 11720 12740
rect 11640 12680 11660 12720
rect 11700 12680 11720 12720
rect 11640 12660 11720 12680
rect 12280 12720 12360 12740
rect 12280 12680 12300 12720
rect 12340 12680 12360 12720
rect 12280 12660 12360 12680
rect 12520 12720 12600 12740
rect 12520 12680 12540 12720
rect 12580 12680 12600 12720
rect 12520 12660 12600 12680
rect 12760 12720 12840 12740
rect 12760 12680 12780 12720
rect 12820 12680 12840 12720
rect 12760 12660 12840 12680
rect 13720 12720 13800 12740
rect 13720 12680 13740 12720
rect 13780 12680 13800 12720
rect 13720 12660 13800 12680
rect 13960 12720 14040 12740
rect 13960 12680 13980 12720
rect 14020 12680 14040 12720
rect 13960 12660 14040 12680
rect 14200 12720 14280 12740
rect 14200 12680 14220 12720
rect 14260 12680 14280 12720
rect 14200 12660 14280 12680
rect 14840 12720 14920 12740
rect 14840 12680 14860 12720
rect 14900 12680 14920 12720
rect 14840 12660 14920 12680
rect 15080 12720 15160 12740
rect 15080 12680 15100 12720
rect 15140 12680 15160 12720
rect 15080 12660 15160 12680
rect 15320 12720 15400 12740
rect 15320 12680 15340 12720
rect 15380 12680 15400 12720
rect 15320 12660 15400 12680
rect 15560 12720 15640 12740
rect 15560 12680 15580 12720
rect 15620 12680 15640 12720
rect 15560 12660 15640 12680
rect 11431 12342 11489 12360
rect 11431 12308 11443 12342
rect 11477 12308 11489 12342
rect 11431 12290 11489 12308
rect 11791 12342 11849 12360
rect 11791 12308 11803 12342
rect 11837 12308 11849 12342
rect 11791 12290 11849 12308
rect 11911 12342 11969 12360
rect 11911 12308 11923 12342
rect 11957 12308 11969 12342
rect 11911 12290 11969 12308
rect 12271 12342 12329 12360
rect 12271 12308 12283 12342
rect 12317 12308 12329 12342
rect 12271 12290 12329 12308
rect 12391 12342 12449 12360
rect 12391 12308 12403 12342
rect 12437 12308 12449 12342
rect 12391 12290 12449 12308
rect 11440 12260 11480 12290
rect 11560 12260 11600 12290
rect 11680 12260 11720 12290
rect 11800 12260 11840 12290
rect 11920 12260 11960 12290
rect 12040 12260 12080 12290
rect 12160 12260 12200 12290
rect 12280 12260 12320 12290
rect 12400 12260 12440 12290
rect 12520 12260 12560 12290
rect 11440 12130 11480 12160
rect 11560 12130 11600 12160
rect 11532 12112 11600 12130
rect 11532 12078 11544 12112
rect 11578 12078 11600 12112
rect 11532 12060 11600 12078
rect 11680 12130 11720 12160
rect 11800 12130 11840 12160
rect 11920 12130 11960 12160
rect 12040 12130 12080 12160
rect 11680 12112 11748 12130
rect 11680 12078 11702 12112
rect 11736 12078 11748 12112
rect 11680 12060 11748 12078
rect 12014 12112 12080 12130
rect 12014 12078 12026 12112
rect 12060 12078 12080 12112
rect 12014 12060 12080 12078
rect 12160 12130 12200 12160
rect 12280 12130 12320 12160
rect 12400 12130 12440 12160
rect 12520 12130 12560 12160
rect 12160 12112 12226 12130
rect 12160 12078 12180 12112
rect 12214 12078 12226 12112
rect 12160 12060 12226 12078
rect 12492 12112 12560 12130
rect 12492 12078 12504 12112
rect 12538 12078 12560 12112
rect 14111 12342 14169 12360
rect 14111 12308 14123 12342
rect 14157 12308 14169 12342
rect 14111 12290 14169 12308
rect 14231 12342 14289 12360
rect 14231 12308 14243 12342
rect 14277 12308 14289 12342
rect 14231 12290 14289 12308
rect 14591 12342 14649 12360
rect 14591 12308 14603 12342
rect 14637 12308 14649 12342
rect 14591 12290 14649 12308
rect 14711 12342 14769 12360
rect 14711 12308 14723 12342
rect 14757 12308 14769 12342
rect 14711 12290 14769 12308
rect 15071 12342 15129 12360
rect 15071 12308 15083 12342
rect 15117 12308 15129 12342
rect 15071 12290 15129 12308
rect 14000 12260 14040 12290
rect 14120 12260 14160 12290
rect 14240 12260 14280 12290
rect 14360 12260 14400 12290
rect 14480 12260 14520 12290
rect 14600 12260 14640 12290
rect 14720 12260 14760 12290
rect 14840 12260 14880 12290
rect 14960 12260 15000 12290
rect 15080 12260 15120 12290
rect 14000 12130 14040 12160
rect 14120 12130 14160 12160
rect 14240 12130 14280 12160
rect 14360 12130 14400 12160
rect 14000 12112 14068 12130
rect 12492 12060 12560 12078
rect 14000 12078 14022 12112
rect 14056 12078 14068 12112
rect 14000 12060 14068 12078
rect 14334 12112 14400 12130
rect 14334 12078 14346 12112
rect 14380 12078 14400 12112
rect 14334 12060 14400 12078
rect 14480 12130 14520 12160
rect 14600 12130 14640 12160
rect 14720 12130 14760 12160
rect 14840 12130 14880 12160
rect 14480 12112 14546 12130
rect 14480 12078 14500 12112
rect 14534 12078 14546 12112
rect 14480 12060 14546 12078
rect 14812 12112 14880 12130
rect 14812 12078 14824 12112
rect 14858 12078 14880 12112
rect 14812 12060 14880 12078
rect 14960 12130 15000 12160
rect 15080 12130 15120 12160
rect 14960 12112 15028 12130
rect 14960 12078 14982 12112
rect 15016 12078 15028 12112
rect 14960 12060 15028 12078
rect 10710 11520 10770 11540
rect 10710 11480 10720 11520
rect 10760 11480 10770 11520
rect 10710 11460 10770 11480
rect 10880 11510 10960 11530
rect 10880 11470 10900 11510
rect 10940 11470 10960 11510
rect 11370 11510 11430 11530
rect 11370 11470 11380 11510
rect 11420 11470 11430 11510
rect 11600 11510 11680 11530
rect 11600 11470 11620 11510
rect 11660 11470 11680 11510
rect 12090 11510 12150 11530
rect 12090 11470 12100 11510
rect 12140 11470 12150 11510
rect 12320 11510 12400 11530
rect 12320 11470 12340 11510
rect 12380 11470 12400 11510
rect 12750 11510 12810 11530
rect 12750 11470 12760 11510
rect 12800 11470 12810 11510
rect 10600 11420 10640 11450
rect 10720 11420 10760 11460
rect 10840 11440 11240 11470
rect 10840 11420 10880 11440
rect 10960 11420 11000 11440
rect 11080 11420 11120 11440
rect 11200 11420 11240 11440
rect 11320 11440 11480 11470
rect 11320 11420 11360 11440
rect 11440 11420 11480 11440
rect 11560 11440 11960 11470
rect 11560 11420 11600 11440
rect 11680 11420 11720 11440
rect 11800 11420 11840 11440
rect 11920 11420 11960 11440
rect 12040 11440 12200 11470
rect 12040 11420 12080 11440
rect 12160 11420 12200 11440
rect 12280 11440 12680 11470
rect 12750 11450 12810 11470
rect 13750 11510 13810 11530
rect 13750 11470 13760 11510
rect 13800 11470 13810 11510
rect 14160 11510 14240 11530
rect 14160 11470 14180 11510
rect 14220 11470 14240 11510
rect 14410 11510 14470 11530
rect 14410 11470 14420 11510
rect 14460 11470 14470 11510
rect 14880 11510 14960 11530
rect 14880 11470 14900 11510
rect 14940 11470 14960 11510
rect 15130 11510 15190 11530
rect 15130 11470 15140 11510
rect 15180 11470 15190 11510
rect 15600 11510 15680 11530
rect 15600 11470 15620 11510
rect 15660 11470 15680 11510
rect 15790 11520 15850 11540
rect 15790 11480 15800 11520
rect 15840 11480 15850 11520
rect 13750 11450 13810 11470
rect 12280 11420 12320 11440
rect 12400 11420 12440 11440
rect 12520 11420 12560 11440
rect 12640 11420 12680 11440
rect 12760 11420 12800 11450
rect 12880 11420 12920 11450
rect 13640 11420 13680 11450
rect 13760 11420 13800 11450
rect 13880 11440 14280 11470
rect 13880 11420 13920 11440
rect 14000 11420 14040 11440
rect 14120 11420 14160 11440
rect 14240 11420 14280 11440
rect 14360 11440 14520 11470
rect 14360 11420 14400 11440
rect 14480 11420 14520 11440
rect 14600 11440 15000 11470
rect 14600 11420 14640 11440
rect 14720 11420 14760 11440
rect 14840 11420 14880 11440
rect 14960 11420 15000 11440
rect 15080 11440 15240 11470
rect 15080 11420 15120 11440
rect 15200 11420 15240 11440
rect 15320 11440 15720 11470
rect 15790 11460 15850 11480
rect 15320 11420 15360 11440
rect 15440 11420 15480 11440
rect 15560 11420 15600 11440
rect 15680 11420 15720 11440
rect 15800 11420 15840 11460
rect 15920 11420 15960 11450
rect 10600 11190 10640 11220
rect 10720 11190 10760 11220
rect 10840 11190 10880 11220
rect 10960 11190 11000 11220
rect 11080 11190 11120 11220
rect 11200 11190 11240 11220
rect 11320 11190 11360 11220
rect 11440 11190 11480 11220
rect 11560 11190 11600 11220
rect 11680 11190 11720 11220
rect 11800 11190 11840 11220
rect 11920 11190 11960 11220
rect 12040 11190 12080 11220
rect 12160 11190 12200 11220
rect 12280 11190 12320 11220
rect 12400 11190 12440 11220
rect 12520 11190 12560 11220
rect 12640 11190 12680 11220
rect 12760 11190 12800 11220
rect 12880 11190 12920 11220
rect 13640 11190 13680 11220
rect 13760 11190 13800 11220
rect 13880 11190 13920 11220
rect 14000 11190 14040 11220
rect 14120 11190 14160 11220
rect 14240 11190 14280 11220
rect 14360 11190 14400 11220
rect 14480 11190 14520 11220
rect 14600 11190 14640 11220
rect 14720 11190 14760 11220
rect 14840 11190 14880 11220
rect 14960 11190 15000 11220
rect 15080 11190 15120 11220
rect 15200 11190 15240 11220
rect 15320 11190 15360 11220
rect 15440 11190 15480 11220
rect 15560 11190 15600 11220
rect 15680 11190 15720 11220
rect 15800 11190 15840 11220
rect 15920 11190 15960 11220
rect 10530 11170 10640 11190
rect 10530 11130 10540 11170
rect 10580 11160 10640 11170
rect 12880 11170 12990 11190
rect 12880 11160 12940 11170
rect 10580 11130 10590 11160
rect 10530 11110 10590 11130
rect 12930 11130 12940 11160
rect 12980 11130 12990 11170
rect 12930 11110 12990 11130
rect 13570 11170 13680 11190
rect 13570 11130 13580 11170
rect 13620 11160 13680 11170
rect 15920 11170 16030 11190
rect 15920 11160 15980 11170
rect 13620 11130 13630 11160
rect 13570 11110 13630 11130
rect 15970 11130 15980 11160
rect 16020 11130 16030 11170
rect 15970 11110 16030 11130
rect 11900 10350 11970 10370
rect 11900 10310 11910 10350
rect 11950 10310 11970 10350
rect 11900 10290 11970 10310
rect 12070 10350 12150 10370
rect 12070 10310 12090 10350
rect 12130 10310 12150 10350
rect 12070 10290 12150 10310
rect 12250 10350 12330 10370
rect 12250 10310 12270 10350
rect 12310 10310 12330 10350
rect 12250 10290 12330 10310
rect 12430 10350 12510 10370
rect 12430 10310 12450 10350
rect 12490 10310 12510 10350
rect 12430 10290 12510 10310
rect 12610 10350 12690 10370
rect 12610 10310 12630 10350
rect 12670 10310 12690 10350
rect 12610 10290 12690 10310
rect 12790 10350 12870 10370
rect 12790 10310 12810 10350
rect 12850 10310 12870 10350
rect 12790 10290 12870 10310
rect 12970 10350 13050 10370
rect 12970 10310 12990 10350
rect 13030 10310 13050 10350
rect 12970 10290 13050 10310
rect 13150 10350 13220 10370
rect 13150 10310 13170 10350
rect 13210 10310 13220 10350
rect 13150 10290 13220 10310
rect 13340 10350 13410 10370
rect 13340 10310 13350 10350
rect 13390 10310 13410 10350
rect 13340 10290 13410 10310
rect 13510 10350 13590 10370
rect 13510 10310 13530 10350
rect 13570 10310 13590 10350
rect 13510 10290 13590 10310
rect 13690 10350 13770 10370
rect 13690 10310 13710 10350
rect 13750 10310 13770 10350
rect 13690 10290 13770 10310
rect 13870 10350 13950 10370
rect 13870 10310 13890 10350
rect 13930 10310 13950 10350
rect 13870 10290 13950 10310
rect 14050 10350 14130 10370
rect 14050 10310 14070 10350
rect 14110 10310 14130 10350
rect 14050 10290 14130 10310
rect 14230 10350 14310 10370
rect 14230 10310 14250 10350
rect 14290 10310 14310 10350
rect 14230 10290 14310 10310
rect 14410 10350 14490 10370
rect 14410 10310 14430 10350
rect 14470 10310 14490 10350
rect 14410 10290 14490 10310
rect 14590 10350 14660 10370
rect 14590 10310 14610 10350
rect 14650 10310 14660 10350
rect 14590 10300 14660 10310
rect 11700 10260 11800 10290
rect 11880 10260 11980 10290
rect 12060 10260 12160 10290
rect 12240 10260 12340 10290
rect 12420 10260 12520 10290
rect 12600 10260 12700 10290
rect 12780 10260 12880 10290
rect 12960 10260 13060 10290
rect 13140 10260 13240 10290
rect 13320 10260 13420 10290
rect 13500 10260 13600 10290
rect 13680 10260 13780 10290
rect 13860 10260 13960 10290
rect 14040 10260 14140 10290
rect 14220 10260 14320 10290
rect 14400 10260 14500 10290
rect 14580 10260 14680 10300
rect 14760 10260 14860 10290
rect 15710 10150 15790 10170
rect 15710 10110 15730 10150
rect 15770 10110 15790 10150
rect 15570 10060 15600 10090
rect 15680 10080 15820 10110
rect 15680 10060 15710 10080
rect 15790 10060 15820 10080
rect 15900 10060 15930 10090
rect 15570 9840 15600 9860
rect 15500 9810 15600 9840
rect 15680 9830 15710 9860
rect 15790 9830 15820 9860
rect 15900 9840 15930 9860
rect 15900 9810 16000 9840
rect 15500 9770 15510 9810
rect 15550 9770 15560 9810
rect 15500 9750 15560 9770
rect 15940 9770 15950 9810
rect 15990 9770 16000 9810
rect 15940 9750 16000 9770
rect 11700 9630 11800 9660
rect 11880 9630 11980 9660
rect 12060 9630 12160 9660
rect 12240 9630 12340 9660
rect 12420 9630 12520 9660
rect 12600 9630 12700 9660
rect 12780 9630 12880 9660
rect 12960 9630 13060 9660
rect 13140 9630 13240 9660
rect 13320 9630 13420 9660
rect 13500 9630 13600 9660
rect 13680 9630 13780 9660
rect 13860 9630 13960 9660
rect 14040 9630 14140 9660
rect 14220 9630 14320 9660
rect 14400 9630 14500 9660
rect 14580 9630 14680 9660
rect 14760 9630 14860 9660
rect 11620 9610 11800 9630
rect 11620 9570 11640 9610
rect 11680 9600 11800 9610
rect 14760 9610 14940 9630
rect 14760 9600 14880 9610
rect 11680 9570 11700 9600
rect 11620 9550 11700 9570
rect 14860 9570 14880 9600
rect 14920 9570 14940 9610
rect 14860 9550 14940 9570
rect 11806 9342 11864 9360
rect 11806 9308 11818 9342
rect 11852 9308 11864 9342
rect 11806 9290 11864 9308
rect 11916 9342 11974 9360
rect 11916 9308 11928 9342
rect 11962 9308 11974 9342
rect 11916 9290 11974 9308
rect 12026 9342 12084 9360
rect 12026 9308 12038 9342
rect 12072 9308 12084 9342
rect 12026 9290 12084 9308
rect 12136 9342 12194 9360
rect 12136 9308 12148 9342
rect 12182 9308 12194 9342
rect 12136 9290 12194 9308
rect 12246 9342 12304 9360
rect 12246 9308 12258 9342
rect 12292 9308 12304 9342
rect 12246 9290 12304 9308
rect 12356 9342 12414 9360
rect 12356 9308 12368 9342
rect 12402 9308 12414 9342
rect 12356 9290 12414 9308
rect 12466 9342 12524 9360
rect 12466 9308 12478 9342
rect 12512 9308 12524 9342
rect 12466 9290 12524 9308
rect 12576 9342 12634 9360
rect 12576 9308 12588 9342
rect 12622 9308 12634 9342
rect 12576 9290 12634 9308
rect 12686 9342 12744 9360
rect 12686 9308 12698 9342
rect 12732 9308 12744 9342
rect 12686 9290 12744 9308
rect 12796 9342 12854 9360
rect 12796 9308 12808 9342
rect 12842 9308 12854 9342
rect 12796 9290 12854 9308
rect 13706 9342 13764 9360
rect 13706 9308 13718 9342
rect 13752 9308 13764 9342
rect 13706 9290 13764 9308
rect 13816 9342 13874 9360
rect 13816 9308 13828 9342
rect 13862 9308 13874 9342
rect 13816 9290 13874 9308
rect 13926 9342 13984 9360
rect 13926 9308 13938 9342
rect 13972 9308 13984 9342
rect 13926 9290 13984 9308
rect 14036 9342 14094 9360
rect 14036 9308 14048 9342
rect 14082 9308 14094 9342
rect 14036 9290 14094 9308
rect 14146 9342 14204 9360
rect 14146 9308 14158 9342
rect 14192 9308 14204 9342
rect 14146 9290 14204 9308
rect 14256 9342 14314 9360
rect 14256 9308 14268 9342
rect 14302 9308 14314 9342
rect 14256 9290 14314 9308
rect 14366 9342 14424 9360
rect 14366 9308 14378 9342
rect 14412 9308 14424 9342
rect 14366 9290 14424 9308
rect 14476 9342 14534 9360
rect 14476 9308 14488 9342
rect 14522 9308 14534 9342
rect 14476 9290 14534 9308
rect 14586 9342 14644 9360
rect 14586 9308 14598 9342
rect 14632 9308 14644 9342
rect 14586 9290 14644 9308
rect 14696 9342 14754 9360
rect 14696 9308 14708 9342
rect 14742 9308 14754 9342
rect 14696 9290 14754 9308
rect 11710 9260 11740 9290
rect 11820 9260 11850 9290
rect 11930 9260 11960 9290
rect 12040 9260 12070 9290
rect 12150 9260 12180 9290
rect 12260 9260 12290 9290
rect 12370 9260 12400 9290
rect 12480 9260 12510 9290
rect 12590 9260 12620 9290
rect 12700 9260 12730 9290
rect 12810 9260 12840 9290
rect 12920 9260 12950 9290
rect 13610 9260 13640 9290
rect 13720 9260 13750 9290
rect 13830 9260 13860 9290
rect 13940 9260 13970 9290
rect 14050 9260 14080 9290
rect 14160 9260 14190 9290
rect 14270 9260 14300 9290
rect 14380 9260 14410 9290
rect 14490 9260 14520 9290
rect 14600 9260 14630 9290
rect 14710 9260 14740 9290
rect 14820 9260 14850 9290
rect 11710 9030 11740 9060
rect 11820 9030 11850 9060
rect 11930 9030 11960 9060
rect 12040 9030 12070 9060
rect 12150 9030 12180 9060
rect 12260 9030 12290 9060
rect 12370 9030 12400 9060
rect 12480 9030 12510 9060
rect 12590 9030 12620 9060
rect 12700 9030 12730 9060
rect 12810 9030 12840 9060
rect 12920 9030 12950 9060
rect 13610 9030 13640 9060
rect 13720 9030 13750 9060
rect 13830 9030 13860 9060
rect 13940 9030 13970 9060
rect 14050 9030 14080 9060
rect 14160 9030 14190 9060
rect 14270 9030 14300 9060
rect 14380 9030 14410 9060
rect 14490 9030 14520 9060
rect 14600 9030 14630 9060
rect 14710 9030 14740 9060
rect 14820 9030 14850 9060
rect 11630 9010 11740 9030
rect 11630 8970 11650 9010
rect 11690 9000 11740 9010
rect 12920 9010 13030 9030
rect 12920 9000 12970 9010
rect 11690 8970 11710 9000
rect 11630 8950 11710 8970
rect 12950 8970 12970 9000
rect 13010 8970 13030 9010
rect 12950 8950 13030 8970
rect 13530 9010 13640 9030
rect 13530 8970 13550 9010
rect 13590 9000 13640 9010
rect 14820 9010 14930 9030
rect 14820 9000 14870 9010
rect 13590 8970 13610 9000
rect 13530 8950 13610 8970
rect 14850 8970 14870 9000
rect 14910 8970 14930 9010
rect 14850 8950 14930 8970
<< polycont >>
rect 11340 13590 11380 13630
rect 11500 13590 11540 13630
rect 11660 13590 11700 13630
rect 11820 13590 11860 13630
rect 11980 13590 12020 13630
rect 12140 13590 12180 13630
rect 12300 13590 12340 13630
rect 12460 13590 12500 13630
rect 12620 13590 12660 13630
rect 12780 13590 12820 13630
rect 12940 13590 12980 13630
rect 13100 13590 13140 13630
rect 13420 13590 13460 13630
rect 13580 13590 13620 13630
rect 13740 13590 13780 13630
rect 13900 13590 13940 13630
rect 14060 13590 14100 13630
rect 14220 13590 14260 13630
rect 14380 13590 14420 13630
rect 14540 13590 14580 13630
rect 14700 13590 14740 13630
rect 14860 13590 14900 13630
rect 15020 13590 15060 13630
rect 15180 13590 15220 13630
rect 10940 12680 10980 12720
rect 11180 12680 11220 12720
rect 11420 12680 11460 12720
rect 11660 12680 11700 12720
rect 12300 12680 12340 12720
rect 12540 12680 12580 12720
rect 12780 12680 12820 12720
rect 13740 12680 13780 12720
rect 13980 12680 14020 12720
rect 14220 12680 14260 12720
rect 14860 12680 14900 12720
rect 15100 12680 15140 12720
rect 15340 12680 15380 12720
rect 15580 12680 15620 12720
rect 11443 12308 11477 12342
rect 11803 12308 11837 12342
rect 11923 12308 11957 12342
rect 12283 12308 12317 12342
rect 12403 12308 12437 12342
rect 11544 12078 11578 12112
rect 11702 12078 11736 12112
rect 12026 12078 12060 12112
rect 12180 12078 12214 12112
rect 12504 12078 12538 12112
rect 14123 12308 14157 12342
rect 14243 12308 14277 12342
rect 14603 12308 14637 12342
rect 14723 12308 14757 12342
rect 15083 12308 15117 12342
rect 14022 12078 14056 12112
rect 14346 12078 14380 12112
rect 14500 12078 14534 12112
rect 14824 12078 14858 12112
rect 14982 12078 15016 12112
rect 10720 11480 10760 11520
rect 10900 11470 10940 11510
rect 11380 11470 11420 11510
rect 11620 11470 11660 11510
rect 12100 11470 12140 11510
rect 12340 11470 12380 11510
rect 12760 11470 12800 11510
rect 13760 11470 13800 11510
rect 14180 11470 14220 11510
rect 14420 11470 14460 11510
rect 14900 11470 14940 11510
rect 15140 11470 15180 11510
rect 15620 11470 15660 11510
rect 15800 11480 15840 11520
rect 10540 11130 10580 11170
rect 12940 11130 12980 11170
rect 13580 11130 13620 11170
rect 15980 11130 16020 11170
rect 11910 10310 11950 10350
rect 12090 10310 12130 10350
rect 12270 10310 12310 10350
rect 12450 10310 12490 10350
rect 12630 10310 12670 10350
rect 12810 10310 12850 10350
rect 12990 10310 13030 10350
rect 13170 10310 13210 10350
rect 13350 10310 13390 10350
rect 13530 10310 13570 10350
rect 13710 10310 13750 10350
rect 13890 10310 13930 10350
rect 14070 10310 14110 10350
rect 14250 10310 14290 10350
rect 14430 10310 14470 10350
rect 14610 10310 14650 10350
rect 15730 10110 15770 10150
rect 15510 9770 15550 9810
rect 15950 9770 15990 9810
rect 11640 9570 11680 9610
rect 14880 9570 14920 9610
rect 11818 9308 11852 9342
rect 11928 9308 11962 9342
rect 12038 9308 12072 9342
rect 12148 9308 12182 9342
rect 12258 9308 12292 9342
rect 12368 9308 12402 9342
rect 12478 9308 12512 9342
rect 12588 9308 12622 9342
rect 12698 9308 12732 9342
rect 12808 9308 12842 9342
rect 13718 9308 13752 9342
rect 13828 9308 13862 9342
rect 13938 9308 13972 9342
rect 14048 9308 14082 9342
rect 14158 9308 14192 9342
rect 14268 9308 14302 9342
rect 14378 9308 14412 9342
rect 14488 9308 14522 9342
rect 14598 9308 14632 9342
rect 14708 9308 14742 9342
rect 11650 8970 11690 9010
rect 12970 8970 13010 9010
rect 13550 8970 13590 9010
rect 14870 8970 14910 9010
<< xpolycontact >>
rect 8760 18018 8898 18450
rect 8760 16632 8898 17064
rect 9574 18024 9644 18456
rect 9574 15062 9644 15494
rect 10686 18026 10756 18458
rect 10354 16286 10424 16718
rect 15674 18026 15744 18458
rect 16006 16286 16076 16718
rect 16784 18024 16854 18456
rect 16784 15952 16854 16384
rect 17540 18018 17678 18450
rect 17540 16632 17678 17064
rect 11542 14344 11974 14414
rect 14582 14344 15014 14414
<< ppolyres >>
rect 8760 17064 8898 18018
rect 16784 16384 16854 18024
rect 17540 17064 17678 18018
rect 11974 14344 14582 14414
<< xpolyres >>
rect 9574 15494 9644 18024
rect 10354 17852 10590 17922
rect 10354 16718 10424 17852
rect 10520 16892 10590 17852
rect 10686 16892 10756 18026
rect 10520 16822 10756 16892
rect 15674 16892 15744 18026
rect 15840 17852 16076 17922
rect 15840 16892 15910 17852
rect 15674 16822 15910 16892
rect 16006 16718 16076 17852
<< locali >>
rect 13240 19070 13320 19090
rect 13240 19030 13260 19070
rect 13300 19030 13320 19070
rect 13240 18990 13320 19030
rect 13240 18950 13260 18990
rect 13300 18950 13320 18990
rect 13240 18910 13320 18950
rect 13240 18870 13260 18910
rect 13300 18870 13320 18910
rect 12560 18784 12640 18790
rect 13240 18784 13320 18870
rect 13920 18784 14000 18790
rect 11276 18752 15284 18784
rect 11276 18718 11410 18752
rect 11444 18718 11500 18752
rect 11534 18718 11590 18752
rect 11624 18718 11680 18752
rect 11714 18718 11770 18752
rect 11804 18718 11860 18752
rect 11894 18718 11950 18752
rect 11984 18718 12040 18752
rect 12074 18718 12130 18752
rect 12164 18718 12220 18752
rect 12254 18718 12310 18752
rect 12344 18718 12400 18752
rect 12434 18718 12770 18752
rect 12804 18718 12860 18752
rect 12894 18718 12950 18752
rect 12984 18718 13040 18752
rect 13074 18718 13130 18752
rect 13164 18718 13220 18752
rect 13254 18718 13310 18752
rect 13344 18718 13400 18752
rect 13434 18718 13490 18752
rect 13524 18718 13580 18752
rect 13614 18718 13670 18752
rect 13704 18718 13760 18752
rect 13794 18718 14130 18752
rect 14164 18718 14220 18752
rect 14254 18718 14310 18752
rect 14344 18718 14400 18752
rect 14434 18718 14490 18752
rect 14524 18718 14580 18752
rect 14614 18718 14670 18752
rect 14704 18718 14760 18752
rect 14794 18718 14850 18752
rect 14884 18718 14940 18752
rect 14974 18718 15030 18752
rect 15064 18718 15120 18752
rect 15154 18718 15284 18752
rect 11276 18685 15284 18718
rect 11276 18668 11375 18685
rect 11276 18634 11309 18668
rect 11343 18634 11375 18668
rect 8790 18590 8870 18610
rect 9570 18600 9650 18620
rect 9570 18595 9590 18600
rect 9630 18595 9650 18600
rect 10680 18610 10760 18630
rect 10680 18597 10700 18610
rect 10740 18597 10760 18610
rect 8790 18589 8810 18590
rect 8850 18589 8870 18590
rect 8603 18555 8699 18589
rect 8959 18555 9055 18589
rect 8603 18493 8637 18555
rect 8790 18550 8810 18555
rect 8850 18550 8870 18555
rect 8790 18530 8870 18550
rect 9021 18493 9055 18555
rect 8603 16527 8637 16589
rect 9021 16527 9055 16589
rect 8603 16493 8699 16527
rect 8959 16493 9055 16527
rect 9383 18561 9479 18595
rect 9739 18561 9835 18595
rect 9383 18499 9417 18561
rect 9570 18560 9590 18561
rect 9630 18560 9650 18561
rect 9570 18540 9650 18560
rect 9801 18499 9835 18561
rect 9383 14957 9417 15019
rect 10163 18563 10259 18597
rect 10851 18563 10947 18597
rect 10163 18501 10197 18563
rect 10680 18550 10760 18563
rect 10913 18501 10947 18563
rect 10163 16181 10197 16243
rect 11276 18578 11375 18634
rect 12465 18668 12735 18685
rect 12465 18634 12496 18668
rect 12530 18634 12669 18668
rect 12703 18634 12735 18668
rect 11276 18544 11309 18578
rect 11343 18544 11375 18578
rect 11276 18488 11375 18544
rect 11276 18454 11309 18488
rect 11343 18454 11375 18488
rect 11276 18398 11375 18454
rect 11276 18364 11309 18398
rect 11343 18364 11375 18398
rect 11276 18308 11375 18364
rect 11276 18274 11309 18308
rect 11343 18274 11375 18308
rect 11276 18218 11375 18274
rect 11276 18184 11309 18218
rect 11343 18184 11375 18218
rect 11276 18128 11375 18184
rect 11276 18094 11309 18128
rect 11343 18094 11375 18128
rect 11276 18038 11375 18094
rect 11276 18004 11309 18038
rect 11343 18004 11375 18038
rect 11276 17948 11375 18004
rect 11276 17914 11309 17948
rect 11343 17914 11375 17948
rect 11276 17858 11375 17914
rect 11276 17824 11309 17858
rect 11343 17824 11375 17858
rect 11276 17768 11375 17824
rect 11276 17740 11309 17768
rect 11270 17734 11309 17740
rect 11343 17740 11375 17768
rect 11439 18602 12401 18621
rect 11439 18568 11550 18602
rect 11584 18568 11640 18602
rect 11674 18568 11730 18602
rect 11764 18568 11820 18602
rect 11854 18568 11910 18602
rect 11944 18568 12000 18602
rect 12034 18568 12090 18602
rect 12124 18568 12180 18602
rect 12214 18568 12270 18602
rect 12304 18568 12401 18602
rect 11439 18549 12401 18568
rect 11439 18508 11511 18549
rect 11439 18474 11458 18508
rect 11492 18474 11511 18508
rect 12329 18489 12401 18549
rect 11439 18418 11511 18474
rect 11439 18384 11458 18418
rect 11492 18384 11511 18418
rect 11439 18328 11511 18384
rect 11439 18294 11458 18328
rect 11492 18294 11511 18328
rect 11439 18238 11511 18294
rect 11439 18204 11458 18238
rect 11492 18204 11511 18238
rect 11439 18148 11511 18204
rect 11439 18114 11458 18148
rect 11492 18114 11511 18148
rect 11439 18058 11511 18114
rect 11439 18024 11458 18058
rect 11492 18024 11511 18058
rect 11439 17968 11511 18024
rect 11439 17934 11458 17968
rect 11492 17934 11511 17968
rect 11439 17878 11511 17934
rect 11439 17844 11458 17878
rect 11492 17844 11511 17878
rect 11439 17788 11511 17844
rect 11573 18426 12267 18487
rect 11573 18392 11632 18426
rect 11666 18414 11722 18426
rect 11694 18392 11722 18414
rect 11756 18414 11812 18426
rect 11756 18392 11760 18414
rect 11573 18380 11660 18392
rect 11694 18380 11760 18392
rect 11794 18392 11812 18414
rect 11846 18414 11902 18426
rect 11846 18392 11860 18414
rect 11794 18380 11860 18392
rect 11894 18392 11902 18414
rect 11936 18414 11992 18426
rect 12026 18414 12082 18426
rect 12116 18414 12172 18426
rect 11936 18392 11960 18414
rect 12026 18392 12060 18414
rect 12116 18392 12160 18414
rect 12206 18392 12267 18426
rect 11894 18380 11960 18392
rect 11994 18380 12060 18392
rect 12094 18380 12160 18392
rect 12194 18380 12267 18392
rect 11573 18336 12267 18380
rect 11573 18302 11632 18336
rect 11666 18314 11722 18336
rect 11694 18302 11722 18314
rect 11756 18314 11812 18336
rect 11756 18302 11760 18314
rect 11573 18280 11660 18302
rect 11694 18280 11760 18302
rect 11794 18302 11812 18314
rect 11846 18314 11902 18336
rect 11846 18302 11860 18314
rect 11794 18280 11860 18302
rect 11894 18302 11902 18314
rect 11936 18314 11992 18336
rect 12026 18314 12082 18336
rect 12116 18314 12172 18336
rect 11936 18302 11960 18314
rect 12026 18302 12060 18314
rect 12116 18302 12160 18314
rect 12206 18302 12267 18336
rect 11894 18280 11960 18302
rect 11994 18280 12060 18302
rect 12094 18280 12160 18302
rect 12194 18280 12267 18302
rect 11573 18246 12267 18280
rect 11573 18212 11632 18246
rect 11666 18214 11722 18246
rect 11694 18212 11722 18214
rect 11756 18214 11812 18246
rect 11756 18212 11760 18214
rect 11573 18180 11660 18212
rect 11694 18180 11760 18212
rect 11794 18212 11812 18214
rect 11846 18214 11902 18246
rect 11846 18212 11860 18214
rect 11794 18180 11860 18212
rect 11894 18212 11902 18214
rect 11936 18214 11992 18246
rect 12026 18214 12082 18246
rect 12116 18214 12172 18246
rect 11936 18212 11960 18214
rect 12026 18212 12060 18214
rect 12116 18212 12160 18214
rect 12206 18212 12267 18246
rect 11894 18180 11960 18212
rect 11994 18180 12060 18212
rect 12094 18180 12160 18212
rect 12194 18180 12267 18212
rect 11573 18156 12267 18180
rect 11573 18122 11632 18156
rect 11666 18122 11722 18156
rect 11756 18122 11812 18156
rect 11846 18122 11902 18156
rect 11936 18122 11992 18156
rect 12026 18122 12082 18156
rect 12116 18122 12172 18156
rect 12206 18122 12267 18156
rect 11573 18114 12267 18122
rect 11573 18080 11660 18114
rect 11694 18080 11760 18114
rect 11794 18080 11860 18114
rect 11894 18080 11960 18114
rect 11994 18080 12060 18114
rect 12094 18080 12160 18114
rect 12194 18080 12267 18114
rect 11573 18066 12267 18080
rect 11573 18032 11632 18066
rect 11666 18032 11722 18066
rect 11756 18032 11812 18066
rect 11846 18032 11902 18066
rect 11936 18032 11992 18066
rect 12026 18032 12082 18066
rect 12116 18032 12172 18066
rect 12206 18032 12267 18066
rect 11573 18014 12267 18032
rect 11573 17980 11660 18014
rect 11694 17980 11760 18014
rect 11794 17980 11860 18014
rect 11894 17980 11960 18014
rect 11994 17980 12060 18014
rect 12094 17980 12160 18014
rect 12194 17980 12267 18014
rect 11573 17976 12267 17980
rect 11573 17942 11632 17976
rect 11666 17942 11722 17976
rect 11756 17942 11812 17976
rect 11846 17942 11902 17976
rect 11936 17942 11992 17976
rect 12026 17942 12082 17976
rect 12116 17942 12172 17976
rect 12206 17942 12267 17976
rect 11573 17914 12267 17942
rect 11573 17886 11660 17914
rect 11694 17886 11760 17914
rect 11573 17852 11632 17886
rect 11694 17880 11722 17886
rect 11666 17852 11722 17880
rect 11756 17880 11760 17886
rect 11794 17886 11860 17914
rect 11794 17880 11812 17886
rect 11756 17852 11812 17880
rect 11846 17880 11860 17886
rect 11894 17886 11960 17914
rect 11994 17886 12060 17914
rect 12094 17886 12160 17914
rect 12194 17886 12267 17914
rect 11894 17880 11902 17886
rect 11846 17852 11902 17880
rect 11936 17880 11960 17886
rect 12026 17880 12060 17886
rect 12116 17880 12160 17886
rect 11936 17852 11992 17880
rect 12026 17852 12082 17880
rect 12116 17852 12172 17880
rect 12206 17852 12267 17886
rect 11573 17793 12267 17852
rect 12329 18455 12348 18489
rect 12382 18455 12401 18489
rect 12329 18399 12401 18455
rect 12329 18365 12348 18399
rect 12382 18365 12401 18399
rect 12329 18309 12401 18365
rect 12329 18275 12348 18309
rect 12382 18275 12401 18309
rect 12329 18219 12401 18275
rect 12329 18185 12348 18219
rect 12382 18185 12401 18219
rect 12329 18129 12401 18185
rect 12329 18095 12348 18129
rect 12382 18095 12401 18129
rect 12329 18039 12401 18095
rect 12329 18005 12348 18039
rect 12382 18005 12401 18039
rect 12329 17949 12401 18005
rect 12329 17915 12348 17949
rect 12382 17915 12401 17949
rect 12329 17859 12401 17915
rect 12329 17825 12348 17859
rect 12382 17825 12401 17859
rect 11439 17754 11458 17788
rect 11492 17754 11511 17788
rect 11439 17740 11511 17754
rect 12329 17769 12401 17825
rect 12329 17740 12348 17769
rect 11343 17735 12348 17740
rect 12382 17740 12401 17769
rect 12465 18578 12735 18634
rect 13825 18668 14095 18685
rect 13825 18634 13856 18668
rect 13890 18634 14029 18668
rect 14063 18634 14095 18668
rect 12465 18544 12496 18578
rect 12530 18544 12669 18578
rect 12703 18544 12735 18578
rect 12465 18488 12735 18544
rect 12465 18454 12496 18488
rect 12530 18454 12669 18488
rect 12703 18454 12735 18488
rect 12465 18398 12735 18454
rect 12465 18364 12496 18398
rect 12530 18364 12669 18398
rect 12703 18364 12735 18398
rect 12465 18308 12735 18364
rect 12465 18274 12496 18308
rect 12530 18274 12669 18308
rect 12703 18274 12735 18308
rect 12465 18218 12735 18274
rect 12465 18184 12496 18218
rect 12530 18184 12669 18218
rect 12703 18184 12735 18218
rect 12465 18128 12735 18184
rect 12465 18094 12496 18128
rect 12530 18094 12669 18128
rect 12703 18094 12735 18128
rect 12465 18038 12735 18094
rect 12465 18004 12496 18038
rect 12530 18004 12669 18038
rect 12703 18004 12735 18038
rect 12465 17948 12735 18004
rect 12465 17914 12496 17948
rect 12530 17914 12669 17948
rect 12703 17914 12735 17948
rect 12465 17858 12735 17914
rect 12465 17824 12496 17858
rect 12530 17824 12669 17858
rect 12703 17824 12735 17858
rect 12465 17768 12735 17824
rect 12465 17740 12496 17768
rect 12382 17735 12496 17740
rect 11343 17734 12496 17735
rect 12530 17734 12669 17768
rect 12703 17740 12735 17768
rect 12799 18602 13761 18621
rect 12799 18568 12910 18602
rect 12944 18568 13000 18602
rect 13034 18568 13090 18602
rect 13124 18568 13180 18602
rect 13214 18568 13270 18602
rect 13304 18568 13360 18602
rect 13394 18568 13450 18602
rect 13484 18568 13540 18602
rect 13574 18568 13630 18602
rect 13664 18568 13761 18602
rect 12799 18549 13761 18568
rect 12799 18508 12871 18549
rect 12799 18474 12818 18508
rect 12852 18474 12871 18508
rect 13689 18489 13761 18549
rect 12799 18418 12871 18474
rect 12799 18384 12818 18418
rect 12852 18384 12871 18418
rect 12799 18328 12871 18384
rect 12799 18294 12818 18328
rect 12852 18294 12871 18328
rect 12799 18238 12871 18294
rect 12799 18204 12818 18238
rect 12852 18204 12871 18238
rect 12799 18148 12871 18204
rect 12799 18114 12818 18148
rect 12852 18114 12871 18148
rect 12799 18058 12871 18114
rect 12799 18024 12818 18058
rect 12852 18024 12871 18058
rect 12799 17968 12871 18024
rect 12799 17934 12818 17968
rect 12852 17934 12871 17968
rect 12799 17878 12871 17934
rect 12799 17844 12818 17878
rect 12852 17844 12871 17878
rect 12799 17788 12871 17844
rect 12933 18426 13627 18487
rect 12933 18392 12992 18426
rect 13026 18414 13082 18426
rect 13054 18392 13082 18414
rect 13116 18414 13172 18426
rect 13116 18392 13120 18414
rect 12933 18380 13020 18392
rect 13054 18380 13120 18392
rect 13154 18392 13172 18414
rect 13206 18414 13262 18426
rect 13206 18392 13220 18414
rect 13154 18380 13220 18392
rect 13254 18392 13262 18414
rect 13296 18414 13352 18426
rect 13386 18414 13442 18426
rect 13476 18414 13532 18426
rect 13296 18392 13320 18414
rect 13386 18392 13420 18414
rect 13476 18392 13520 18414
rect 13566 18392 13627 18426
rect 13254 18380 13320 18392
rect 13354 18380 13420 18392
rect 13454 18380 13520 18392
rect 13554 18380 13627 18392
rect 12933 18336 13627 18380
rect 12933 18302 12992 18336
rect 13026 18314 13082 18336
rect 13054 18302 13082 18314
rect 13116 18314 13172 18336
rect 13116 18302 13120 18314
rect 12933 18280 13020 18302
rect 13054 18280 13120 18302
rect 13154 18302 13172 18314
rect 13206 18314 13262 18336
rect 13206 18302 13220 18314
rect 13154 18280 13220 18302
rect 13254 18302 13262 18314
rect 13296 18314 13352 18336
rect 13386 18314 13442 18336
rect 13476 18314 13532 18336
rect 13296 18302 13320 18314
rect 13386 18302 13420 18314
rect 13476 18302 13520 18314
rect 13566 18302 13627 18336
rect 13254 18280 13320 18302
rect 13354 18280 13420 18302
rect 13454 18280 13520 18302
rect 13554 18280 13627 18302
rect 12933 18246 13627 18280
rect 12933 18212 12992 18246
rect 13026 18214 13082 18246
rect 13054 18212 13082 18214
rect 13116 18214 13172 18246
rect 13116 18212 13120 18214
rect 12933 18180 13020 18212
rect 13054 18180 13120 18212
rect 13154 18212 13172 18214
rect 13206 18214 13262 18246
rect 13206 18212 13220 18214
rect 13154 18180 13220 18212
rect 13254 18212 13262 18214
rect 13296 18214 13352 18246
rect 13386 18214 13442 18246
rect 13476 18214 13532 18246
rect 13296 18212 13320 18214
rect 13386 18212 13420 18214
rect 13476 18212 13520 18214
rect 13566 18212 13627 18246
rect 13254 18180 13320 18212
rect 13354 18180 13420 18212
rect 13454 18180 13520 18212
rect 13554 18180 13627 18212
rect 12933 18156 13627 18180
rect 12933 18122 12992 18156
rect 13026 18122 13082 18156
rect 13116 18122 13172 18156
rect 13206 18122 13262 18156
rect 13296 18122 13352 18156
rect 13386 18122 13442 18156
rect 13476 18122 13532 18156
rect 13566 18122 13627 18156
rect 12933 18114 13627 18122
rect 12933 18080 13020 18114
rect 13054 18080 13120 18114
rect 13154 18080 13220 18114
rect 13254 18080 13320 18114
rect 13354 18080 13420 18114
rect 13454 18080 13520 18114
rect 13554 18080 13627 18114
rect 12933 18066 13627 18080
rect 12933 18032 12992 18066
rect 13026 18032 13082 18066
rect 13116 18032 13172 18066
rect 13206 18032 13262 18066
rect 13296 18032 13352 18066
rect 13386 18032 13442 18066
rect 13476 18032 13532 18066
rect 13566 18032 13627 18066
rect 12933 18014 13627 18032
rect 12933 17980 13020 18014
rect 13054 17980 13120 18014
rect 13154 17980 13220 18014
rect 13254 17980 13320 18014
rect 13354 17980 13420 18014
rect 13454 17980 13520 18014
rect 13554 17980 13627 18014
rect 12933 17976 13627 17980
rect 12933 17942 12992 17976
rect 13026 17942 13082 17976
rect 13116 17942 13172 17976
rect 13206 17942 13262 17976
rect 13296 17942 13352 17976
rect 13386 17942 13442 17976
rect 13476 17942 13532 17976
rect 13566 17942 13627 17976
rect 12933 17914 13627 17942
rect 12933 17886 13020 17914
rect 13054 17886 13120 17914
rect 12933 17852 12992 17886
rect 13054 17880 13082 17886
rect 13026 17852 13082 17880
rect 13116 17880 13120 17886
rect 13154 17886 13220 17914
rect 13154 17880 13172 17886
rect 13116 17852 13172 17880
rect 13206 17880 13220 17886
rect 13254 17886 13320 17914
rect 13354 17886 13420 17914
rect 13454 17886 13520 17914
rect 13554 17886 13627 17914
rect 13254 17880 13262 17886
rect 13206 17852 13262 17880
rect 13296 17880 13320 17886
rect 13386 17880 13420 17886
rect 13476 17880 13520 17886
rect 13296 17852 13352 17880
rect 13386 17852 13442 17880
rect 13476 17852 13532 17880
rect 13566 17852 13627 17886
rect 12933 17793 13627 17852
rect 13689 18455 13708 18489
rect 13742 18455 13761 18489
rect 13689 18399 13761 18455
rect 13689 18365 13708 18399
rect 13742 18365 13761 18399
rect 13689 18309 13761 18365
rect 13689 18275 13708 18309
rect 13742 18275 13761 18309
rect 13689 18219 13761 18275
rect 13689 18185 13708 18219
rect 13742 18185 13761 18219
rect 13689 18129 13761 18185
rect 13689 18095 13708 18129
rect 13742 18095 13761 18129
rect 13689 18039 13761 18095
rect 13689 18005 13708 18039
rect 13742 18005 13761 18039
rect 13689 17949 13761 18005
rect 13689 17915 13708 17949
rect 13742 17915 13761 17949
rect 13689 17859 13761 17915
rect 13689 17825 13708 17859
rect 13742 17825 13761 17859
rect 12799 17754 12818 17788
rect 12852 17754 12871 17788
rect 12799 17740 12871 17754
rect 13689 17769 13761 17825
rect 13689 17740 13708 17769
rect 12703 17735 13708 17740
rect 13742 17740 13761 17769
rect 13825 18578 14095 18634
rect 15185 18668 15284 18685
rect 15185 18634 15216 18668
rect 15250 18634 15284 18668
rect 13825 18544 13856 18578
rect 13890 18544 14029 18578
rect 14063 18544 14095 18578
rect 13825 18488 14095 18544
rect 13825 18454 13856 18488
rect 13890 18454 14029 18488
rect 14063 18454 14095 18488
rect 13825 18398 14095 18454
rect 13825 18364 13856 18398
rect 13890 18364 14029 18398
rect 14063 18364 14095 18398
rect 13825 18308 14095 18364
rect 13825 18274 13856 18308
rect 13890 18274 14029 18308
rect 14063 18274 14095 18308
rect 13825 18218 14095 18274
rect 13825 18184 13856 18218
rect 13890 18184 14029 18218
rect 14063 18184 14095 18218
rect 13825 18128 14095 18184
rect 13825 18094 13856 18128
rect 13890 18094 14029 18128
rect 14063 18094 14095 18128
rect 13825 18038 14095 18094
rect 13825 18004 13856 18038
rect 13890 18004 14029 18038
rect 14063 18004 14095 18038
rect 13825 17948 14095 18004
rect 13825 17914 13856 17948
rect 13890 17914 14029 17948
rect 14063 17914 14095 17948
rect 13825 17858 14095 17914
rect 13825 17824 13856 17858
rect 13890 17824 14029 17858
rect 14063 17824 14095 17858
rect 13825 17768 14095 17824
rect 13825 17740 13856 17768
rect 13742 17735 13856 17740
rect 12703 17734 13856 17735
rect 13890 17734 14029 17768
rect 14063 17740 14095 17768
rect 14159 18602 15121 18621
rect 14159 18568 14270 18602
rect 14304 18568 14360 18602
rect 14394 18568 14450 18602
rect 14484 18568 14540 18602
rect 14574 18568 14630 18602
rect 14664 18568 14720 18602
rect 14754 18568 14810 18602
rect 14844 18568 14900 18602
rect 14934 18568 14990 18602
rect 15024 18568 15121 18602
rect 14159 18549 15121 18568
rect 14159 18508 14231 18549
rect 14159 18474 14178 18508
rect 14212 18474 14231 18508
rect 15049 18489 15121 18549
rect 14159 18418 14231 18474
rect 14159 18384 14178 18418
rect 14212 18384 14231 18418
rect 14159 18328 14231 18384
rect 14159 18294 14178 18328
rect 14212 18294 14231 18328
rect 14159 18238 14231 18294
rect 14159 18204 14178 18238
rect 14212 18204 14231 18238
rect 14159 18148 14231 18204
rect 14159 18114 14178 18148
rect 14212 18114 14231 18148
rect 14159 18058 14231 18114
rect 14159 18024 14178 18058
rect 14212 18024 14231 18058
rect 14159 17968 14231 18024
rect 14159 17934 14178 17968
rect 14212 17934 14231 17968
rect 14159 17878 14231 17934
rect 14159 17844 14178 17878
rect 14212 17844 14231 17878
rect 14159 17788 14231 17844
rect 14293 18426 14987 18487
rect 14293 18392 14352 18426
rect 14386 18414 14442 18426
rect 14414 18392 14442 18414
rect 14476 18414 14532 18426
rect 14476 18392 14480 18414
rect 14293 18380 14380 18392
rect 14414 18380 14480 18392
rect 14514 18392 14532 18414
rect 14566 18414 14622 18426
rect 14566 18392 14580 18414
rect 14514 18380 14580 18392
rect 14614 18392 14622 18414
rect 14656 18414 14712 18426
rect 14746 18414 14802 18426
rect 14836 18414 14892 18426
rect 14656 18392 14680 18414
rect 14746 18392 14780 18414
rect 14836 18392 14880 18414
rect 14926 18392 14987 18426
rect 14614 18380 14680 18392
rect 14714 18380 14780 18392
rect 14814 18380 14880 18392
rect 14914 18380 14987 18392
rect 14293 18336 14987 18380
rect 14293 18302 14352 18336
rect 14386 18314 14442 18336
rect 14414 18302 14442 18314
rect 14476 18314 14532 18336
rect 14476 18302 14480 18314
rect 14293 18280 14380 18302
rect 14414 18280 14480 18302
rect 14514 18302 14532 18314
rect 14566 18314 14622 18336
rect 14566 18302 14580 18314
rect 14514 18280 14580 18302
rect 14614 18302 14622 18314
rect 14656 18314 14712 18336
rect 14746 18314 14802 18336
rect 14836 18314 14892 18336
rect 14656 18302 14680 18314
rect 14746 18302 14780 18314
rect 14836 18302 14880 18314
rect 14926 18302 14987 18336
rect 14614 18280 14680 18302
rect 14714 18280 14780 18302
rect 14814 18280 14880 18302
rect 14914 18280 14987 18302
rect 14293 18246 14987 18280
rect 14293 18212 14352 18246
rect 14386 18214 14442 18246
rect 14414 18212 14442 18214
rect 14476 18214 14532 18246
rect 14476 18212 14480 18214
rect 14293 18180 14380 18212
rect 14414 18180 14480 18212
rect 14514 18212 14532 18214
rect 14566 18214 14622 18246
rect 14566 18212 14580 18214
rect 14514 18180 14580 18212
rect 14614 18212 14622 18214
rect 14656 18214 14712 18246
rect 14746 18214 14802 18246
rect 14836 18214 14892 18246
rect 14656 18212 14680 18214
rect 14746 18212 14780 18214
rect 14836 18212 14880 18214
rect 14926 18212 14987 18246
rect 14614 18180 14680 18212
rect 14714 18180 14780 18212
rect 14814 18180 14880 18212
rect 14914 18180 14987 18212
rect 14293 18156 14987 18180
rect 14293 18122 14352 18156
rect 14386 18122 14442 18156
rect 14476 18122 14532 18156
rect 14566 18122 14622 18156
rect 14656 18122 14712 18156
rect 14746 18122 14802 18156
rect 14836 18122 14892 18156
rect 14926 18122 14987 18156
rect 14293 18114 14987 18122
rect 14293 18080 14380 18114
rect 14414 18080 14480 18114
rect 14514 18080 14580 18114
rect 14614 18080 14680 18114
rect 14714 18080 14780 18114
rect 14814 18080 14880 18114
rect 14914 18080 14987 18114
rect 14293 18066 14987 18080
rect 14293 18032 14352 18066
rect 14386 18032 14442 18066
rect 14476 18032 14532 18066
rect 14566 18032 14622 18066
rect 14656 18032 14712 18066
rect 14746 18032 14802 18066
rect 14836 18032 14892 18066
rect 14926 18032 14987 18066
rect 14293 18014 14987 18032
rect 14293 17980 14380 18014
rect 14414 17980 14480 18014
rect 14514 17980 14580 18014
rect 14614 17980 14680 18014
rect 14714 17980 14780 18014
rect 14814 17980 14880 18014
rect 14914 17980 14987 18014
rect 14293 17976 14987 17980
rect 14293 17942 14352 17976
rect 14386 17942 14442 17976
rect 14476 17942 14532 17976
rect 14566 17942 14622 17976
rect 14656 17942 14712 17976
rect 14746 17942 14802 17976
rect 14836 17942 14892 17976
rect 14926 17942 14987 17976
rect 14293 17914 14987 17942
rect 14293 17886 14380 17914
rect 14414 17886 14480 17914
rect 14293 17852 14352 17886
rect 14414 17880 14442 17886
rect 14386 17852 14442 17880
rect 14476 17880 14480 17886
rect 14514 17886 14580 17914
rect 14514 17880 14532 17886
rect 14476 17852 14532 17880
rect 14566 17880 14580 17886
rect 14614 17886 14680 17914
rect 14714 17886 14780 17914
rect 14814 17886 14880 17914
rect 14914 17886 14987 17914
rect 14614 17880 14622 17886
rect 14566 17852 14622 17880
rect 14656 17880 14680 17886
rect 14746 17880 14780 17886
rect 14836 17880 14880 17886
rect 14656 17852 14712 17880
rect 14746 17852 14802 17880
rect 14836 17852 14892 17880
rect 14926 17852 14987 17886
rect 14293 17793 14987 17852
rect 15049 18455 15068 18489
rect 15102 18455 15121 18489
rect 15049 18399 15121 18455
rect 15049 18365 15068 18399
rect 15102 18365 15121 18399
rect 15049 18309 15121 18365
rect 15049 18275 15068 18309
rect 15102 18275 15121 18309
rect 15049 18219 15121 18275
rect 15049 18185 15068 18219
rect 15102 18185 15121 18219
rect 15049 18129 15121 18185
rect 15049 18095 15068 18129
rect 15102 18095 15121 18129
rect 15049 18039 15121 18095
rect 15049 18005 15068 18039
rect 15102 18005 15121 18039
rect 15049 17949 15121 18005
rect 15049 17915 15068 17949
rect 15102 17915 15121 17949
rect 15049 17859 15121 17915
rect 15049 17825 15068 17859
rect 15102 17825 15121 17859
rect 14159 17754 14178 17788
rect 14212 17754 14231 17788
rect 14159 17740 14231 17754
rect 15049 17769 15121 17825
rect 15049 17740 15068 17769
rect 14063 17735 15068 17740
rect 15102 17740 15121 17769
rect 15185 18578 15284 18634
rect 15670 18610 15750 18630
rect 15670 18597 15690 18610
rect 15730 18597 15750 18610
rect 16780 18610 16860 18630
rect 15185 18544 15216 18578
rect 15250 18544 15284 18578
rect 15185 18488 15284 18544
rect 15185 18454 15216 18488
rect 15250 18454 15284 18488
rect 15185 18398 15284 18454
rect 15185 18364 15216 18398
rect 15250 18364 15284 18398
rect 15185 18308 15284 18364
rect 15185 18274 15216 18308
rect 15250 18274 15284 18308
rect 15185 18218 15284 18274
rect 15185 18184 15216 18218
rect 15250 18184 15284 18218
rect 15185 18128 15284 18184
rect 15185 18094 15216 18128
rect 15250 18094 15284 18128
rect 15185 18038 15284 18094
rect 15185 18004 15216 18038
rect 15250 18004 15284 18038
rect 15185 17948 15284 18004
rect 15185 17914 15216 17948
rect 15250 17914 15284 17948
rect 15185 17858 15284 17914
rect 15185 17824 15216 17858
rect 15250 17824 15284 17858
rect 15185 17768 15284 17824
rect 15185 17740 15216 17768
rect 15102 17735 15216 17740
rect 14063 17734 15216 17735
rect 15250 17740 15284 17768
rect 15483 18563 15579 18597
rect 16171 18563 16267 18597
rect 16780 18595 16800 18610
rect 16840 18595 16860 18610
rect 15483 18501 15517 18563
rect 15670 18550 15750 18563
rect 15250 17734 15290 17740
rect 11270 17712 15290 17734
rect 11270 17678 11516 17712
rect 11550 17678 11606 17712
rect 11640 17678 11696 17712
rect 11730 17678 11786 17712
rect 11820 17678 11876 17712
rect 11910 17678 11966 17712
rect 12000 17678 12056 17712
rect 12090 17678 12146 17712
rect 12180 17678 12236 17712
rect 12270 17678 12876 17712
rect 12910 17678 12966 17712
rect 13000 17678 13056 17712
rect 13090 17678 13146 17712
rect 13180 17678 13236 17712
rect 13270 17678 13326 17712
rect 13360 17678 13416 17712
rect 13450 17678 13506 17712
rect 13540 17678 13596 17712
rect 13630 17678 14236 17712
rect 14270 17678 14326 17712
rect 14360 17678 14416 17712
rect 14450 17678 14506 17712
rect 14540 17678 14596 17712
rect 14630 17678 14686 17712
rect 14720 17678 14776 17712
rect 14810 17678 14866 17712
rect 14900 17678 14956 17712
rect 14990 17678 15290 17712
rect 11270 17644 11309 17678
rect 11343 17644 12496 17678
rect 12530 17644 12669 17678
rect 12703 17644 13856 17678
rect 13890 17644 14029 17678
rect 14063 17644 15216 17678
rect 15250 17644 15290 17678
rect 11270 17588 15290 17644
rect 11270 17554 11309 17588
rect 11343 17565 12496 17588
rect 11343 17554 11410 17565
rect 11270 17531 11410 17554
rect 11444 17531 11500 17565
rect 11534 17531 11590 17565
rect 11624 17531 11680 17565
rect 11714 17531 11770 17565
rect 11804 17531 11860 17565
rect 11894 17531 11950 17565
rect 11984 17531 12040 17565
rect 12074 17531 12130 17565
rect 12164 17531 12220 17565
rect 12254 17531 12310 17565
rect 12344 17531 12400 17565
rect 12434 17554 12496 17565
rect 12530 17554 12669 17588
rect 12703 17565 13856 17588
rect 12703 17554 12770 17565
rect 12434 17531 12770 17554
rect 12804 17531 12860 17565
rect 12894 17531 12950 17565
rect 12984 17531 13040 17565
rect 13074 17531 13130 17565
rect 13164 17531 13220 17565
rect 13254 17531 13310 17565
rect 13344 17531 13400 17565
rect 13434 17531 13490 17565
rect 13524 17531 13580 17565
rect 13614 17531 13670 17565
rect 13704 17531 13760 17565
rect 13794 17554 13856 17565
rect 13890 17554 14029 17588
rect 14063 17565 15216 17588
rect 14063 17554 14130 17565
rect 13794 17531 14130 17554
rect 14164 17531 14220 17565
rect 14254 17531 14310 17565
rect 14344 17531 14400 17565
rect 14434 17531 14490 17565
rect 14524 17531 14580 17565
rect 14614 17531 14670 17565
rect 14704 17531 14760 17565
rect 14794 17531 14850 17565
rect 14884 17531 14940 17565
rect 14974 17531 15030 17565
rect 15064 17531 15120 17565
rect 15154 17554 15216 17565
rect 15250 17554 15290 17588
rect 15154 17531 15290 17554
rect 11270 17490 15290 17531
rect 12560 17424 12640 17490
rect 13920 17424 14000 17490
rect 11276 17392 15284 17424
rect 11276 17358 11410 17392
rect 11444 17358 11500 17392
rect 11534 17358 11590 17392
rect 11624 17358 11680 17392
rect 11714 17358 11770 17392
rect 11804 17358 11860 17392
rect 11894 17358 11950 17392
rect 11984 17358 12040 17392
rect 12074 17358 12130 17392
rect 12164 17358 12220 17392
rect 12254 17358 12310 17392
rect 12344 17358 12400 17392
rect 12434 17358 12770 17392
rect 12804 17358 12860 17392
rect 12894 17358 12950 17392
rect 12984 17358 13040 17392
rect 13074 17358 13130 17392
rect 13164 17358 13220 17392
rect 13254 17358 13310 17392
rect 13344 17358 13400 17392
rect 13434 17358 13490 17392
rect 13524 17358 13580 17392
rect 13614 17358 13670 17392
rect 13704 17358 13760 17392
rect 13794 17358 14130 17392
rect 14164 17358 14220 17392
rect 14254 17358 14310 17392
rect 14344 17358 14400 17392
rect 14434 17358 14490 17392
rect 14524 17358 14580 17392
rect 14614 17358 14670 17392
rect 14704 17358 14760 17392
rect 14794 17358 14850 17392
rect 14884 17358 14940 17392
rect 14974 17358 15030 17392
rect 15064 17358 15120 17392
rect 15154 17358 15284 17392
rect 11276 17325 15284 17358
rect 11276 17308 11375 17325
rect 11276 17274 11309 17308
rect 11343 17274 11375 17308
rect 11276 17218 11375 17274
rect 12465 17308 12735 17325
rect 12465 17274 12496 17308
rect 12530 17274 12669 17308
rect 12703 17274 12735 17308
rect 11276 17184 11309 17218
rect 11343 17184 11375 17218
rect 11276 17128 11375 17184
rect 11276 17094 11309 17128
rect 11343 17094 11375 17128
rect 11276 17038 11375 17094
rect 11276 17004 11309 17038
rect 11343 17004 11375 17038
rect 11276 16948 11375 17004
rect 11276 16914 11309 16948
rect 11343 16914 11375 16948
rect 11276 16858 11375 16914
rect 11276 16824 11309 16858
rect 11343 16824 11375 16858
rect 11276 16768 11375 16824
rect 11276 16734 11309 16768
rect 11343 16734 11375 16768
rect 11276 16678 11375 16734
rect 11276 16644 11309 16678
rect 11343 16644 11375 16678
rect 11276 16588 11375 16644
rect 11276 16554 11309 16588
rect 11343 16554 11375 16588
rect 11276 16498 11375 16554
rect 11276 16464 11309 16498
rect 11343 16464 11375 16498
rect 11276 16408 11375 16464
rect 11276 16380 11309 16408
rect 10913 16181 10947 16243
rect 10163 16147 10259 16181
rect 10851 16147 10947 16181
rect 11270 16374 11309 16380
rect 11343 16380 11375 16408
rect 11439 17242 12401 17261
rect 11439 17208 11550 17242
rect 11584 17208 11640 17242
rect 11674 17208 11730 17242
rect 11764 17208 11820 17242
rect 11854 17208 11910 17242
rect 11944 17208 12000 17242
rect 12034 17208 12090 17242
rect 12124 17208 12180 17242
rect 12214 17208 12270 17242
rect 12304 17208 12401 17242
rect 11439 17189 12401 17208
rect 11439 17148 11511 17189
rect 11439 17114 11458 17148
rect 11492 17114 11511 17148
rect 12329 17129 12401 17189
rect 11439 17058 11511 17114
rect 11439 17024 11458 17058
rect 11492 17024 11511 17058
rect 11439 16968 11511 17024
rect 11439 16934 11458 16968
rect 11492 16934 11511 16968
rect 11439 16878 11511 16934
rect 11439 16844 11458 16878
rect 11492 16844 11511 16878
rect 11439 16788 11511 16844
rect 11439 16754 11458 16788
rect 11492 16754 11511 16788
rect 11439 16698 11511 16754
rect 11439 16664 11458 16698
rect 11492 16664 11511 16698
rect 11439 16608 11511 16664
rect 11439 16574 11458 16608
rect 11492 16574 11511 16608
rect 11439 16518 11511 16574
rect 11439 16484 11458 16518
rect 11492 16484 11511 16518
rect 11439 16428 11511 16484
rect 11573 17066 12267 17127
rect 11573 17032 11632 17066
rect 11666 17054 11722 17066
rect 11694 17032 11722 17054
rect 11756 17054 11812 17066
rect 11756 17032 11760 17054
rect 11573 17020 11660 17032
rect 11694 17020 11760 17032
rect 11794 17032 11812 17054
rect 11846 17054 11902 17066
rect 11846 17032 11860 17054
rect 11794 17020 11860 17032
rect 11894 17032 11902 17054
rect 11936 17054 11992 17066
rect 12026 17054 12082 17066
rect 12116 17054 12172 17066
rect 11936 17032 11960 17054
rect 12026 17032 12060 17054
rect 12116 17032 12160 17054
rect 12206 17032 12267 17066
rect 11894 17020 11960 17032
rect 11994 17020 12060 17032
rect 12094 17020 12160 17032
rect 12194 17020 12267 17032
rect 11573 16976 12267 17020
rect 11573 16942 11632 16976
rect 11666 16954 11722 16976
rect 11694 16942 11722 16954
rect 11756 16954 11812 16976
rect 11756 16942 11760 16954
rect 11573 16920 11660 16942
rect 11694 16920 11760 16942
rect 11794 16942 11812 16954
rect 11846 16954 11902 16976
rect 11846 16942 11860 16954
rect 11794 16920 11860 16942
rect 11894 16942 11902 16954
rect 11936 16954 11992 16976
rect 12026 16954 12082 16976
rect 12116 16954 12172 16976
rect 11936 16942 11960 16954
rect 12026 16942 12060 16954
rect 12116 16942 12160 16954
rect 12206 16942 12267 16976
rect 11894 16920 11960 16942
rect 11994 16920 12060 16942
rect 12094 16920 12160 16942
rect 12194 16920 12267 16942
rect 11573 16886 12267 16920
rect 11573 16852 11632 16886
rect 11666 16854 11722 16886
rect 11694 16852 11722 16854
rect 11756 16854 11812 16886
rect 11756 16852 11760 16854
rect 11573 16820 11660 16852
rect 11694 16820 11760 16852
rect 11794 16852 11812 16854
rect 11846 16854 11902 16886
rect 11846 16852 11860 16854
rect 11794 16820 11860 16852
rect 11894 16852 11902 16854
rect 11936 16854 11992 16886
rect 12026 16854 12082 16886
rect 12116 16854 12172 16886
rect 11936 16852 11960 16854
rect 12026 16852 12060 16854
rect 12116 16852 12160 16854
rect 12206 16852 12267 16886
rect 11894 16820 11960 16852
rect 11994 16820 12060 16852
rect 12094 16820 12160 16852
rect 12194 16820 12267 16852
rect 11573 16796 12267 16820
rect 11573 16762 11632 16796
rect 11666 16762 11722 16796
rect 11756 16762 11812 16796
rect 11846 16762 11902 16796
rect 11936 16762 11992 16796
rect 12026 16762 12082 16796
rect 12116 16762 12172 16796
rect 12206 16762 12267 16796
rect 11573 16754 12267 16762
rect 11573 16720 11660 16754
rect 11694 16720 11760 16754
rect 11794 16720 11860 16754
rect 11894 16720 11960 16754
rect 11994 16720 12060 16754
rect 12094 16720 12160 16754
rect 12194 16720 12267 16754
rect 11573 16706 12267 16720
rect 11573 16672 11632 16706
rect 11666 16672 11722 16706
rect 11756 16672 11812 16706
rect 11846 16672 11902 16706
rect 11936 16672 11992 16706
rect 12026 16672 12082 16706
rect 12116 16672 12172 16706
rect 12206 16672 12267 16706
rect 11573 16654 12267 16672
rect 11573 16620 11660 16654
rect 11694 16620 11760 16654
rect 11794 16620 11860 16654
rect 11894 16620 11960 16654
rect 11994 16620 12060 16654
rect 12094 16620 12160 16654
rect 12194 16620 12267 16654
rect 11573 16616 12267 16620
rect 11573 16582 11632 16616
rect 11666 16582 11722 16616
rect 11756 16582 11812 16616
rect 11846 16582 11902 16616
rect 11936 16582 11992 16616
rect 12026 16582 12082 16616
rect 12116 16582 12172 16616
rect 12206 16582 12267 16616
rect 11573 16554 12267 16582
rect 11573 16526 11660 16554
rect 11694 16526 11760 16554
rect 11573 16492 11632 16526
rect 11694 16520 11722 16526
rect 11666 16492 11722 16520
rect 11756 16520 11760 16526
rect 11794 16526 11860 16554
rect 11794 16520 11812 16526
rect 11756 16492 11812 16520
rect 11846 16520 11860 16526
rect 11894 16526 11960 16554
rect 11994 16526 12060 16554
rect 12094 16526 12160 16554
rect 12194 16526 12267 16554
rect 11894 16520 11902 16526
rect 11846 16492 11902 16520
rect 11936 16520 11960 16526
rect 12026 16520 12060 16526
rect 12116 16520 12160 16526
rect 11936 16492 11992 16520
rect 12026 16492 12082 16520
rect 12116 16492 12172 16520
rect 12206 16492 12267 16526
rect 11573 16433 12267 16492
rect 12329 17095 12348 17129
rect 12382 17095 12401 17129
rect 12329 17039 12401 17095
rect 12329 17005 12348 17039
rect 12382 17005 12401 17039
rect 12329 16949 12401 17005
rect 12329 16915 12348 16949
rect 12382 16915 12401 16949
rect 12329 16859 12401 16915
rect 12329 16825 12348 16859
rect 12382 16825 12401 16859
rect 12329 16769 12401 16825
rect 12329 16735 12348 16769
rect 12382 16735 12401 16769
rect 12329 16679 12401 16735
rect 12329 16645 12348 16679
rect 12382 16645 12401 16679
rect 12329 16589 12401 16645
rect 12329 16555 12348 16589
rect 12382 16555 12401 16589
rect 12329 16499 12401 16555
rect 12329 16465 12348 16499
rect 12382 16465 12401 16499
rect 11439 16394 11458 16428
rect 11492 16394 11511 16428
rect 11439 16380 11511 16394
rect 12329 16409 12401 16465
rect 12329 16380 12348 16409
rect 11343 16375 12348 16380
rect 12382 16380 12401 16409
rect 12465 17218 12735 17274
rect 13825 17308 14095 17325
rect 13825 17274 13856 17308
rect 13890 17274 14029 17308
rect 14063 17274 14095 17308
rect 12465 17184 12496 17218
rect 12530 17184 12669 17218
rect 12703 17184 12735 17218
rect 12465 17128 12735 17184
rect 12465 17094 12496 17128
rect 12530 17094 12669 17128
rect 12703 17094 12735 17128
rect 12465 17038 12735 17094
rect 12465 17004 12496 17038
rect 12530 17004 12669 17038
rect 12703 17004 12735 17038
rect 12465 16948 12735 17004
rect 12465 16914 12496 16948
rect 12530 16914 12669 16948
rect 12703 16914 12735 16948
rect 12465 16858 12735 16914
rect 12465 16824 12496 16858
rect 12530 16824 12669 16858
rect 12703 16824 12735 16858
rect 12465 16768 12735 16824
rect 12465 16734 12496 16768
rect 12530 16734 12669 16768
rect 12703 16734 12735 16768
rect 12465 16678 12735 16734
rect 12465 16644 12496 16678
rect 12530 16644 12669 16678
rect 12703 16644 12735 16678
rect 12465 16588 12735 16644
rect 12465 16554 12496 16588
rect 12530 16554 12669 16588
rect 12703 16554 12735 16588
rect 12465 16498 12735 16554
rect 12465 16464 12496 16498
rect 12530 16464 12669 16498
rect 12703 16464 12735 16498
rect 12465 16408 12735 16464
rect 12465 16380 12496 16408
rect 12382 16375 12496 16380
rect 11343 16374 12496 16375
rect 12530 16374 12669 16408
rect 12703 16380 12735 16408
rect 12799 17242 13761 17261
rect 12799 17208 12910 17242
rect 12944 17208 13000 17242
rect 13034 17208 13090 17242
rect 13124 17208 13180 17242
rect 13214 17208 13270 17242
rect 13304 17208 13360 17242
rect 13394 17208 13450 17242
rect 13484 17208 13540 17242
rect 13574 17208 13630 17242
rect 13664 17208 13761 17242
rect 12799 17189 13761 17208
rect 12799 17148 12871 17189
rect 12799 17114 12818 17148
rect 12852 17114 12871 17148
rect 13689 17129 13761 17189
rect 12799 17058 12871 17114
rect 12799 17024 12818 17058
rect 12852 17024 12871 17058
rect 12799 16968 12871 17024
rect 12799 16934 12818 16968
rect 12852 16934 12871 16968
rect 12799 16878 12871 16934
rect 12799 16844 12818 16878
rect 12852 16844 12871 16878
rect 12799 16788 12871 16844
rect 12799 16754 12818 16788
rect 12852 16754 12871 16788
rect 12799 16698 12871 16754
rect 12799 16664 12818 16698
rect 12852 16664 12871 16698
rect 12799 16608 12871 16664
rect 12799 16574 12818 16608
rect 12852 16574 12871 16608
rect 12799 16518 12871 16574
rect 12799 16484 12818 16518
rect 12852 16484 12871 16518
rect 12799 16428 12871 16484
rect 12933 17066 13627 17127
rect 12933 17032 12992 17066
rect 13026 17054 13082 17066
rect 13054 17032 13082 17054
rect 13116 17054 13172 17066
rect 13116 17032 13120 17054
rect 12933 17020 13020 17032
rect 13054 17020 13120 17032
rect 13154 17032 13172 17054
rect 13206 17054 13262 17066
rect 13206 17032 13220 17054
rect 13154 17020 13220 17032
rect 13254 17032 13262 17054
rect 13296 17054 13352 17066
rect 13386 17054 13442 17066
rect 13476 17054 13532 17066
rect 13296 17032 13320 17054
rect 13386 17032 13420 17054
rect 13476 17032 13520 17054
rect 13566 17032 13627 17066
rect 13254 17020 13320 17032
rect 13354 17020 13420 17032
rect 13454 17020 13520 17032
rect 13554 17020 13627 17032
rect 12933 16976 13627 17020
rect 12933 16942 12992 16976
rect 13026 16954 13082 16976
rect 13054 16942 13082 16954
rect 13116 16954 13172 16976
rect 13116 16942 13120 16954
rect 12933 16920 13020 16942
rect 13054 16920 13120 16942
rect 13154 16942 13172 16954
rect 13206 16954 13262 16976
rect 13206 16942 13220 16954
rect 13154 16920 13220 16942
rect 13254 16942 13262 16954
rect 13296 16954 13352 16976
rect 13386 16954 13442 16976
rect 13476 16954 13532 16976
rect 13296 16942 13320 16954
rect 13386 16942 13420 16954
rect 13476 16942 13520 16954
rect 13566 16942 13627 16976
rect 13254 16920 13320 16942
rect 13354 16920 13420 16942
rect 13454 16920 13520 16942
rect 13554 16920 13627 16942
rect 12933 16886 13627 16920
rect 12933 16852 12992 16886
rect 13026 16854 13082 16886
rect 13054 16852 13082 16854
rect 13116 16854 13172 16886
rect 13116 16852 13120 16854
rect 12933 16820 13020 16852
rect 13054 16820 13120 16852
rect 13154 16852 13172 16854
rect 13206 16854 13262 16886
rect 13206 16852 13220 16854
rect 13154 16820 13220 16852
rect 13254 16852 13262 16854
rect 13296 16854 13352 16886
rect 13386 16854 13442 16886
rect 13476 16854 13532 16886
rect 13296 16852 13320 16854
rect 13386 16852 13420 16854
rect 13476 16852 13520 16854
rect 13566 16852 13627 16886
rect 13254 16820 13320 16852
rect 13354 16820 13420 16852
rect 13454 16820 13520 16852
rect 13554 16820 13627 16852
rect 12933 16796 13627 16820
rect 12933 16762 12992 16796
rect 13026 16762 13082 16796
rect 13116 16762 13172 16796
rect 13206 16762 13262 16796
rect 13296 16762 13352 16796
rect 13386 16762 13442 16796
rect 13476 16762 13532 16796
rect 13566 16762 13627 16796
rect 12933 16754 13627 16762
rect 12933 16720 13020 16754
rect 13054 16720 13120 16754
rect 13154 16720 13220 16754
rect 13254 16720 13320 16754
rect 13354 16720 13420 16754
rect 13454 16720 13520 16754
rect 13554 16720 13627 16754
rect 12933 16706 13627 16720
rect 12933 16672 12992 16706
rect 13026 16672 13082 16706
rect 13116 16672 13172 16706
rect 13206 16672 13262 16706
rect 13296 16672 13352 16706
rect 13386 16672 13442 16706
rect 13476 16672 13532 16706
rect 13566 16672 13627 16706
rect 12933 16654 13627 16672
rect 12933 16620 13020 16654
rect 13054 16620 13120 16654
rect 13154 16620 13220 16654
rect 13254 16620 13320 16654
rect 13354 16620 13420 16654
rect 13454 16620 13520 16654
rect 13554 16620 13627 16654
rect 12933 16616 13627 16620
rect 12933 16582 12992 16616
rect 13026 16582 13082 16616
rect 13116 16582 13172 16616
rect 13206 16582 13262 16616
rect 13296 16582 13352 16616
rect 13386 16582 13442 16616
rect 13476 16582 13532 16616
rect 13566 16582 13627 16616
rect 12933 16554 13627 16582
rect 12933 16526 13020 16554
rect 13054 16526 13120 16554
rect 12933 16492 12992 16526
rect 13054 16520 13082 16526
rect 13026 16492 13082 16520
rect 13116 16520 13120 16526
rect 13154 16526 13220 16554
rect 13154 16520 13172 16526
rect 13116 16492 13172 16520
rect 13206 16520 13220 16526
rect 13254 16526 13320 16554
rect 13354 16526 13420 16554
rect 13454 16526 13520 16554
rect 13554 16526 13627 16554
rect 13254 16520 13262 16526
rect 13206 16492 13262 16520
rect 13296 16520 13320 16526
rect 13386 16520 13420 16526
rect 13476 16520 13520 16526
rect 13296 16492 13352 16520
rect 13386 16492 13442 16520
rect 13476 16492 13532 16520
rect 13566 16492 13627 16526
rect 12933 16433 13627 16492
rect 13689 17095 13708 17129
rect 13742 17095 13761 17129
rect 13689 17039 13761 17095
rect 13689 17005 13708 17039
rect 13742 17005 13761 17039
rect 13689 16949 13761 17005
rect 13689 16915 13708 16949
rect 13742 16915 13761 16949
rect 13689 16859 13761 16915
rect 13689 16825 13708 16859
rect 13742 16825 13761 16859
rect 13689 16769 13761 16825
rect 13689 16735 13708 16769
rect 13742 16735 13761 16769
rect 13689 16679 13761 16735
rect 13689 16645 13708 16679
rect 13742 16645 13761 16679
rect 13689 16589 13761 16645
rect 13689 16555 13708 16589
rect 13742 16555 13761 16589
rect 13689 16499 13761 16555
rect 13689 16465 13708 16499
rect 13742 16465 13761 16499
rect 12799 16394 12818 16428
rect 12852 16394 12871 16428
rect 12799 16380 12871 16394
rect 13689 16409 13761 16465
rect 13689 16380 13708 16409
rect 12703 16375 13708 16380
rect 13742 16380 13761 16409
rect 13825 17218 14095 17274
rect 15185 17308 15284 17325
rect 15185 17274 15216 17308
rect 15250 17274 15284 17308
rect 13825 17184 13856 17218
rect 13890 17184 14029 17218
rect 14063 17184 14095 17218
rect 13825 17128 14095 17184
rect 13825 17094 13856 17128
rect 13890 17094 14029 17128
rect 14063 17094 14095 17128
rect 13825 17038 14095 17094
rect 13825 17004 13856 17038
rect 13890 17004 14029 17038
rect 14063 17004 14095 17038
rect 13825 16948 14095 17004
rect 13825 16914 13856 16948
rect 13890 16914 14029 16948
rect 14063 16914 14095 16948
rect 13825 16858 14095 16914
rect 13825 16824 13856 16858
rect 13890 16824 14029 16858
rect 14063 16824 14095 16858
rect 13825 16768 14095 16824
rect 13825 16734 13856 16768
rect 13890 16734 14029 16768
rect 14063 16734 14095 16768
rect 13825 16678 14095 16734
rect 13825 16644 13856 16678
rect 13890 16644 14029 16678
rect 14063 16644 14095 16678
rect 13825 16588 14095 16644
rect 13825 16554 13856 16588
rect 13890 16554 14029 16588
rect 14063 16554 14095 16588
rect 13825 16498 14095 16554
rect 13825 16464 13856 16498
rect 13890 16464 14029 16498
rect 14063 16464 14095 16498
rect 13825 16408 14095 16464
rect 13825 16380 13856 16408
rect 13742 16375 13856 16380
rect 12703 16374 13856 16375
rect 13890 16374 14029 16408
rect 14063 16380 14095 16408
rect 14159 17242 15121 17261
rect 14159 17208 14270 17242
rect 14304 17208 14360 17242
rect 14394 17208 14450 17242
rect 14484 17208 14540 17242
rect 14574 17208 14630 17242
rect 14664 17208 14720 17242
rect 14754 17208 14810 17242
rect 14844 17208 14900 17242
rect 14934 17208 14990 17242
rect 15024 17208 15121 17242
rect 14159 17189 15121 17208
rect 14159 17148 14231 17189
rect 14159 17114 14178 17148
rect 14212 17114 14231 17148
rect 15049 17129 15121 17189
rect 14159 17058 14231 17114
rect 14159 17024 14178 17058
rect 14212 17024 14231 17058
rect 14159 16968 14231 17024
rect 14159 16934 14178 16968
rect 14212 16934 14231 16968
rect 14159 16878 14231 16934
rect 14159 16844 14178 16878
rect 14212 16844 14231 16878
rect 14159 16788 14231 16844
rect 14159 16754 14178 16788
rect 14212 16754 14231 16788
rect 14159 16698 14231 16754
rect 14159 16664 14178 16698
rect 14212 16664 14231 16698
rect 14159 16608 14231 16664
rect 14159 16574 14178 16608
rect 14212 16574 14231 16608
rect 14159 16518 14231 16574
rect 14159 16484 14178 16518
rect 14212 16484 14231 16518
rect 14159 16428 14231 16484
rect 14293 17066 14987 17127
rect 14293 17032 14352 17066
rect 14386 17054 14442 17066
rect 14414 17032 14442 17054
rect 14476 17054 14532 17066
rect 14476 17032 14480 17054
rect 14293 17020 14380 17032
rect 14414 17020 14480 17032
rect 14514 17032 14532 17054
rect 14566 17054 14622 17066
rect 14566 17032 14580 17054
rect 14514 17020 14580 17032
rect 14614 17032 14622 17054
rect 14656 17054 14712 17066
rect 14746 17054 14802 17066
rect 14836 17054 14892 17066
rect 14656 17032 14680 17054
rect 14746 17032 14780 17054
rect 14836 17032 14880 17054
rect 14926 17032 14987 17066
rect 14614 17020 14680 17032
rect 14714 17020 14780 17032
rect 14814 17020 14880 17032
rect 14914 17020 14987 17032
rect 14293 16976 14987 17020
rect 14293 16942 14352 16976
rect 14386 16954 14442 16976
rect 14414 16942 14442 16954
rect 14476 16954 14532 16976
rect 14476 16942 14480 16954
rect 14293 16920 14380 16942
rect 14414 16920 14480 16942
rect 14514 16942 14532 16954
rect 14566 16954 14622 16976
rect 14566 16942 14580 16954
rect 14514 16920 14580 16942
rect 14614 16942 14622 16954
rect 14656 16954 14712 16976
rect 14746 16954 14802 16976
rect 14836 16954 14892 16976
rect 14656 16942 14680 16954
rect 14746 16942 14780 16954
rect 14836 16942 14880 16954
rect 14926 16942 14987 16976
rect 14614 16920 14680 16942
rect 14714 16920 14780 16942
rect 14814 16920 14880 16942
rect 14914 16920 14987 16942
rect 14293 16886 14987 16920
rect 14293 16852 14352 16886
rect 14386 16854 14442 16886
rect 14414 16852 14442 16854
rect 14476 16854 14532 16886
rect 14476 16852 14480 16854
rect 14293 16820 14380 16852
rect 14414 16820 14480 16852
rect 14514 16852 14532 16854
rect 14566 16854 14622 16886
rect 14566 16852 14580 16854
rect 14514 16820 14580 16852
rect 14614 16852 14622 16854
rect 14656 16854 14712 16886
rect 14746 16854 14802 16886
rect 14836 16854 14892 16886
rect 14656 16852 14680 16854
rect 14746 16852 14780 16854
rect 14836 16852 14880 16854
rect 14926 16852 14987 16886
rect 14614 16820 14680 16852
rect 14714 16820 14780 16852
rect 14814 16820 14880 16852
rect 14914 16820 14987 16852
rect 14293 16796 14987 16820
rect 14293 16762 14352 16796
rect 14386 16762 14442 16796
rect 14476 16762 14532 16796
rect 14566 16762 14622 16796
rect 14656 16762 14712 16796
rect 14746 16762 14802 16796
rect 14836 16762 14892 16796
rect 14926 16762 14987 16796
rect 14293 16754 14987 16762
rect 14293 16720 14380 16754
rect 14414 16720 14480 16754
rect 14514 16720 14580 16754
rect 14614 16720 14680 16754
rect 14714 16720 14780 16754
rect 14814 16720 14880 16754
rect 14914 16720 14987 16754
rect 14293 16706 14987 16720
rect 14293 16672 14352 16706
rect 14386 16672 14442 16706
rect 14476 16672 14532 16706
rect 14566 16672 14622 16706
rect 14656 16672 14712 16706
rect 14746 16672 14802 16706
rect 14836 16672 14892 16706
rect 14926 16672 14987 16706
rect 14293 16654 14987 16672
rect 14293 16620 14380 16654
rect 14414 16620 14480 16654
rect 14514 16620 14580 16654
rect 14614 16620 14680 16654
rect 14714 16620 14780 16654
rect 14814 16620 14880 16654
rect 14914 16620 14987 16654
rect 14293 16616 14987 16620
rect 14293 16582 14352 16616
rect 14386 16582 14442 16616
rect 14476 16582 14532 16616
rect 14566 16582 14622 16616
rect 14656 16582 14712 16616
rect 14746 16582 14802 16616
rect 14836 16582 14892 16616
rect 14926 16582 14987 16616
rect 14293 16554 14987 16582
rect 14293 16526 14380 16554
rect 14414 16526 14480 16554
rect 14293 16492 14352 16526
rect 14414 16520 14442 16526
rect 14386 16492 14442 16520
rect 14476 16520 14480 16526
rect 14514 16526 14580 16554
rect 14514 16520 14532 16526
rect 14476 16492 14532 16520
rect 14566 16520 14580 16526
rect 14614 16526 14680 16554
rect 14714 16526 14780 16554
rect 14814 16526 14880 16554
rect 14914 16526 14987 16554
rect 14614 16520 14622 16526
rect 14566 16492 14622 16520
rect 14656 16520 14680 16526
rect 14746 16520 14780 16526
rect 14836 16520 14880 16526
rect 14656 16492 14712 16520
rect 14746 16492 14802 16520
rect 14836 16492 14892 16520
rect 14926 16492 14987 16526
rect 14293 16433 14987 16492
rect 15049 17095 15068 17129
rect 15102 17095 15121 17129
rect 15049 17039 15121 17095
rect 15049 17005 15068 17039
rect 15102 17005 15121 17039
rect 15049 16949 15121 17005
rect 15049 16915 15068 16949
rect 15102 16915 15121 16949
rect 15049 16859 15121 16915
rect 15049 16825 15068 16859
rect 15102 16825 15121 16859
rect 15049 16769 15121 16825
rect 15049 16735 15068 16769
rect 15102 16735 15121 16769
rect 15049 16679 15121 16735
rect 15049 16645 15068 16679
rect 15102 16645 15121 16679
rect 15049 16589 15121 16645
rect 15049 16555 15068 16589
rect 15102 16555 15121 16589
rect 15049 16499 15121 16555
rect 15049 16465 15068 16499
rect 15102 16465 15121 16499
rect 14159 16394 14178 16428
rect 14212 16394 14231 16428
rect 14159 16380 14231 16394
rect 15049 16409 15121 16465
rect 15049 16380 15068 16409
rect 14063 16375 15068 16380
rect 15102 16380 15121 16409
rect 15185 17218 15284 17274
rect 15185 17184 15216 17218
rect 15250 17184 15284 17218
rect 15185 17128 15284 17184
rect 15185 17094 15216 17128
rect 15250 17094 15284 17128
rect 15185 17038 15284 17094
rect 15185 17004 15216 17038
rect 15250 17004 15284 17038
rect 15185 16948 15284 17004
rect 15185 16914 15216 16948
rect 15250 16914 15284 16948
rect 15185 16858 15284 16914
rect 15185 16824 15216 16858
rect 15250 16824 15284 16858
rect 15185 16768 15284 16824
rect 15185 16734 15216 16768
rect 15250 16734 15284 16768
rect 15185 16678 15284 16734
rect 15185 16644 15216 16678
rect 15250 16644 15284 16678
rect 15185 16588 15284 16644
rect 15185 16554 15216 16588
rect 15250 16554 15284 16588
rect 15185 16498 15284 16554
rect 15185 16464 15216 16498
rect 15250 16464 15284 16498
rect 15185 16408 15284 16464
rect 15185 16380 15216 16408
rect 15102 16375 15216 16380
rect 14063 16374 15216 16375
rect 15250 16380 15284 16408
rect 15250 16374 15290 16380
rect 11270 16352 15290 16374
rect 11270 16318 11516 16352
rect 11550 16318 11606 16352
rect 11640 16318 11696 16352
rect 11730 16318 11786 16352
rect 11820 16318 11876 16352
rect 11910 16318 11966 16352
rect 12000 16318 12056 16352
rect 12090 16318 12146 16352
rect 12180 16318 12236 16352
rect 12270 16318 12876 16352
rect 12910 16318 12966 16352
rect 13000 16318 13056 16352
rect 13090 16318 13146 16352
rect 13180 16318 13236 16352
rect 13270 16318 13326 16352
rect 13360 16318 13416 16352
rect 13450 16318 13506 16352
rect 13540 16318 13596 16352
rect 13630 16318 14236 16352
rect 14270 16318 14326 16352
rect 14360 16318 14416 16352
rect 14450 16318 14506 16352
rect 14540 16318 14596 16352
rect 14630 16318 14686 16352
rect 14720 16318 14776 16352
rect 14810 16318 14866 16352
rect 14900 16318 14956 16352
rect 14990 16318 15290 16352
rect 11270 16284 11309 16318
rect 11343 16284 12496 16318
rect 12530 16284 12669 16318
rect 12703 16284 13856 16318
rect 13890 16284 14029 16318
rect 14063 16284 15216 16318
rect 15250 16284 15290 16318
rect 11270 16228 15290 16284
rect 11270 16194 11309 16228
rect 11343 16205 12496 16228
rect 11343 16194 11410 16205
rect 11270 16171 11410 16194
rect 11444 16171 11500 16205
rect 11534 16171 11590 16205
rect 11624 16171 11680 16205
rect 11714 16171 11770 16205
rect 11804 16171 11860 16205
rect 11894 16171 11950 16205
rect 11984 16171 12040 16205
rect 12074 16171 12130 16205
rect 12164 16171 12220 16205
rect 12254 16171 12310 16205
rect 12344 16171 12400 16205
rect 12434 16194 12496 16205
rect 12530 16194 12669 16228
rect 12703 16205 13856 16228
rect 12703 16194 12770 16205
rect 12434 16171 12770 16194
rect 12804 16171 12860 16205
rect 12894 16171 12950 16205
rect 12984 16171 13040 16205
rect 13074 16171 13130 16205
rect 13164 16171 13220 16205
rect 13254 16171 13310 16205
rect 13344 16171 13400 16205
rect 13434 16171 13490 16205
rect 13524 16171 13580 16205
rect 13614 16171 13670 16205
rect 13704 16171 13760 16205
rect 13794 16194 13856 16205
rect 13890 16194 14029 16228
rect 14063 16205 15216 16228
rect 14063 16194 14130 16205
rect 13794 16171 14130 16194
rect 14164 16171 14220 16205
rect 14254 16171 14310 16205
rect 14344 16171 14400 16205
rect 14434 16171 14490 16205
rect 14524 16171 14580 16205
rect 14614 16171 14670 16205
rect 14704 16171 14760 16205
rect 14794 16171 14850 16205
rect 14884 16171 14940 16205
rect 14974 16171 15030 16205
rect 15064 16171 15120 16205
rect 15154 16194 15216 16205
rect 15250 16194 15290 16228
rect 15154 16171 15290 16194
rect 11270 16130 15290 16171
rect 16233 18501 16267 18563
rect 15483 16181 15517 16243
rect 16233 16181 16267 16243
rect 15483 16147 15579 16181
rect 16171 16147 16267 16181
rect 16593 18561 16689 18595
rect 16949 18561 17045 18595
rect 17570 18590 17650 18610
rect 17570 18589 17590 18590
rect 17630 18589 17650 18590
rect 16593 18499 16627 18561
rect 16780 18550 16860 18561
rect 12560 16064 12640 16130
rect 13920 16064 14000 16130
rect 11276 16032 15284 16064
rect 11276 15998 11410 16032
rect 11444 15998 11500 16032
rect 11534 15998 11590 16032
rect 11624 15998 11680 16032
rect 11714 15998 11770 16032
rect 11804 15998 11860 16032
rect 11894 15998 11950 16032
rect 11984 15998 12040 16032
rect 12074 15998 12130 16032
rect 12164 15998 12220 16032
rect 12254 15998 12310 16032
rect 12344 15998 12400 16032
rect 12434 15998 12770 16032
rect 12804 15998 12860 16032
rect 12894 15998 12950 16032
rect 12984 15998 13040 16032
rect 13074 15998 13130 16032
rect 13164 15998 13220 16032
rect 13254 15998 13310 16032
rect 13344 15998 13400 16032
rect 13434 15998 13490 16032
rect 13524 15998 13580 16032
rect 13614 15998 13670 16032
rect 13704 15998 13760 16032
rect 13794 15998 14130 16032
rect 14164 15998 14220 16032
rect 14254 15998 14310 16032
rect 14344 15998 14400 16032
rect 14434 15998 14490 16032
rect 14524 15998 14580 16032
rect 14614 15998 14670 16032
rect 14704 15998 14760 16032
rect 14794 15998 14850 16032
rect 14884 15998 14940 16032
rect 14974 15998 15030 16032
rect 15064 15998 15120 16032
rect 15154 15998 15284 16032
rect 11276 15965 15284 15998
rect 11276 15948 11375 15965
rect 11276 15914 11309 15948
rect 11343 15914 11375 15948
rect 11276 15858 11375 15914
rect 12465 15948 12735 15965
rect 12465 15914 12496 15948
rect 12530 15914 12669 15948
rect 12703 15914 12735 15948
rect 11276 15824 11309 15858
rect 11343 15824 11375 15858
rect 11276 15768 11375 15824
rect 11276 15734 11309 15768
rect 11343 15734 11375 15768
rect 11276 15678 11375 15734
rect 11276 15644 11309 15678
rect 11343 15644 11375 15678
rect 11276 15588 11375 15644
rect 11276 15554 11309 15588
rect 11343 15554 11375 15588
rect 11276 15498 11375 15554
rect 11276 15464 11309 15498
rect 11343 15464 11375 15498
rect 11276 15408 11375 15464
rect 11276 15374 11309 15408
rect 11343 15374 11375 15408
rect 11276 15318 11375 15374
rect 11276 15284 11309 15318
rect 11343 15284 11375 15318
rect 11276 15228 11375 15284
rect 11276 15194 11309 15228
rect 11343 15194 11375 15228
rect 11276 15138 11375 15194
rect 11276 15104 11309 15138
rect 11343 15104 11375 15138
rect 11276 15048 11375 15104
rect 11276 15020 11309 15048
rect 9801 14957 9835 15019
rect 9383 14923 9479 14957
rect 9739 14923 9835 14957
rect 11270 15014 11309 15020
rect 11343 15020 11375 15048
rect 11439 15882 12401 15901
rect 11439 15848 11550 15882
rect 11584 15848 11640 15882
rect 11674 15848 11730 15882
rect 11764 15848 11820 15882
rect 11854 15848 11910 15882
rect 11944 15848 12000 15882
rect 12034 15848 12090 15882
rect 12124 15848 12180 15882
rect 12214 15848 12270 15882
rect 12304 15848 12401 15882
rect 11439 15829 12401 15848
rect 11439 15788 11511 15829
rect 11439 15754 11458 15788
rect 11492 15754 11511 15788
rect 12329 15769 12401 15829
rect 11439 15698 11511 15754
rect 11439 15664 11458 15698
rect 11492 15664 11511 15698
rect 11439 15608 11511 15664
rect 11439 15574 11458 15608
rect 11492 15574 11511 15608
rect 11439 15518 11511 15574
rect 11439 15484 11458 15518
rect 11492 15484 11511 15518
rect 11439 15428 11511 15484
rect 11439 15394 11458 15428
rect 11492 15394 11511 15428
rect 11439 15338 11511 15394
rect 11439 15304 11458 15338
rect 11492 15304 11511 15338
rect 11439 15248 11511 15304
rect 11439 15214 11458 15248
rect 11492 15214 11511 15248
rect 11439 15158 11511 15214
rect 11439 15124 11458 15158
rect 11492 15124 11511 15158
rect 11439 15068 11511 15124
rect 11573 15706 12267 15767
rect 11573 15672 11632 15706
rect 11666 15694 11722 15706
rect 11694 15672 11722 15694
rect 11756 15694 11812 15706
rect 11756 15672 11760 15694
rect 11573 15660 11660 15672
rect 11694 15660 11760 15672
rect 11794 15672 11812 15694
rect 11846 15694 11902 15706
rect 11846 15672 11860 15694
rect 11794 15660 11860 15672
rect 11894 15672 11902 15694
rect 11936 15694 11992 15706
rect 12026 15694 12082 15706
rect 12116 15694 12172 15706
rect 11936 15672 11960 15694
rect 12026 15672 12060 15694
rect 12116 15672 12160 15694
rect 12206 15672 12267 15706
rect 11894 15660 11960 15672
rect 11994 15660 12060 15672
rect 12094 15660 12160 15672
rect 12194 15660 12267 15672
rect 11573 15616 12267 15660
rect 11573 15582 11632 15616
rect 11666 15594 11722 15616
rect 11694 15582 11722 15594
rect 11756 15594 11812 15616
rect 11756 15582 11760 15594
rect 11573 15560 11660 15582
rect 11694 15560 11760 15582
rect 11794 15582 11812 15594
rect 11846 15594 11902 15616
rect 11846 15582 11860 15594
rect 11794 15560 11860 15582
rect 11894 15582 11902 15594
rect 11936 15594 11992 15616
rect 12026 15594 12082 15616
rect 12116 15594 12172 15616
rect 11936 15582 11960 15594
rect 12026 15582 12060 15594
rect 12116 15582 12160 15594
rect 12206 15582 12267 15616
rect 11894 15560 11960 15582
rect 11994 15560 12060 15582
rect 12094 15560 12160 15582
rect 12194 15560 12267 15582
rect 11573 15526 12267 15560
rect 11573 15492 11632 15526
rect 11666 15494 11722 15526
rect 11694 15492 11722 15494
rect 11756 15494 11812 15526
rect 11756 15492 11760 15494
rect 11573 15460 11660 15492
rect 11694 15460 11760 15492
rect 11794 15492 11812 15494
rect 11846 15494 11902 15526
rect 11846 15492 11860 15494
rect 11794 15460 11860 15492
rect 11894 15492 11902 15494
rect 11936 15494 11992 15526
rect 12026 15494 12082 15526
rect 12116 15494 12172 15526
rect 11936 15492 11960 15494
rect 12026 15492 12060 15494
rect 12116 15492 12160 15494
rect 12206 15492 12267 15526
rect 11894 15460 11960 15492
rect 11994 15460 12060 15492
rect 12094 15460 12160 15492
rect 12194 15460 12267 15492
rect 11573 15436 12267 15460
rect 11573 15402 11632 15436
rect 11666 15402 11722 15436
rect 11756 15402 11812 15436
rect 11846 15402 11902 15436
rect 11936 15402 11992 15436
rect 12026 15402 12082 15436
rect 12116 15402 12172 15436
rect 12206 15402 12267 15436
rect 11573 15394 12267 15402
rect 11573 15360 11660 15394
rect 11694 15360 11760 15394
rect 11794 15360 11860 15394
rect 11894 15360 11960 15394
rect 11994 15360 12060 15394
rect 12094 15360 12160 15394
rect 12194 15360 12267 15394
rect 11573 15346 12267 15360
rect 11573 15312 11632 15346
rect 11666 15312 11722 15346
rect 11756 15312 11812 15346
rect 11846 15312 11902 15346
rect 11936 15312 11992 15346
rect 12026 15312 12082 15346
rect 12116 15312 12172 15346
rect 12206 15312 12267 15346
rect 11573 15294 12267 15312
rect 11573 15260 11660 15294
rect 11694 15260 11760 15294
rect 11794 15260 11860 15294
rect 11894 15260 11960 15294
rect 11994 15260 12060 15294
rect 12094 15260 12160 15294
rect 12194 15260 12267 15294
rect 11573 15256 12267 15260
rect 11573 15222 11632 15256
rect 11666 15222 11722 15256
rect 11756 15222 11812 15256
rect 11846 15222 11902 15256
rect 11936 15222 11992 15256
rect 12026 15222 12082 15256
rect 12116 15222 12172 15256
rect 12206 15222 12267 15256
rect 11573 15194 12267 15222
rect 11573 15166 11660 15194
rect 11694 15166 11760 15194
rect 11573 15132 11632 15166
rect 11694 15160 11722 15166
rect 11666 15132 11722 15160
rect 11756 15160 11760 15166
rect 11794 15166 11860 15194
rect 11794 15160 11812 15166
rect 11756 15132 11812 15160
rect 11846 15160 11860 15166
rect 11894 15166 11960 15194
rect 11994 15166 12060 15194
rect 12094 15166 12160 15194
rect 12194 15166 12267 15194
rect 11894 15160 11902 15166
rect 11846 15132 11902 15160
rect 11936 15160 11960 15166
rect 12026 15160 12060 15166
rect 12116 15160 12160 15166
rect 11936 15132 11992 15160
rect 12026 15132 12082 15160
rect 12116 15132 12172 15160
rect 12206 15132 12267 15166
rect 11573 15073 12267 15132
rect 12329 15735 12348 15769
rect 12382 15735 12401 15769
rect 12329 15679 12401 15735
rect 12329 15645 12348 15679
rect 12382 15645 12401 15679
rect 12329 15589 12401 15645
rect 12329 15555 12348 15589
rect 12382 15555 12401 15589
rect 12329 15499 12401 15555
rect 12329 15465 12348 15499
rect 12382 15465 12401 15499
rect 12329 15409 12401 15465
rect 12329 15375 12348 15409
rect 12382 15375 12401 15409
rect 12329 15319 12401 15375
rect 12329 15285 12348 15319
rect 12382 15285 12401 15319
rect 12329 15229 12401 15285
rect 12329 15195 12348 15229
rect 12382 15195 12401 15229
rect 12329 15139 12401 15195
rect 12329 15105 12348 15139
rect 12382 15105 12401 15139
rect 11439 15034 11458 15068
rect 11492 15034 11511 15068
rect 11439 15020 11511 15034
rect 12329 15049 12401 15105
rect 12329 15020 12348 15049
rect 11343 15015 12348 15020
rect 12382 15020 12401 15049
rect 12465 15858 12735 15914
rect 13825 15948 14095 15965
rect 13825 15914 13856 15948
rect 13890 15914 14029 15948
rect 14063 15914 14095 15948
rect 12465 15824 12496 15858
rect 12530 15824 12669 15858
rect 12703 15824 12735 15858
rect 12465 15768 12735 15824
rect 12465 15734 12496 15768
rect 12530 15734 12669 15768
rect 12703 15734 12735 15768
rect 12465 15678 12735 15734
rect 12465 15644 12496 15678
rect 12530 15644 12669 15678
rect 12703 15644 12735 15678
rect 12465 15588 12735 15644
rect 12465 15554 12496 15588
rect 12530 15554 12669 15588
rect 12703 15554 12735 15588
rect 12465 15498 12735 15554
rect 12465 15464 12496 15498
rect 12530 15464 12669 15498
rect 12703 15464 12735 15498
rect 12465 15408 12735 15464
rect 12465 15374 12496 15408
rect 12530 15374 12669 15408
rect 12703 15374 12735 15408
rect 12465 15318 12735 15374
rect 12465 15284 12496 15318
rect 12530 15284 12669 15318
rect 12703 15284 12735 15318
rect 12465 15228 12735 15284
rect 12465 15194 12496 15228
rect 12530 15194 12669 15228
rect 12703 15194 12735 15228
rect 12465 15138 12735 15194
rect 12465 15104 12496 15138
rect 12530 15104 12669 15138
rect 12703 15104 12735 15138
rect 12465 15048 12735 15104
rect 12465 15020 12496 15048
rect 12382 15015 12496 15020
rect 11343 15014 12496 15015
rect 12530 15014 12669 15048
rect 12703 15020 12735 15048
rect 12799 15882 13761 15901
rect 12799 15848 12910 15882
rect 12944 15848 13000 15882
rect 13034 15848 13090 15882
rect 13124 15848 13180 15882
rect 13214 15848 13270 15882
rect 13304 15848 13360 15882
rect 13394 15848 13450 15882
rect 13484 15848 13540 15882
rect 13574 15848 13630 15882
rect 13664 15848 13761 15882
rect 12799 15829 13761 15848
rect 12799 15788 12871 15829
rect 12799 15754 12818 15788
rect 12852 15754 12871 15788
rect 13689 15769 13761 15829
rect 12799 15698 12871 15754
rect 12799 15664 12818 15698
rect 12852 15664 12871 15698
rect 12799 15608 12871 15664
rect 12799 15574 12818 15608
rect 12852 15574 12871 15608
rect 12799 15518 12871 15574
rect 12799 15484 12818 15518
rect 12852 15484 12871 15518
rect 12799 15428 12871 15484
rect 12799 15394 12818 15428
rect 12852 15394 12871 15428
rect 12799 15338 12871 15394
rect 12799 15304 12818 15338
rect 12852 15304 12871 15338
rect 12799 15248 12871 15304
rect 12799 15214 12818 15248
rect 12852 15214 12871 15248
rect 12799 15158 12871 15214
rect 12799 15124 12818 15158
rect 12852 15124 12871 15158
rect 12799 15068 12871 15124
rect 12933 15706 13627 15767
rect 12933 15672 12992 15706
rect 13026 15694 13082 15706
rect 13054 15672 13082 15694
rect 13116 15694 13172 15706
rect 13116 15672 13120 15694
rect 12933 15660 13020 15672
rect 13054 15660 13120 15672
rect 13154 15672 13172 15694
rect 13206 15694 13262 15706
rect 13206 15672 13220 15694
rect 13154 15660 13220 15672
rect 13254 15672 13262 15694
rect 13296 15694 13352 15706
rect 13386 15694 13442 15706
rect 13476 15694 13532 15706
rect 13296 15672 13320 15694
rect 13386 15672 13420 15694
rect 13476 15672 13520 15694
rect 13566 15672 13627 15706
rect 13254 15660 13320 15672
rect 13354 15660 13420 15672
rect 13454 15660 13520 15672
rect 13554 15660 13627 15672
rect 12933 15616 13627 15660
rect 12933 15582 12992 15616
rect 13026 15594 13082 15616
rect 13054 15582 13082 15594
rect 13116 15594 13172 15616
rect 13116 15582 13120 15594
rect 12933 15560 13020 15582
rect 13054 15560 13120 15582
rect 13154 15582 13172 15594
rect 13206 15594 13262 15616
rect 13206 15582 13220 15594
rect 13154 15560 13220 15582
rect 13254 15582 13262 15594
rect 13296 15594 13352 15616
rect 13386 15594 13442 15616
rect 13476 15594 13532 15616
rect 13296 15582 13320 15594
rect 13386 15582 13420 15594
rect 13476 15582 13520 15594
rect 13566 15582 13627 15616
rect 13254 15560 13320 15582
rect 13354 15560 13420 15582
rect 13454 15560 13520 15582
rect 13554 15560 13627 15582
rect 12933 15526 13627 15560
rect 12933 15492 12992 15526
rect 13026 15494 13082 15526
rect 13054 15492 13082 15494
rect 13116 15494 13172 15526
rect 13116 15492 13120 15494
rect 12933 15460 13020 15492
rect 13054 15460 13120 15492
rect 13154 15492 13172 15494
rect 13206 15494 13262 15526
rect 13206 15492 13220 15494
rect 13154 15460 13220 15492
rect 13254 15492 13262 15494
rect 13296 15494 13352 15526
rect 13386 15494 13442 15526
rect 13476 15494 13532 15526
rect 13296 15492 13320 15494
rect 13386 15492 13420 15494
rect 13476 15492 13520 15494
rect 13566 15492 13627 15526
rect 13254 15460 13320 15492
rect 13354 15460 13420 15492
rect 13454 15460 13520 15492
rect 13554 15460 13627 15492
rect 12933 15436 13627 15460
rect 12933 15402 12992 15436
rect 13026 15402 13082 15436
rect 13116 15402 13172 15436
rect 13206 15402 13262 15436
rect 13296 15402 13352 15436
rect 13386 15402 13442 15436
rect 13476 15402 13532 15436
rect 13566 15402 13627 15436
rect 12933 15394 13627 15402
rect 12933 15360 13020 15394
rect 13054 15360 13120 15394
rect 13154 15360 13220 15394
rect 13254 15360 13320 15394
rect 13354 15360 13420 15394
rect 13454 15360 13520 15394
rect 13554 15360 13627 15394
rect 12933 15346 13627 15360
rect 12933 15312 12992 15346
rect 13026 15312 13082 15346
rect 13116 15312 13172 15346
rect 13206 15312 13262 15346
rect 13296 15312 13352 15346
rect 13386 15312 13442 15346
rect 13476 15312 13532 15346
rect 13566 15312 13627 15346
rect 12933 15294 13627 15312
rect 12933 15260 13020 15294
rect 13054 15260 13120 15294
rect 13154 15260 13220 15294
rect 13254 15260 13320 15294
rect 13354 15260 13420 15294
rect 13454 15260 13520 15294
rect 13554 15260 13627 15294
rect 12933 15256 13627 15260
rect 12933 15222 12992 15256
rect 13026 15222 13082 15256
rect 13116 15222 13172 15256
rect 13206 15222 13262 15256
rect 13296 15222 13352 15256
rect 13386 15222 13442 15256
rect 13476 15222 13532 15256
rect 13566 15222 13627 15256
rect 12933 15194 13627 15222
rect 12933 15166 13020 15194
rect 13054 15166 13120 15194
rect 12933 15132 12992 15166
rect 13054 15160 13082 15166
rect 13026 15132 13082 15160
rect 13116 15160 13120 15166
rect 13154 15166 13220 15194
rect 13154 15160 13172 15166
rect 13116 15132 13172 15160
rect 13206 15160 13220 15166
rect 13254 15166 13320 15194
rect 13354 15166 13420 15194
rect 13454 15166 13520 15194
rect 13554 15166 13627 15194
rect 13254 15160 13262 15166
rect 13206 15132 13262 15160
rect 13296 15160 13320 15166
rect 13386 15160 13420 15166
rect 13476 15160 13520 15166
rect 13296 15132 13352 15160
rect 13386 15132 13442 15160
rect 13476 15132 13532 15160
rect 13566 15132 13627 15166
rect 12933 15073 13627 15132
rect 13689 15735 13708 15769
rect 13742 15735 13761 15769
rect 13689 15679 13761 15735
rect 13689 15645 13708 15679
rect 13742 15645 13761 15679
rect 13689 15589 13761 15645
rect 13689 15555 13708 15589
rect 13742 15555 13761 15589
rect 13689 15499 13761 15555
rect 13689 15465 13708 15499
rect 13742 15465 13761 15499
rect 13689 15409 13761 15465
rect 13689 15375 13708 15409
rect 13742 15375 13761 15409
rect 13689 15319 13761 15375
rect 13689 15285 13708 15319
rect 13742 15285 13761 15319
rect 13689 15229 13761 15285
rect 13689 15195 13708 15229
rect 13742 15195 13761 15229
rect 13689 15139 13761 15195
rect 13689 15105 13708 15139
rect 13742 15105 13761 15139
rect 12799 15034 12818 15068
rect 12852 15034 12871 15068
rect 12799 15020 12871 15034
rect 13689 15049 13761 15105
rect 13689 15020 13708 15049
rect 12703 15015 13708 15020
rect 13742 15020 13761 15049
rect 13825 15858 14095 15914
rect 15185 15948 15284 15965
rect 15185 15914 15216 15948
rect 15250 15914 15284 15948
rect 13825 15824 13856 15858
rect 13890 15824 14029 15858
rect 14063 15824 14095 15858
rect 13825 15768 14095 15824
rect 13825 15734 13856 15768
rect 13890 15734 14029 15768
rect 14063 15734 14095 15768
rect 13825 15678 14095 15734
rect 13825 15644 13856 15678
rect 13890 15644 14029 15678
rect 14063 15644 14095 15678
rect 13825 15588 14095 15644
rect 13825 15554 13856 15588
rect 13890 15554 14029 15588
rect 14063 15554 14095 15588
rect 13825 15498 14095 15554
rect 13825 15464 13856 15498
rect 13890 15464 14029 15498
rect 14063 15464 14095 15498
rect 13825 15408 14095 15464
rect 13825 15374 13856 15408
rect 13890 15374 14029 15408
rect 14063 15374 14095 15408
rect 13825 15318 14095 15374
rect 13825 15284 13856 15318
rect 13890 15284 14029 15318
rect 14063 15284 14095 15318
rect 13825 15228 14095 15284
rect 13825 15194 13856 15228
rect 13890 15194 14029 15228
rect 14063 15194 14095 15228
rect 13825 15138 14095 15194
rect 13825 15104 13856 15138
rect 13890 15104 14029 15138
rect 14063 15104 14095 15138
rect 13825 15048 14095 15104
rect 13825 15020 13856 15048
rect 13742 15015 13856 15020
rect 12703 15014 13856 15015
rect 13890 15014 14029 15048
rect 14063 15020 14095 15048
rect 14159 15882 15121 15901
rect 14159 15848 14270 15882
rect 14304 15848 14360 15882
rect 14394 15848 14450 15882
rect 14484 15848 14540 15882
rect 14574 15848 14630 15882
rect 14664 15848 14720 15882
rect 14754 15848 14810 15882
rect 14844 15848 14900 15882
rect 14934 15848 14990 15882
rect 15024 15848 15121 15882
rect 14159 15829 15121 15848
rect 14159 15788 14231 15829
rect 14159 15754 14178 15788
rect 14212 15754 14231 15788
rect 15049 15769 15121 15829
rect 14159 15698 14231 15754
rect 14159 15664 14178 15698
rect 14212 15664 14231 15698
rect 14159 15608 14231 15664
rect 14159 15574 14178 15608
rect 14212 15574 14231 15608
rect 14159 15518 14231 15574
rect 14159 15484 14178 15518
rect 14212 15484 14231 15518
rect 14159 15428 14231 15484
rect 14159 15394 14178 15428
rect 14212 15394 14231 15428
rect 14159 15338 14231 15394
rect 14159 15304 14178 15338
rect 14212 15304 14231 15338
rect 14159 15248 14231 15304
rect 14159 15214 14178 15248
rect 14212 15214 14231 15248
rect 14159 15158 14231 15214
rect 14159 15124 14178 15158
rect 14212 15124 14231 15158
rect 14159 15068 14231 15124
rect 14293 15706 14987 15767
rect 14293 15672 14352 15706
rect 14386 15694 14442 15706
rect 14414 15672 14442 15694
rect 14476 15694 14532 15706
rect 14476 15672 14480 15694
rect 14293 15660 14380 15672
rect 14414 15660 14480 15672
rect 14514 15672 14532 15694
rect 14566 15694 14622 15706
rect 14566 15672 14580 15694
rect 14514 15660 14580 15672
rect 14614 15672 14622 15694
rect 14656 15694 14712 15706
rect 14746 15694 14802 15706
rect 14836 15694 14892 15706
rect 14656 15672 14680 15694
rect 14746 15672 14780 15694
rect 14836 15672 14880 15694
rect 14926 15672 14987 15706
rect 14614 15660 14680 15672
rect 14714 15660 14780 15672
rect 14814 15660 14880 15672
rect 14914 15660 14987 15672
rect 14293 15616 14987 15660
rect 14293 15582 14352 15616
rect 14386 15594 14442 15616
rect 14414 15582 14442 15594
rect 14476 15594 14532 15616
rect 14476 15582 14480 15594
rect 14293 15560 14380 15582
rect 14414 15560 14480 15582
rect 14514 15582 14532 15594
rect 14566 15594 14622 15616
rect 14566 15582 14580 15594
rect 14514 15560 14580 15582
rect 14614 15582 14622 15594
rect 14656 15594 14712 15616
rect 14746 15594 14802 15616
rect 14836 15594 14892 15616
rect 14656 15582 14680 15594
rect 14746 15582 14780 15594
rect 14836 15582 14880 15594
rect 14926 15582 14987 15616
rect 14614 15560 14680 15582
rect 14714 15560 14780 15582
rect 14814 15560 14880 15582
rect 14914 15560 14987 15582
rect 14293 15526 14987 15560
rect 14293 15492 14352 15526
rect 14386 15494 14442 15526
rect 14414 15492 14442 15494
rect 14476 15494 14532 15526
rect 14476 15492 14480 15494
rect 14293 15460 14380 15492
rect 14414 15460 14480 15492
rect 14514 15492 14532 15494
rect 14566 15494 14622 15526
rect 14566 15492 14580 15494
rect 14514 15460 14580 15492
rect 14614 15492 14622 15494
rect 14656 15494 14712 15526
rect 14746 15494 14802 15526
rect 14836 15494 14892 15526
rect 14656 15492 14680 15494
rect 14746 15492 14780 15494
rect 14836 15492 14880 15494
rect 14926 15492 14987 15526
rect 14614 15460 14680 15492
rect 14714 15460 14780 15492
rect 14814 15460 14880 15492
rect 14914 15460 14987 15492
rect 14293 15436 14987 15460
rect 14293 15402 14352 15436
rect 14386 15402 14442 15436
rect 14476 15402 14532 15436
rect 14566 15402 14622 15436
rect 14656 15402 14712 15436
rect 14746 15402 14802 15436
rect 14836 15402 14892 15436
rect 14926 15402 14987 15436
rect 14293 15394 14987 15402
rect 14293 15360 14380 15394
rect 14414 15360 14480 15394
rect 14514 15360 14580 15394
rect 14614 15360 14680 15394
rect 14714 15360 14780 15394
rect 14814 15360 14880 15394
rect 14914 15360 14987 15394
rect 14293 15346 14987 15360
rect 14293 15312 14352 15346
rect 14386 15312 14442 15346
rect 14476 15312 14532 15346
rect 14566 15312 14622 15346
rect 14656 15312 14712 15346
rect 14746 15312 14802 15346
rect 14836 15312 14892 15346
rect 14926 15312 14987 15346
rect 14293 15294 14987 15312
rect 14293 15260 14380 15294
rect 14414 15260 14480 15294
rect 14514 15260 14580 15294
rect 14614 15260 14680 15294
rect 14714 15260 14780 15294
rect 14814 15260 14880 15294
rect 14914 15260 14987 15294
rect 14293 15256 14987 15260
rect 14293 15222 14352 15256
rect 14386 15222 14442 15256
rect 14476 15222 14532 15256
rect 14566 15222 14622 15256
rect 14656 15222 14712 15256
rect 14746 15222 14802 15256
rect 14836 15222 14892 15256
rect 14926 15222 14987 15256
rect 14293 15194 14987 15222
rect 14293 15166 14380 15194
rect 14414 15166 14480 15194
rect 14293 15132 14352 15166
rect 14414 15160 14442 15166
rect 14386 15132 14442 15160
rect 14476 15160 14480 15166
rect 14514 15166 14580 15194
rect 14514 15160 14532 15166
rect 14476 15132 14532 15160
rect 14566 15160 14580 15166
rect 14614 15166 14680 15194
rect 14714 15166 14780 15194
rect 14814 15166 14880 15194
rect 14914 15166 14987 15194
rect 14614 15160 14622 15166
rect 14566 15132 14622 15160
rect 14656 15160 14680 15166
rect 14746 15160 14780 15166
rect 14836 15160 14880 15166
rect 14656 15132 14712 15160
rect 14746 15132 14802 15160
rect 14836 15132 14892 15160
rect 14926 15132 14987 15166
rect 14293 15073 14987 15132
rect 15049 15735 15068 15769
rect 15102 15735 15121 15769
rect 15049 15679 15121 15735
rect 15049 15645 15068 15679
rect 15102 15645 15121 15679
rect 15049 15589 15121 15645
rect 15049 15555 15068 15589
rect 15102 15555 15121 15589
rect 15049 15499 15121 15555
rect 15049 15465 15068 15499
rect 15102 15465 15121 15499
rect 15049 15409 15121 15465
rect 15049 15375 15068 15409
rect 15102 15375 15121 15409
rect 15049 15319 15121 15375
rect 15049 15285 15068 15319
rect 15102 15285 15121 15319
rect 15049 15229 15121 15285
rect 15049 15195 15068 15229
rect 15102 15195 15121 15229
rect 15049 15139 15121 15195
rect 15049 15105 15068 15139
rect 15102 15105 15121 15139
rect 14159 15034 14178 15068
rect 14212 15034 14231 15068
rect 14159 15020 14231 15034
rect 15049 15049 15121 15105
rect 15049 15020 15068 15049
rect 14063 15015 15068 15020
rect 15102 15020 15121 15049
rect 15185 15858 15284 15914
rect 15185 15824 15216 15858
rect 15250 15824 15284 15858
rect 15185 15768 15284 15824
rect 17011 18499 17045 18561
rect 16593 15847 16627 15909
rect 17383 18555 17479 18589
rect 17739 18555 17835 18589
rect 17383 18493 17417 18555
rect 17570 18550 17590 18555
rect 17630 18550 17650 18555
rect 17570 18530 17650 18550
rect 17801 18493 17835 18555
rect 17383 16527 17417 16589
rect 17801 16527 17835 16589
rect 17383 16493 17479 16527
rect 17739 16493 17835 16527
rect 17011 15847 17045 15909
rect 16593 15813 16689 15847
rect 16949 15813 17045 15847
rect 15185 15734 15216 15768
rect 15250 15734 15284 15768
rect 15185 15678 15284 15734
rect 15185 15644 15216 15678
rect 15250 15644 15284 15678
rect 15185 15588 15284 15644
rect 15185 15554 15216 15588
rect 15250 15554 15284 15588
rect 15185 15498 15284 15554
rect 15185 15464 15216 15498
rect 15250 15464 15284 15498
rect 15185 15408 15284 15464
rect 15185 15374 15216 15408
rect 15250 15374 15284 15408
rect 15185 15318 15284 15374
rect 15185 15284 15216 15318
rect 15250 15284 15284 15318
rect 15185 15228 15284 15284
rect 15185 15194 15216 15228
rect 15250 15194 15284 15228
rect 15185 15138 15284 15194
rect 15185 15104 15216 15138
rect 15250 15104 15284 15138
rect 15185 15048 15284 15104
rect 15185 15020 15216 15048
rect 15102 15015 15216 15020
rect 14063 15014 15216 15015
rect 15250 15020 15284 15048
rect 15250 15014 15290 15020
rect 11270 14992 15290 15014
rect 11270 14958 11516 14992
rect 11550 14958 11606 14992
rect 11640 14958 11696 14992
rect 11730 14958 11786 14992
rect 11820 14958 11876 14992
rect 11910 14958 11966 14992
rect 12000 14958 12056 14992
rect 12090 14958 12146 14992
rect 12180 14958 12236 14992
rect 12270 14958 12876 14992
rect 12910 14958 12966 14992
rect 13000 14958 13056 14992
rect 13090 14958 13146 14992
rect 13180 14958 13236 14992
rect 13270 14958 13326 14992
rect 13360 14958 13416 14992
rect 13450 14958 13506 14992
rect 13540 14958 13596 14992
rect 13630 14958 14236 14992
rect 14270 14958 14326 14992
rect 14360 14958 14416 14992
rect 14450 14958 14506 14992
rect 14540 14958 14596 14992
rect 14630 14958 14686 14992
rect 14720 14958 14776 14992
rect 14810 14958 14866 14992
rect 14900 14958 14956 14992
rect 14990 14958 15290 14992
rect 11270 14924 11309 14958
rect 11343 14924 12496 14958
rect 12530 14924 12669 14958
rect 12703 14924 13856 14958
rect 13890 14924 14029 14958
rect 14063 14924 15216 14958
rect 15250 14924 15290 14958
rect 11270 14868 15290 14924
rect 11270 14834 11309 14868
rect 11343 14845 12496 14868
rect 11343 14834 11410 14845
rect 11270 14811 11410 14834
rect 11444 14811 11500 14845
rect 11534 14811 11590 14845
rect 11624 14811 11680 14845
rect 11714 14811 11770 14845
rect 11804 14811 11860 14845
rect 11894 14811 11950 14845
rect 11984 14811 12040 14845
rect 12074 14811 12130 14845
rect 12164 14811 12220 14845
rect 12254 14811 12310 14845
rect 12344 14811 12400 14845
rect 12434 14834 12496 14845
rect 12530 14834 12669 14868
rect 12703 14845 13856 14868
rect 12703 14834 12770 14845
rect 12434 14811 12770 14834
rect 12804 14811 12860 14845
rect 12894 14811 12950 14845
rect 12984 14811 13040 14845
rect 13074 14811 13130 14845
rect 13164 14811 13220 14845
rect 13254 14811 13310 14845
rect 13344 14811 13400 14845
rect 13434 14811 13490 14845
rect 13524 14811 13580 14845
rect 13614 14811 13670 14845
rect 13704 14811 13760 14845
rect 13794 14834 13856 14845
rect 13890 14834 14029 14868
rect 14063 14845 15216 14868
rect 14063 14834 14130 14845
rect 13794 14811 14130 14834
rect 14164 14811 14220 14845
rect 14254 14811 14310 14845
rect 14344 14811 14400 14845
rect 14434 14811 14490 14845
rect 14524 14811 14580 14845
rect 14614 14811 14670 14845
rect 14704 14811 14760 14845
rect 14794 14811 14850 14845
rect 14884 14811 14940 14845
rect 14974 14811 15030 14845
rect 15064 14811 15120 14845
rect 15154 14834 15216 14845
rect 15250 14834 15290 14868
rect 15154 14811 15290 14834
rect 11270 14770 15290 14811
rect 11403 14571 11499 14605
rect 15057 14571 15153 14605
rect 11403 14509 11437 14571
rect 15119 14509 15153 14571
rect 11403 14187 11437 14249
rect 15119 14187 15153 14249
rect 11403 14153 11499 14187
rect 15057 14153 15153 14187
rect 11170 13850 11230 13870
rect 11170 13820 11180 13850
rect 11080 13810 11180 13820
rect 11220 13810 11230 13850
rect 11080 13800 11230 13810
rect 11080 13760 11100 13800
rect 11140 13760 11230 13800
rect 11080 13750 11230 13760
rect 11080 13740 11180 13750
rect 11170 13710 11180 13740
rect 11220 13710 11230 13750
rect 11170 13690 11230 13710
rect 13250 13850 13310 13870
rect 13250 13810 13260 13850
rect 13300 13810 13310 13850
rect 13250 13750 13310 13810
rect 13250 13710 13260 13750
rect 13300 13710 13310 13750
rect 13250 13690 13310 13710
rect 15330 13860 15470 13870
rect 15330 13850 15550 13860
rect 15330 13810 15340 13850
rect 15380 13810 15420 13850
rect 15460 13840 15550 13850
rect 15460 13810 15490 13840
rect 15330 13800 15490 13810
rect 15530 13800 15550 13840
rect 15330 13760 15550 13800
rect 15330 13750 15490 13760
rect 15330 13710 15340 13750
rect 15380 13710 15420 13750
rect 15460 13720 15490 13750
rect 15530 13720 15550 13760
rect 15460 13710 15550 13720
rect 15330 13700 15550 13710
rect 15330 13690 15470 13700
rect 11180 13650 11220 13690
rect 13260 13650 13300 13690
rect 11160 13630 11240 13650
rect 11160 13590 11180 13630
rect 11220 13590 11240 13630
rect 11160 13570 11240 13590
rect 11320 13630 11400 13650
rect 11320 13590 11340 13630
rect 11380 13590 11400 13630
rect 11320 13570 11400 13590
rect 11480 13630 11560 13650
rect 11480 13590 11500 13630
rect 11540 13590 11560 13630
rect 11480 13570 11560 13590
rect 11640 13630 11720 13650
rect 11640 13590 11660 13630
rect 11700 13590 11720 13630
rect 11640 13570 11720 13590
rect 11800 13630 11880 13650
rect 11800 13590 11820 13630
rect 11860 13590 11880 13630
rect 11800 13570 11880 13590
rect 11960 13630 12040 13650
rect 11960 13590 11980 13630
rect 12020 13590 12040 13630
rect 11960 13570 12040 13590
rect 12120 13630 12200 13650
rect 12120 13590 12140 13630
rect 12180 13590 12200 13630
rect 12120 13570 12200 13590
rect 12280 13630 12360 13650
rect 12280 13590 12300 13630
rect 12340 13590 12360 13630
rect 12280 13570 12360 13590
rect 12440 13630 12520 13650
rect 12440 13590 12460 13630
rect 12500 13590 12520 13630
rect 12440 13570 12520 13590
rect 12600 13630 12680 13650
rect 12600 13590 12620 13630
rect 12660 13590 12680 13630
rect 12600 13570 12680 13590
rect 12760 13630 12840 13650
rect 12760 13590 12780 13630
rect 12820 13590 12840 13630
rect 12760 13570 12840 13590
rect 12920 13630 13000 13650
rect 12920 13590 12940 13630
rect 12980 13590 13000 13630
rect 12920 13570 13000 13590
rect 13080 13630 13160 13650
rect 13080 13590 13100 13630
rect 13140 13590 13160 13630
rect 13080 13570 13160 13590
rect 13240 13630 13320 13650
rect 13240 13590 13260 13630
rect 13300 13590 13320 13630
rect 13240 13570 13320 13590
rect 13400 13630 13480 13650
rect 13400 13590 13420 13630
rect 13460 13590 13480 13630
rect 13400 13570 13480 13590
rect 13560 13630 13640 13650
rect 13560 13590 13580 13630
rect 13620 13590 13640 13630
rect 13560 13570 13640 13590
rect 13720 13630 13800 13650
rect 13720 13590 13740 13630
rect 13780 13590 13800 13630
rect 13720 13570 13800 13590
rect 13880 13630 13960 13650
rect 13880 13590 13900 13630
rect 13940 13590 13960 13630
rect 13880 13570 13960 13590
rect 14040 13630 14120 13650
rect 14040 13590 14060 13630
rect 14100 13590 14120 13630
rect 14040 13570 14120 13590
rect 14200 13630 14280 13650
rect 14200 13590 14220 13630
rect 14260 13590 14280 13630
rect 14200 13570 14280 13590
rect 14360 13630 14440 13650
rect 14360 13590 14380 13630
rect 14420 13590 14440 13630
rect 14360 13570 14440 13590
rect 14520 13630 14600 13650
rect 14520 13590 14540 13630
rect 14580 13590 14600 13630
rect 14520 13570 14600 13590
rect 14680 13630 14760 13650
rect 14680 13590 14700 13630
rect 14740 13590 14760 13630
rect 14680 13570 14760 13590
rect 14840 13630 14920 13650
rect 14840 13590 14860 13630
rect 14900 13590 14920 13630
rect 14840 13570 14920 13590
rect 15000 13630 15080 13650
rect 15000 13590 15020 13630
rect 15060 13590 15080 13630
rect 15000 13570 15080 13590
rect 15160 13630 15240 13650
rect 15160 13590 15180 13630
rect 15220 13590 15240 13630
rect 15160 13570 15240 13590
rect 11900 13360 11980 13380
rect 11900 13320 11920 13360
rect 11960 13320 11980 13360
rect 11900 13260 11980 13320
rect 14580 13360 14660 13380
rect 14580 13320 14600 13360
rect 14640 13320 14660 13360
rect 14580 13260 14660 13320
rect 10750 13240 10810 13260
rect 10750 13200 10760 13240
rect 10800 13200 10810 13240
rect 10750 13140 10810 13200
rect 10750 13100 10760 13140
rect 10800 13100 10810 13140
rect 10750 13040 10810 13100
rect 10750 13000 10760 13040
rect 10800 13000 10810 13040
rect 10750 12940 10810 13000
rect 10750 12900 10760 12940
rect 10800 12900 10810 12940
rect 10750 12840 10810 12900
rect 10750 12800 10760 12840
rect 10800 12800 10810 12840
rect 10750 12780 10810 12800
rect 11830 13240 12050 13260
rect 11830 13200 11840 13240
rect 11880 13200 11920 13240
rect 11960 13200 12000 13240
rect 12040 13200 12050 13240
rect 11830 13140 12050 13200
rect 11830 13100 11840 13140
rect 11880 13100 11920 13140
rect 11960 13100 12000 13140
rect 12040 13100 12050 13140
rect 11830 13040 12050 13100
rect 11830 13000 11840 13040
rect 11880 13000 11920 13040
rect 11960 13000 12000 13040
rect 12040 13000 12050 13040
rect 11830 12940 12050 13000
rect 11830 12900 11840 12940
rect 11880 12900 11920 12940
rect 11960 12900 12000 12940
rect 12040 12900 12050 12940
rect 11830 12840 12050 12900
rect 11830 12800 11840 12840
rect 11880 12800 11920 12840
rect 11960 12800 12000 12840
rect 12040 12800 12050 12840
rect 11830 12780 12050 12800
rect 13070 13240 13130 13260
rect 13070 13200 13080 13240
rect 13120 13200 13130 13240
rect 13070 13140 13130 13200
rect 13070 13100 13080 13140
rect 13120 13100 13130 13140
rect 13070 13040 13130 13100
rect 13070 13000 13080 13040
rect 13120 13000 13130 13040
rect 13070 12940 13130 13000
rect 13070 12900 13080 12940
rect 13120 12900 13130 12940
rect 13070 12840 13130 12900
rect 13070 12800 13080 12840
rect 13120 12800 13130 12840
rect 10740 12760 10820 12780
rect 10740 12720 10760 12760
rect 10800 12720 10820 12760
rect 13070 12750 13130 12800
rect 10740 12700 10820 12720
rect 10920 12720 11000 12740
rect 10920 12680 10940 12720
rect 10980 12680 11000 12720
rect 10920 12660 11000 12680
rect 11160 12720 11240 12740
rect 11160 12680 11180 12720
rect 11220 12680 11240 12720
rect 11160 12660 11240 12680
rect 11400 12720 11480 12740
rect 11400 12680 11420 12720
rect 11460 12680 11480 12720
rect 11400 12660 11480 12680
rect 11640 12720 11720 12740
rect 11640 12680 11660 12720
rect 11700 12680 11720 12720
rect 11640 12660 11720 12680
rect 12280 12720 12360 12740
rect 12280 12680 12300 12720
rect 12340 12680 12360 12720
rect 12280 12660 12360 12680
rect 12520 12720 12600 12740
rect 12520 12680 12540 12720
rect 12580 12680 12600 12720
rect 12520 12660 12600 12680
rect 12760 12720 12840 12740
rect 12760 12680 12780 12720
rect 12820 12680 12840 12720
rect 13070 12710 13080 12750
rect 13120 12710 13130 12750
rect 13070 12690 13130 12710
rect 13430 13240 13490 13260
rect 13430 13200 13440 13240
rect 13480 13200 13490 13240
rect 13430 13140 13490 13200
rect 13430 13100 13440 13140
rect 13480 13100 13490 13140
rect 13430 13040 13490 13100
rect 13430 13000 13440 13040
rect 13480 13000 13490 13040
rect 13430 12940 13490 13000
rect 13430 12900 13440 12940
rect 13480 12900 13490 12940
rect 13430 12840 13490 12900
rect 13430 12800 13440 12840
rect 13480 12800 13490 12840
rect 13430 12750 13490 12800
rect 14510 13240 14730 13260
rect 14510 13200 14520 13240
rect 14560 13200 14600 13240
rect 14640 13200 14680 13240
rect 14720 13200 14730 13240
rect 14510 13140 14730 13200
rect 14510 13100 14520 13140
rect 14560 13100 14600 13140
rect 14640 13100 14680 13140
rect 14720 13100 14730 13140
rect 14510 13040 14730 13100
rect 14510 13000 14520 13040
rect 14560 13000 14600 13040
rect 14640 13000 14680 13040
rect 14720 13000 14730 13040
rect 14510 12940 14730 13000
rect 14510 12900 14520 12940
rect 14560 12900 14600 12940
rect 14640 12900 14680 12940
rect 14720 12900 14730 12940
rect 14510 12840 14730 12900
rect 14510 12800 14520 12840
rect 14560 12800 14600 12840
rect 14640 12800 14680 12840
rect 14720 12800 14730 12840
rect 14510 12780 14730 12800
rect 15750 13240 15810 13260
rect 15750 13200 15760 13240
rect 15800 13200 15810 13240
rect 15750 13140 15810 13200
rect 15750 13100 15760 13140
rect 15800 13100 15810 13140
rect 15750 13040 15810 13100
rect 15750 13000 15760 13040
rect 15800 13000 15810 13040
rect 15750 12940 15810 13000
rect 15750 12900 15760 12940
rect 15800 12900 15810 12940
rect 15750 12840 15810 12900
rect 15750 12800 15760 12840
rect 15800 12800 15810 12840
rect 15750 12780 15810 12800
rect 13430 12710 13440 12750
rect 13480 12710 13490 12750
rect 13430 12690 13490 12710
rect 13720 12720 13800 12740
rect 12760 12660 12840 12680
rect 13720 12680 13740 12720
rect 13780 12680 13800 12720
rect 13720 12660 13800 12680
rect 13960 12720 14040 12740
rect 13960 12680 13980 12720
rect 14020 12680 14040 12720
rect 13960 12660 14040 12680
rect 14200 12720 14280 12740
rect 14200 12680 14220 12720
rect 14260 12680 14280 12720
rect 14200 12660 14280 12680
rect 14840 12720 14920 12740
rect 14840 12680 14860 12720
rect 14900 12680 14920 12720
rect 14840 12660 14920 12680
rect 15080 12720 15160 12740
rect 15080 12680 15100 12720
rect 15140 12680 15160 12720
rect 15080 12660 15160 12680
rect 15320 12720 15400 12740
rect 15320 12680 15340 12720
rect 15380 12680 15400 12720
rect 15320 12660 15400 12680
rect 15560 12720 15640 12740
rect 15560 12680 15580 12720
rect 15620 12680 15640 12720
rect 15560 12660 15640 12680
rect 11431 12342 11489 12360
rect 11431 12308 11443 12342
rect 11477 12308 11489 12342
rect 11431 12290 11489 12308
rect 11791 12342 11849 12360
rect 11791 12308 11803 12342
rect 11837 12308 11849 12342
rect 11791 12290 11849 12308
rect 11911 12342 11969 12360
rect 11911 12308 11923 12342
rect 11957 12308 11969 12342
rect 11911 12290 11969 12308
rect 12271 12342 12329 12360
rect 12271 12308 12283 12342
rect 12317 12308 12329 12342
rect 12271 12290 12329 12308
rect 12391 12342 12449 12360
rect 12391 12308 12403 12342
rect 12437 12308 12449 12342
rect 14111 12342 14169 12360
rect 12391 12290 12449 12308
rect 12800 12320 12880 12340
rect 12800 12280 12820 12320
rect 12860 12280 12880 12320
rect 11370 12230 11430 12250
rect 11370 12190 11380 12230
rect 11420 12190 11430 12230
rect 11370 12170 11430 12190
rect 11490 12230 11550 12250
rect 11490 12190 11500 12230
rect 11540 12190 11550 12230
rect 11490 12170 11550 12190
rect 11610 12230 11670 12250
rect 11610 12190 11620 12230
rect 11660 12190 11670 12230
rect 11610 12170 11670 12190
rect 11730 12230 11790 12250
rect 11730 12190 11740 12230
rect 11780 12190 11790 12230
rect 11730 12170 11790 12190
rect 11850 12230 11910 12250
rect 11850 12190 11860 12230
rect 11900 12190 11910 12230
rect 11850 12170 11910 12190
rect 11970 12230 12030 12250
rect 11970 12190 11980 12230
rect 12020 12190 12030 12230
rect 11970 12170 12030 12190
rect 12090 12230 12150 12250
rect 12090 12190 12100 12230
rect 12140 12190 12150 12230
rect 12090 12170 12150 12190
rect 12210 12230 12270 12250
rect 12210 12190 12220 12230
rect 12260 12190 12270 12230
rect 12210 12170 12270 12190
rect 12330 12230 12390 12250
rect 12330 12190 12340 12230
rect 12380 12190 12390 12230
rect 12330 12170 12390 12190
rect 12450 12230 12510 12250
rect 12450 12190 12460 12230
rect 12500 12190 12510 12230
rect 12450 12170 12510 12190
rect 12570 12230 12630 12250
rect 12570 12190 12580 12230
rect 12620 12190 12630 12230
rect 12570 12170 12630 12190
rect 12800 12240 12880 12280
rect 12800 12200 12820 12240
rect 12860 12200 12880 12240
rect 12800 12160 12880 12200
rect 11532 12112 11590 12130
rect 11532 12078 11544 12112
rect 11578 12078 11590 12112
rect 11532 12060 11590 12078
rect 11690 12112 11748 12130
rect 11690 12078 11702 12112
rect 11736 12078 11748 12112
rect 11690 12060 11748 12078
rect 12014 12112 12072 12130
rect 12014 12078 12026 12112
rect 12060 12078 12072 12112
rect 12014 12060 12072 12078
rect 12168 12112 12226 12130
rect 12168 12078 12180 12112
rect 12214 12078 12226 12112
rect 12168 12060 12226 12078
rect 12492 12112 12550 12130
rect 12492 12078 12504 12112
rect 12538 12078 12550 12112
rect 12800 12120 12820 12160
rect 12860 12120 12880 12160
rect 12800 12100 12880 12120
rect 13680 12320 13760 12340
rect 13680 12280 13700 12320
rect 13740 12280 13760 12320
rect 14111 12308 14123 12342
rect 14157 12308 14169 12342
rect 14111 12290 14169 12308
rect 14231 12342 14289 12360
rect 14231 12308 14243 12342
rect 14277 12308 14289 12342
rect 14231 12290 14289 12308
rect 14591 12342 14649 12360
rect 14591 12308 14603 12342
rect 14637 12308 14649 12342
rect 14591 12290 14649 12308
rect 14711 12342 14769 12360
rect 14711 12308 14723 12342
rect 14757 12308 14769 12342
rect 14711 12290 14769 12308
rect 15071 12342 15129 12360
rect 15071 12308 15083 12342
rect 15117 12308 15129 12342
rect 15071 12290 15129 12308
rect 13680 12240 13760 12280
rect 13680 12200 13700 12240
rect 13740 12200 13760 12240
rect 13680 12160 13760 12200
rect 13930 12230 13990 12250
rect 13930 12190 13940 12230
rect 13980 12190 13990 12230
rect 13930 12170 13990 12190
rect 14050 12230 14110 12250
rect 14050 12190 14060 12230
rect 14100 12190 14110 12230
rect 14050 12170 14110 12190
rect 14170 12230 14230 12250
rect 14170 12190 14180 12230
rect 14220 12190 14230 12230
rect 14170 12170 14230 12190
rect 14290 12230 14350 12250
rect 14290 12190 14300 12230
rect 14340 12190 14350 12230
rect 14290 12170 14350 12190
rect 14410 12230 14470 12250
rect 14410 12190 14420 12230
rect 14460 12190 14470 12230
rect 14410 12170 14470 12190
rect 14530 12230 14590 12250
rect 14530 12190 14540 12230
rect 14580 12190 14590 12230
rect 14530 12170 14590 12190
rect 14650 12230 14710 12250
rect 14650 12190 14660 12230
rect 14700 12190 14710 12230
rect 14650 12170 14710 12190
rect 14770 12230 14830 12250
rect 14770 12190 14780 12230
rect 14820 12190 14830 12230
rect 14770 12170 14830 12190
rect 14890 12230 14950 12250
rect 14890 12190 14900 12230
rect 14940 12190 14950 12230
rect 14890 12170 14950 12190
rect 15010 12230 15070 12250
rect 15010 12190 15020 12230
rect 15060 12190 15070 12230
rect 15010 12170 15070 12190
rect 15130 12230 15190 12250
rect 15130 12190 15140 12230
rect 15180 12190 15190 12230
rect 15130 12170 15190 12190
rect 13680 12120 13700 12160
rect 13740 12120 13760 12160
rect 13680 12100 13760 12120
rect 14010 12112 14068 12130
rect 12492 12060 12550 12078
rect 14010 12078 14022 12112
rect 14056 12078 14068 12112
rect 14010 12060 14068 12078
rect 14334 12112 14392 12130
rect 14334 12078 14346 12112
rect 14380 12078 14392 12112
rect 14334 12060 14392 12078
rect 14488 12112 14546 12130
rect 14488 12078 14500 12112
rect 14534 12078 14546 12112
rect 14488 12060 14546 12078
rect 14812 12112 14870 12130
rect 14812 12078 14824 12112
rect 14858 12078 14870 12112
rect 14812 12060 14870 12078
rect 14970 12112 15028 12130
rect 14970 12078 14982 12112
rect 15016 12078 15028 12112
rect 14970 12060 15028 12078
rect 10710 11520 10770 11540
rect 10710 11480 10720 11520
rect 10760 11480 10770 11520
rect 10710 11460 10770 11480
rect 10880 11510 10960 11530
rect 10880 11470 10900 11510
rect 10940 11470 10960 11510
rect 10880 11450 10960 11470
rect 11370 11510 11430 11530
rect 11370 11470 11380 11510
rect 11420 11470 11430 11510
rect 11370 11450 11430 11470
rect 11600 11510 11680 11530
rect 11600 11470 11620 11510
rect 11660 11470 11680 11510
rect 11600 11450 11680 11470
rect 12090 11510 12150 11530
rect 12090 11470 12100 11510
rect 12140 11470 12150 11510
rect 12090 11450 12150 11470
rect 12320 11510 12400 11530
rect 12320 11470 12340 11510
rect 12380 11470 12400 11510
rect 12320 11450 12400 11470
rect 12750 11510 12810 11530
rect 12750 11470 12760 11510
rect 12800 11470 12810 11510
rect 12750 11450 12810 11470
rect 13750 11510 13810 11530
rect 13750 11470 13760 11510
rect 13800 11470 13810 11510
rect 13750 11450 13810 11470
rect 14160 11510 14240 11530
rect 14160 11470 14180 11510
rect 14220 11470 14240 11510
rect 14160 11450 14240 11470
rect 14410 11510 14470 11530
rect 14410 11470 14420 11510
rect 14460 11470 14470 11510
rect 14410 11450 14470 11470
rect 14880 11510 14960 11530
rect 14880 11470 14900 11510
rect 14940 11470 14960 11510
rect 14880 11450 14960 11470
rect 15130 11510 15190 11530
rect 15130 11470 15140 11510
rect 15180 11470 15190 11510
rect 15130 11450 15190 11470
rect 15600 11510 15680 11530
rect 15600 11470 15620 11510
rect 15660 11470 15680 11510
rect 15600 11450 15680 11470
rect 15790 11520 15850 11540
rect 15790 11480 15800 11520
rect 15840 11480 15850 11520
rect 15790 11460 15850 11480
rect 10450 11390 10590 11410
rect 10450 11350 10460 11390
rect 10500 11350 10540 11390
rect 10580 11350 10590 11390
rect 10450 11290 10590 11350
rect 10450 11250 10460 11290
rect 10500 11250 10540 11290
rect 10580 11250 10590 11290
rect 10450 11230 10590 11250
rect 10650 11390 10710 11410
rect 10650 11350 10660 11390
rect 10700 11350 10710 11390
rect 10650 11290 10710 11350
rect 10650 11250 10660 11290
rect 10700 11250 10710 11290
rect 10650 11230 10710 11250
rect 10770 11390 10830 11410
rect 10770 11350 10780 11390
rect 10820 11350 10830 11390
rect 10770 11290 10830 11350
rect 10770 11250 10780 11290
rect 10820 11250 10830 11290
rect 10770 11230 10830 11250
rect 10890 11390 10950 11410
rect 10890 11350 10900 11390
rect 10940 11350 10950 11390
rect 10890 11290 10950 11350
rect 10890 11250 10900 11290
rect 10940 11250 10950 11290
rect 10890 11230 10950 11250
rect 11010 11390 11070 11410
rect 11010 11350 11020 11390
rect 11060 11350 11070 11390
rect 11010 11290 11070 11350
rect 11010 11250 11020 11290
rect 11060 11250 11070 11290
rect 11010 11230 11070 11250
rect 11130 11390 11190 11410
rect 11130 11350 11140 11390
rect 11180 11350 11190 11390
rect 11130 11290 11190 11350
rect 11130 11250 11140 11290
rect 11180 11250 11190 11290
rect 11130 11230 11190 11250
rect 11250 11390 11310 11410
rect 11250 11350 11260 11390
rect 11300 11350 11310 11390
rect 11250 11290 11310 11350
rect 11250 11250 11260 11290
rect 11300 11250 11310 11290
rect 11250 11230 11310 11250
rect 11370 11390 11430 11410
rect 11370 11350 11380 11390
rect 11420 11350 11430 11390
rect 11370 11290 11430 11350
rect 11370 11250 11380 11290
rect 11420 11250 11430 11290
rect 11370 11230 11430 11250
rect 11490 11390 11550 11410
rect 11490 11350 11500 11390
rect 11540 11350 11550 11390
rect 11490 11290 11550 11350
rect 11490 11250 11500 11290
rect 11540 11250 11550 11290
rect 11490 11230 11550 11250
rect 11610 11390 11670 11410
rect 11610 11350 11620 11390
rect 11660 11350 11670 11390
rect 11610 11290 11670 11350
rect 11610 11250 11620 11290
rect 11660 11250 11670 11290
rect 11610 11230 11670 11250
rect 11730 11390 11790 11410
rect 11730 11350 11740 11390
rect 11780 11350 11790 11390
rect 11730 11290 11790 11350
rect 11730 11250 11740 11290
rect 11780 11250 11790 11290
rect 11730 11230 11790 11250
rect 11850 11390 11910 11410
rect 11850 11350 11860 11390
rect 11900 11350 11910 11390
rect 11850 11290 11910 11350
rect 11850 11250 11860 11290
rect 11900 11250 11910 11290
rect 11850 11230 11910 11250
rect 11970 11390 12030 11410
rect 11970 11350 11980 11390
rect 12020 11350 12030 11390
rect 11970 11290 12030 11350
rect 11970 11250 11980 11290
rect 12020 11250 12030 11290
rect 11970 11230 12030 11250
rect 12090 11390 12150 11410
rect 12090 11350 12100 11390
rect 12140 11350 12150 11390
rect 12090 11290 12150 11350
rect 12090 11250 12100 11290
rect 12140 11250 12150 11290
rect 12090 11230 12150 11250
rect 12210 11390 12270 11410
rect 12210 11350 12220 11390
rect 12260 11350 12270 11390
rect 12210 11290 12270 11350
rect 12210 11250 12220 11290
rect 12260 11250 12270 11290
rect 12210 11230 12270 11250
rect 12330 11390 12390 11410
rect 12330 11350 12340 11390
rect 12380 11350 12390 11390
rect 12330 11290 12390 11350
rect 12330 11250 12340 11290
rect 12380 11250 12390 11290
rect 12330 11230 12390 11250
rect 12450 11390 12510 11410
rect 12450 11350 12460 11390
rect 12500 11350 12510 11390
rect 12450 11290 12510 11350
rect 12450 11250 12460 11290
rect 12500 11250 12510 11290
rect 12450 11230 12510 11250
rect 12570 11390 12630 11410
rect 12570 11350 12580 11390
rect 12620 11350 12630 11390
rect 12570 11290 12630 11350
rect 12570 11250 12580 11290
rect 12620 11250 12630 11290
rect 12570 11230 12630 11250
rect 12690 11390 12750 11410
rect 12690 11350 12700 11390
rect 12740 11350 12750 11390
rect 12690 11290 12750 11350
rect 12690 11250 12700 11290
rect 12740 11250 12750 11290
rect 12690 11230 12750 11250
rect 12810 11390 12870 11410
rect 12810 11350 12820 11390
rect 12860 11350 12870 11390
rect 12810 11290 12870 11350
rect 12810 11250 12820 11290
rect 12860 11250 12870 11290
rect 12810 11230 12870 11250
rect 12930 11390 13070 11410
rect 12930 11350 12940 11390
rect 12980 11350 13020 11390
rect 13060 11350 13070 11390
rect 12930 11290 13070 11350
rect 12930 11250 12940 11290
rect 12980 11250 13020 11290
rect 13060 11250 13070 11290
rect 12930 11230 13070 11250
rect 13490 11390 13630 11410
rect 13490 11350 13500 11390
rect 13540 11350 13580 11390
rect 13620 11350 13630 11390
rect 13490 11290 13630 11350
rect 13490 11250 13500 11290
rect 13540 11250 13580 11290
rect 13620 11250 13630 11290
rect 13490 11230 13630 11250
rect 13690 11390 13750 11410
rect 13690 11350 13700 11390
rect 13740 11350 13750 11390
rect 13690 11290 13750 11350
rect 13690 11250 13700 11290
rect 13740 11250 13750 11290
rect 13690 11230 13750 11250
rect 13810 11390 13870 11410
rect 13810 11350 13820 11390
rect 13860 11350 13870 11390
rect 13810 11290 13870 11350
rect 13810 11250 13820 11290
rect 13860 11250 13870 11290
rect 13810 11230 13870 11250
rect 13930 11390 13990 11410
rect 13930 11350 13940 11390
rect 13980 11350 13990 11390
rect 13930 11290 13990 11350
rect 13930 11250 13940 11290
rect 13980 11250 13990 11290
rect 13930 11230 13990 11250
rect 14050 11390 14110 11410
rect 14050 11350 14060 11390
rect 14100 11350 14110 11390
rect 14050 11290 14110 11350
rect 14050 11250 14060 11290
rect 14100 11250 14110 11290
rect 14050 11230 14110 11250
rect 14170 11390 14230 11410
rect 14170 11350 14180 11390
rect 14220 11350 14230 11390
rect 14170 11290 14230 11350
rect 14170 11250 14180 11290
rect 14220 11250 14230 11290
rect 14170 11230 14230 11250
rect 14290 11390 14350 11410
rect 14290 11350 14300 11390
rect 14340 11350 14350 11390
rect 14290 11290 14350 11350
rect 14290 11250 14300 11290
rect 14340 11250 14350 11290
rect 14290 11230 14350 11250
rect 14410 11390 14470 11410
rect 14410 11350 14420 11390
rect 14460 11350 14470 11390
rect 14410 11290 14470 11350
rect 14410 11250 14420 11290
rect 14460 11250 14470 11290
rect 14410 11230 14470 11250
rect 14530 11390 14590 11410
rect 14530 11350 14540 11390
rect 14580 11350 14590 11390
rect 14530 11290 14590 11350
rect 14530 11250 14540 11290
rect 14580 11250 14590 11290
rect 14530 11230 14590 11250
rect 14650 11390 14710 11410
rect 14650 11350 14660 11390
rect 14700 11350 14710 11390
rect 14650 11290 14710 11350
rect 14650 11250 14660 11290
rect 14700 11250 14710 11290
rect 14650 11230 14710 11250
rect 14770 11390 14830 11410
rect 14770 11350 14780 11390
rect 14820 11350 14830 11390
rect 14770 11290 14830 11350
rect 14770 11250 14780 11290
rect 14820 11250 14830 11290
rect 14770 11230 14830 11250
rect 14890 11390 14950 11410
rect 14890 11350 14900 11390
rect 14940 11350 14950 11390
rect 14890 11290 14950 11350
rect 14890 11250 14900 11290
rect 14940 11250 14950 11290
rect 14890 11230 14950 11250
rect 15010 11390 15070 11410
rect 15010 11350 15020 11390
rect 15060 11350 15070 11390
rect 15010 11290 15070 11350
rect 15010 11250 15020 11290
rect 15060 11250 15070 11290
rect 15010 11230 15070 11250
rect 15130 11390 15190 11410
rect 15130 11350 15140 11390
rect 15180 11350 15190 11390
rect 15130 11290 15190 11350
rect 15130 11250 15140 11290
rect 15180 11250 15190 11290
rect 15130 11230 15190 11250
rect 15250 11390 15310 11410
rect 15250 11350 15260 11390
rect 15300 11350 15310 11390
rect 15250 11290 15310 11350
rect 15250 11250 15260 11290
rect 15300 11250 15310 11290
rect 15250 11230 15310 11250
rect 15370 11390 15430 11410
rect 15370 11350 15380 11390
rect 15420 11350 15430 11390
rect 15370 11290 15430 11350
rect 15370 11250 15380 11290
rect 15420 11250 15430 11290
rect 15370 11230 15430 11250
rect 15490 11390 15550 11410
rect 15490 11350 15500 11390
rect 15540 11350 15550 11390
rect 15490 11290 15550 11350
rect 15490 11250 15500 11290
rect 15540 11250 15550 11290
rect 15490 11230 15550 11250
rect 15610 11390 15670 11410
rect 15610 11350 15620 11390
rect 15660 11350 15670 11390
rect 15610 11290 15670 11350
rect 15610 11250 15620 11290
rect 15660 11250 15670 11290
rect 15610 11230 15670 11250
rect 15730 11390 15790 11410
rect 15730 11350 15740 11390
rect 15780 11350 15790 11390
rect 15730 11290 15790 11350
rect 15730 11250 15740 11290
rect 15780 11250 15790 11290
rect 15730 11230 15790 11250
rect 15850 11390 15910 11410
rect 15850 11350 15860 11390
rect 15900 11350 15910 11390
rect 15850 11290 15910 11350
rect 15850 11250 15860 11290
rect 15900 11250 15910 11290
rect 15850 11230 15910 11250
rect 15970 11390 16110 11410
rect 15970 11350 15980 11390
rect 16020 11350 16060 11390
rect 16100 11350 16110 11390
rect 15970 11290 16110 11350
rect 15970 11250 15980 11290
rect 16020 11250 16060 11290
rect 16100 11250 16110 11290
rect 15970 11230 16110 11250
rect 10530 11170 10590 11190
rect 10530 11130 10540 11170
rect 10580 11130 10590 11170
rect 10530 11110 10590 11130
rect 12930 11170 12990 11190
rect 12930 11130 12940 11170
rect 12980 11130 12990 11170
rect 12930 11110 12990 11130
rect 13570 11170 13630 11190
rect 13570 11130 13580 11170
rect 13620 11130 13630 11170
rect 13570 11110 13630 11130
rect 15970 11170 16030 11190
rect 15970 11130 15980 11170
rect 16020 11130 16030 11170
rect 15970 11110 16030 11130
rect 11900 10350 11970 10370
rect 11900 10310 11910 10350
rect 11950 10310 11970 10350
rect 11900 10290 11970 10310
rect 12070 10350 12150 10370
rect 12070 10310 12090 10350
rect 12130 10310 12150 10350
rect 12070 10290 12150 10310
rect 12250 10350 12330 10370
rect 12250 10310 12270 10350
rect 12310 10310 12330 10350
rect 12250 10290 12330 10310
rect 12430 10350 12510 10370
rect 12430 10310 12450 10350
rect 12490 10310 12510 10350
rect 12430 10290 12510 10310
rect 12610 10350 12690 10370
rect 12610 10310 12630 10350
rect 12670 10310 12690 10350
rect 12610 10290 12690 10310
rect 12790 10350 12870 10370
rect 12790 10310 12810 10350
rect 12850 10310 12870 10350
rect 12790 10290 12870 10310
rect 12970 10350 13050 10370
rect 12970 10310 12990 10350
rect 13030 10310 13050 10350
rect 12970 10290 13050 10310
rect 13150 10350 13220 10370
rect 13150 10310 13170 10350
rect 13210 10310 13220 10350
rect 13150 10290 13220 10310
rect 13340 10350 13410 10370
rect 13340 10310 13350 10350
rect 13390 10310 13410 10350
rect 13340 10290 13410 10310
rect 13510 10350 13590 10370
rect 13510 10310 13530 10350
rect 13570 10310 13590 10350
rect 13510 10290 13590 10310
rect 13690 10350 13770 10370
rect 13690 10310 13710 10350
rect 13750 10310 13770 10350
rect 13690 10290 13770 10310
rect 13870 10350 13950 10370
rect 13870 10310 13890 10350
rect 13930 10310 13950 10350
rect 13870 10290 13950 10310
rect 14050 10350 14130 10370
rect 14050 10310 14070 10350
rect 14110 10310 14130 10350
rect 14050 10290 14130 10310
rect 14230 10350 14310 10370
rect 14230 10310 14250 10350
rect 14290 10310 14310 10350
rect 14230 10290 14310 10310
rect 14410 10350 14490 10370
rect 14410 10310 14430 10350
rect 14470 10310 14490 10350
rect 14410 10290 14490 10310
rect 14590 10350 14660 10370
rect 14590 10310 14610 10350
rect 14650 10310 14660 10350
rect 14590 10290 14660 10310
rect 11550 10230 11690 10250
rect 11550 10190 11560 10230
rect 11600 10190 11640 10230
rect 11680 10190 11690 10230
rect 11550 10130 11690 10190
rect 11550 10090 11560 10130
rect 11600 10090 11640 10130
rect 11680 10090 11690 10130
rect 11550 10030 11690 10090
rect 11550 9990 11560 10030
rect 11600 9990 11640 10030
rect 11680 9990 11690 10030
rect 11550 9930 11690 9990
rect 11550 9890 11560 9930
rect 11600 9890 11640 9930
rect 11680 9890 11690 9930
rect 11550 9830 11690 9890
rect 11550 9790 11560 9830
rect 11600 9790 11640 9830
rect 11680 9790 11690 9830
rect 11550 9730 11690 9790
rect 11550 9690 11560 9730
rect 11600 9690 11640 9730
rect 11680 9690 11690 9730
rect 11550 9670 11690 9690
rect 11810 10230 11870 10250
rect 11810 10190 11820 10230
rect 11860 10190 11870 10230
rect 11810 10130 11870 10190
rect 11810 10090 11820 10130
rect 11860 10090 11870 10130
rect 11810 10030 11870 10090
rect 11810 9990 11820 10030
rect 11860 9990 11870 10030
rect 11810 9930 11870 9990
rect 11810 9890 11820 9930
rect 11860 9890 11870 9930
rect 11810 9830 11870 9890
rect 11810 9790 11820 9830
rect 11860 9790 11870 9830
rect 11810 9730 11870 9790
rect 11810 9690 11820 9730
rect 11860 9690 11870 9730
rect 11810 9670 11870 9690
rect 11990 10230 12050 10250
rect 11990 10190 12000 10230
rect 12040 10190 12050 10230
rect 11990 10130 12050 10190
rect 11990 10090 12000 10130
rect 12040 10090 12050 10130
rect 11990 10030 12050 10090
rect 11990 9990 12000 10030
rect 12040 9990 12050 10030
rect 11990 9930 12050 9990
rect 11990 9890 12000 9930
rect 12040 9890 12050 9930
rect 11990 9830 12050 9890
rect 11990 9790 12000 9830
rect 12040 9790 12050 9830
rect 11990 9730 12050 9790
rect 11990 9690 12000 9730
rect 12040 9690 12050 9730
rect 11990 9670 12050 9690
rect 12170 10230 12230 10250
rect 12170 10190 12180 10230
rect 12220 10190 12230 10230
rect 12170 10130 12230 10190
rect 12170 10090 12180 10130
rect 12220 10090 12230 10130
rect 12170 10030 12230 10090
rect 12170 9990 12180 10030
rect 12220 9990 12230 10030
rect 12170 9930 12230 9990
rect 12170 9890 12180 9930
rect 12220 9890 12230 9930
rect 12170 9830 12230 9890
rect 12170 9790 12180 9830
rect 12220 9790 12230 9830
rect 12170 9730 12230 9790
rect 12170 9690 12180 9730
rect 12220 9690 12230 9730
rect 12170 9670 12230 9690
rect 12350 10230 12410 10250
rect 12350 10190 12360 10230
rect 12400 10190 12410 10230
rect 12350 10130 12410 10190
rect 12350 10090 12360 10130
rect 12400 10090 12410 10130
rect 12350 10030 12410 10090
rect 12350 9990 12360 10030
rect 12400 9990 12410 10030
rect 12350 9930 12410 9990
rect 12350 9890 12360 9930
rect 12400 9890 12410 9930
rect 12350 9830 12410 9890
rect 12350 9790 12360 9830
rect 12400 9790 12410 9830
rect 12350 9730 12410 9790
rect 12350 9690 12360 9730
rect 12400 9690 12410 9730
rect 12350 9670 12410 9690
rect 12530 10230 12590 10250
rect 12530 10190 12540 10230
rect 12580 10190 12590 10230
rect 12530 10130 12590 10190
rect 12530 10090 12540 10130
rect 12580 10090 12590 10130
rect 12530 10030 12590 10090
rect 12530 9990 12540 10030
rect 12580 9990 12590 10030
rect 12530 9930 12590 9990
rect 12530 9890 12540 9930
rect 12580 9890 12590 9930
rect 12530 9830 12590 9890
rect 12530 9790 12540 9830
rect 12580 9790 12590 9830
rect 12530 9730 12590 9790
rect 12530 9690 12540 9730
rect 12580 9690 12590 9730
rect 12530 9670 12590 9690
rect 12710 10230 12770 10250
rect 12710 10190 12720 10230
rect 12760 10190 12770 10230
rect 12710 10130 12770 10190
rect 12710 10090 12720 10130
rect 12760 10090 12770 10130
rect 12710 10030 12770 10090
rect 12710 9990 12720 10030
rect 12760 9990 12770 10030
rect 12710 9930 12770 9990
rect 12710 9890 12720 9930
rect 12760 9890 12770 9930
rect 12710 9830 12770 9890
rect 12710 9790 12720 9830
rect 12760 9790 12770 9830
rect 12710 9730 12770 9790
rect 12710 9690 12720 9730
rect 12760 9690 12770 9730
rect 12710 9670 12770 9690
rect 12890 10230 12950 10250
rect 12890 10190 12900 10230
rect 12940 10190 12950 10230
rect 12890 10130 12950 10190
rect 12890 10090 12900 10130
rect 12940 10090 12950 10130
rect 12890 10030 12950 10090
rect 12890 9990 12900 10030
rect 12940 9990 12950 10030
rect 12890 9930 12950 9990
rect 12890 9890 12900 9930
rect 12940 9890 12950 9930
rect 12890 9830 12950 9890
rect 12890 9790 12900 9830
rect 12940 9790 12950 9830
rect 12890 9730 12950 9790
rect 12890 9690 12900 9730
rect 12940 9690 12950 9730
rect 12890 9670 12950 9690
rect 13070 10230 13130 10250
rect 13070 10190 13080 10230
rect 13120 10190 13130 10230
rect 13070 10130 13130 10190
rect 13070 10090 13080 10130
rect 13120 10090 13130 10130
rect 13070 10030 13130 10090
rect 13070 9990 13080 10030
rect 13120 9990 13130 10030
rect 13070 9930 13130 9990
rect 13070 9890 13080 9930
rect 13120 9890 13130 9930
rect 13070 9830 13130 9890
rect 13070 9790 13080 9830
rect 13120 9790 13130 9830
rect 13070 9730 13130 9790
rect 13070 9690 13080 9730
rect 13120 9690 13130 9730
rect 13070 9670 13130 9690
rect 13250 10230 13310 10250
rect 13250 10190 13260 10230
rect 13300 10190 13310 10230
rect 13250 10130 13310 10190
rect 13250 10090 13260 10130
rect 13300 10090 13310 10130
rect 13250 10030 13310 10090
rect 13250 9990 13260 10030
rect 13300 9990 13310 10030
rect 13250 9930 13310 9990
rect 13250 9890 13260 9930
rect 13300 9890 13310 9930
rect 13250 9830 13310 9890
rect 13250 9790 13260 9830
rect 13300 9790 13310 9830
rect 13250 9730 13310 9790
rect 13250 9690 13260 9730
rect 13300 9690 13310 9730
rect 13250 9670 13310 9690
rect 13430 10230 13490 10250
rect 13430 10190 13440 10230
rect 13480 10190 13490 10230
rect 13430 10130 13490 10190
rect 13430 10090 13440 10130
rect 13480 10090 13490 10130
rect 13430 10030 13490 10090
rect 13430 9990 13440 10030
rect 13480 9990 13490 10030
rect 13430 9930 13490 9990
rect 13430 9890 13440 9930
rect 13480 9890 13490 9930
rect 13430 9830 13490 9890
rect 13430 9790 13440 9830
rect 13480 9790 13490 9830
rect 13430 9730 13490 9790
rect 13430 9690 13440 9730
rect 13480 9690 13490 9730
rect 13430 9670 13490 9690
rect 13610 10230 13670 10250
rect 13610 10190 13620 10230
rect 13660 10190 13670 10230
rect 13610 10130 13670 10190
rect 13610 10090 13620 10130
rect 13660 10090 13670 10130
rect 13610 10030 13670 10090
rect 13610 9990 13620 10030
rect 13660 9990 13670 10030
rect 13610 9930 13670 9990
rect 13610 9890 13620 9930
rect 13660 9890 13670 9930
rect 13610 9830 13670 9890
rect 13610 9790 13620 9830
rect 13660 9790 13670 9830
rect 13610 9730 13670 9790
rect 13610 9690 13620 9730
rect 13660 9690 13670 9730
rect 13610 9670 13670 9690
rect 13790 10230 13850 10250
rect 13790 10190 13800 10230
rect 13840 10190 13850 10230
rect 13790 10130 13850 10190
rect 13790 10090 13800 10130
rect 13840 10090 13850 10130
rect 13790 10030 13850 10090
rect 13790 9990 13800 10030
rect 13840 9990 13850 10030
rect 13790 9930 13850 9990
rect 13790 9890 13800 9930
rect 13840 9890 13850 9930
rect 13790 9830 13850 9890
rect 13790 9790 13800 9830
rect 13840 9790 13850 9830
rect 13790 9730 13850 9790
rect 13790 9690 13800 9730
rect 13840 9690 13850 9730
rect 13790 9670 13850 9690
rect 13970 10230 14030 10250
rect 13970 10190 13980 10230
rect 14020 10190 14030 10230
rect 13970 10130 14030 10190
rect 13970 10090 13980 10130
rect 14020 10090 14030 10130
rect 13970 10030 14030 10090
rect 13970 9990 13980 10030
rect 14020 9990 14030 10030
rect 13970 9930 14030 9990
rect 13970 9890 13980 9930
rect 14020 9890 14030 9930
rect 13970 9830 14030 9890
rect 13970 9790 13980 9830
rect 14020 9790 14030 9830
rect 13970 9730 14030 9790
rect 13970 9690 13980 9730
rect 14020 9690 14030 9730
rect 13970 9670 14030 9690
rect 14150 10230 14210 10250
rect 14150 10190 14160 10230
rect 14200 10190 14210 10230
rect 14150 10130 14210 10190
rect 14150 10090 14160 10130
rect 14200 10090 14210 10130
rect 14150 10030 14210 10090
rect 14150 9990 14160 10030
rect 14200 9990 14210 10030
rect 14150 9930 14210 9990
rect 14150 9890 14160 9930
rect 14200 9890 14210 9930
rect 14150 9830 14210 9890
rect 14150 9790 14160 9830
rect 14200 9790 14210 9830
rect 14150 9730 14210 9790
rect 14150 9690 14160 9730
rect 14200 9690 14210 9730
rect 14150 9670 14210 9690
rect 14330 10230 14390 10250
rect 14330 10190 14340 10230
rect 14380 10190 14390 10230
rect 14330 10130 14390 10190
rect 14330 10090 14340 10130
rect 14380 10090 14390 10130
rect 14330 10030 14390 10090
rect 14330 9990 14340 10030
rect 14380 9990 14390 10030
rect 14330 9930 14390 9990
rect 14330 9890 14340 9930
rect 14380 9890 14390 9930
rect 14330 9830 14390 9890
rect 14330 9790 14340 9830
rect 14380 9790 14390 9830
rect 14330 9730 14390 9790
rect 14330 9690 14340 9730
rect 14380 9690 14390 9730
rect 14330 9670 14390 9690
rect 14510 10230 14570 10250
rect 14510 10190 14520 10230
rect 14560 10190 14570 10230
rect 14510 10130 14570 10190
rect 14510 10090 14520 10130
rect 14560 10090 14570 10130
rect 14510 10030 14570 10090
rect 14510 9990 14520 10030
rect 14560 9990 14570 10030
rect 14510 9930 14570 9990
rect 14510 9890 14520 9930
rect 14560 9890 14570 9930
rect 14510 9830 14570 9890
rect 14510 9790 14520 9830
rect 14560 9790 14570 9830
rect 14510 9730 14570 9790
rect 14510 9690 14520 9730
rect 14560 9690 14570 9730
rect 14510 9670 14570 9690
rect 14690 10230 14750 10250
rect 14690 10190 14700 10230
rect 14740 10190 14750 10230
rect 14690 10130 14750 10190
rect 14690 10090 14700 10130
rect 14740 10090 14750 10130
rect 14690 10030 14750 10090
rect 14690 9990 14700 10030
rect 14740 9990 14750 10030
rect 14690 9930 14750 9990
rect 14690 9890 14700 9930
rect 14740 9890 14750 9930
rect 14690 9830 14750 9890
rect 14690 9790 14700 9830
rect 14740 9790 14750 9830
rect 14690 9730 14750 9790
rect 14690 9690 14700 9730
rect 14740 9690 14750 9730
rect 14690 9670 14750 9690
rect 14870 10230 15010 10250
rect 14870 10190 14880 10230
rect 14920 10190 14960 10230
rect 15000 10190 15010 10230
rect 14870 10130 15010 10190
rect 14870 10090 14880 10130
rect 14920 10090 14960 10130
rect 15000 10090 15010 10130
rect 15590 10150 15670 10170
rect 15590 10110 15610 10150
rect 15650 10110 15670 10150
rect 15590 10090 15670 10110
rect 15710 10150 15790 10170
rect 15710 10110 15730 10150
rect 15770 10110 15790 10150
rect 15710 10090 15790 10110
rect 15830 10150 15910 10170
rect 15830 10110 15850 10150
rect 15890 10110 15910 10150
rect 15830 10090 15910 10110
rect 14870 10030 15010 10090
rect 14870 9990 14880 10030
rect 14920 9990 14960 10030
rect 15000 9990 15010 10030
rect 14870 9930 15010 9990
rect 14870 9890 14880 9930
rect 14920 9890 14960 9930
rect 15000 9890 15010 9930
rect 14870 9830 15010 9890
rect 15410 10030 15560 10050
rect 15410 9990 15420 10030
rect 15460 9990 15510 10030
rect 15550 9990 15560 10030
rect 15410 9930 15560 9990
rect 15410 9890 15420 9930
rect 15460 9890 15510 9930
rect 15550 9890 15560 9930
rect 15410 9870 15560 9890
rect 15610 10030 15670 10050
rect 15610 9990 15620 10030
rect 15660 9990 15670 10030
rect 15610 9930 15670 9990
rect 15610 9890 15620 9930
rect 15660 9890 15670 9930
rect 15610 9870 15670 9890
rect 15720 10030 15780 10050
rect 15720 9990 15730 10030
rect 15770 9990 15780 10030
rect 15720 9930 15780 9990
rect 15720 9890 15730 9930
rect 15770 9890 15780 9930
rect 15720 9870 15780 9890
rect 15830 10030 15890 10050
rect 15830 9990 15840 10030
rect 15880 9990 15890 10030
rect 15830 9930 15890 9990
rect 15830 9890 15840 9930
rect 15880 9890 15890 9930
rect 15830 9870 15890 9890
rect 15940 10030 16080 10050
rect 15940 9990 15950 10030
rect 15990 9990 16030 10030
rect 16070 9990 16080 10030
rect 15940 9930 16080 9990
rect 15940 9890 15950 9930
rect 15990 9890 16030 9930
rect 16070 9890 16080 9930
rect 15940 9870 16080 9890
rect 14870 9790 14880 9830
rect 14920 9790 14960 9830
rect 15000 9790 15010 9830
rect 14870 9730 15010 9790
rect 15490 9810 15570 9830
rect 15490 9770 15510 9810
rect 15550 9770 15570 9810
rect 15490 9750 15570 9770
rect 15710 9810 15790 9830
rect 15710 9770 15730 9810
rect 15770 9770 15790 9810
rect 15710 9750 15790 9770
rect 15940 9810 16000 9830
rect 15940 9770 15950 9810
rect 15990 9770 16000 9810
rect 15940 9750 16000 9770
rect 14870 9690 14880 9730
rect 14920 9690 14960 9730
rect 15000 9690 15010 9730
rect 14870 9670 15010 9690
rect 11640 9630 11680 9670
rect 12000 9630 12040 9670
rect 12360 9630 12400 9670
rect 12720 9630 12760 9670
rect 13080 9630 13120 9670
rect 13440 9630 13480 9670
rect 13800 9630 13840 9670
rect 14160 9630 14200 9670
rect 14520 9630 14560 9670
rect 14880 9630 14920 9670
rect 11620 9610 11700 9630
rect 11620 9570 11640 9610
rect 11680 9570 11700 9610
rect 11620 9550 11700 9570
rect 11980 9610 12060 9630
rect 11980 9570 12000 9610
rect 12040 9570 12060 9610
rect 11980 9550 12060 9570
rect 12340 9610 12420 9630
rect 12340 9570 12360 9610
rect 12400 9570 12420 9610
rect 12340 9550 12420 9570
rect 12700 9610 12780 9630
rect 12700 9570 12720 9610
rect 12760 9570 12780 9610
rect 12700 9550 12780 9570
rect 13060 9610 13140 9630
rect 13060 9570 13080 9610
rect 13120 9570 13140 9610
rect 13060 9550 13140 9570
rect 13420 9610 13500 9630
rect 13420 9570 13440 9610
rect 13480 9570 13500 9610
rect 13420 9550 13500 9570
rect 13780 9610 13860 9630
rect 13780 9570 13800 9610
rect 13840 9570 13860 9610
rect 13780 9550 13860 9570
rect 14140 9610 14220 9630
rect 14140 9570 14160 9610
rect 14200 9570 14220 9610
rect 14140 9550 14220 9570
rect 14500 9610 14580 9630
rect 14500 9570 14520 9610
rect 14560 9570 14580 9610
rect 14500 9550 14580 9570
rect 14860 9610 14940 9630
rect 14860 9570 14880 9610
rect 14920 9570 14940 9610
rect 14860 9550 14940 9570
rect 11806 9342 11864 9360
rect 11806 9308 11818 9342
rect 11852 9308 11864 9342
rect 11806 9290 11864 9308
rect 11916 9342 11974 9360
rect 11916 9308 11928 9342
rect 11962 9308 11974 9342
rect 11916 9290 11974 9308
rect 12026 9342 12084 9360
rect 12026 9308 12038 9342
rect 12072 9308 12084 9342
rect 12026 9290 12084 9308
rect 12136 9342 12194 9360
rect 12136 9308 12148 9342
rect 12182 9308 12194 9342
rect 12136 9290 12194 9308
rect 12246 9342 12304 9360
rect 12246 9308 12258 9342
rect 12292 9308 12304 9342
rect 12246 9290 12304 9308
rect 12356 9342 12414 9360
rect 12356 9308 12368 9342
rect 12402 9308 12414 9342
rect 12356 9290 12414 9308
rect 12466 9342 12524 9360
rect 12466 9308 12478 9342
rect 12512 9308 12524 9342
rect 12466 9290 12524 9308
rect 12576 9342 12634 9360
rect 12576 9308 12588 9342
rect 12622 9308 12634 9342
rect 12576 9290 12634 9308
rect 12686 9342 12744 9360
rect 12686 9308 12698 9342
rect 12732 9308 12744 9342
rect 12686 9290 12744 9308
rect 12796 9342 12854 9360
rect 12796 9308 12808 9342
rect 12842 9308 12854 9342
rect 12796 9290 12854 9308
rect 13706 9342 13764 9360
rect 13706 9308 13718 9342
rect 13752 9308 13764 9342
rect 13706 9290 13764 9308
rect 13816 9342 13874 9360
rect 13816 9308 13828 9342
rect 13862 9308 13874 9342
rect 13816 9290 13874 9308
rect 13926 9342 13984 9360
rect 13926 9308 13938 9342
rect 13972 9308 13984 9342
rect 13926 9290 13984 9308
rect 14036 9342 14094 9360
rect 14036 9308 14048 9342
rect 14082 9308 14094 9342
rect 14036 9290 14094 9308
rect 14146 9342 14204 9360
rect 14146 9308 14158 9342
rect 14192 9308 14204 9342
rect 14146 9290 14204 9308
rect 14256 9342 14314 9360
rect 14256 9308 14268 9342
rect 14302 9308 14314 9342
rect 14256 9290 14314 9308
rect 14366 9342 14424 9360
rect 14366 9308 14378 9342
rect 14412 9308 14424 9342
rect 14366 9290 14424 9308
rect 14476 9342 14534 9360
rect 14476 9308 14488 9342
rect 14522 9308 14534 9342
rect 14476 9290 14534 9308
rect 14586 9342 14644 9360
rect 14586 9308 14598 9342
rect 14632 9308 14644 9342
rect 14586 9290 14644 9308
rect 14696 9342 14754 9360
rect 14696 9308 14708 9342
rect 14742 9308 14754 9342
rect 14696 9290 14754 9308
rect 11560 9230 11700 9250
rect 11560 9190 11570 9230
rect 11610 9190 11650 9230
rect 11690 9190 11700 9230
rect 11560 9130 11700 9190
rect 11560 9090 11570 9130
rect 11610 9090 11650 9130
rect 11690 9090 11700 9130
rect 11560 9070 11700 9090
rect 11750 9230 11810 9250
rect 11750 9190 11760 9230
rect 11800 9190 11810 9230
rect 11750 9130 11810 9190
rect 11750 9090 11760 9130
rect 11800 9090 11810 9130
rect 11750 9070 11810 9090
rect 11860 9230 11920 9250
rect 11860 9190 11870 9230
rect 11910 9190 11920 9230
rect 11860 9130 11920 9190
rect 11860 9090 11870 9130
rect 11910 9090 11920 9130
rect 11860 9070 11920 9090
rect 11970 9230 12030 9250
rect 11970 9190 11980 9230
rect 12020 9190 12030 9230
rect 11970 9130 12030 9190
rect 11970 9090 11980 9130
rect 12020 9090 12030 9130
rect 11970 9070 12030 9090
rect 12080 9230 12140 9250
rect 12080 9190 12090 9230
rect 12130 9190 12140 9230
rect 12080 9130 12140 9190
rect 12080 9090 12090 9130
rect 12130 9090 12140 9130
rect 12080 9070 12140 9090
rect 12190 9230 12250 9250
rect 12190 9190 12200 9230
rect 12240 9190 12250 9230
rect 12190 9130 12250 9190
rect 12190 9090 12200 9130
rect 12240 9090 12250 9130
rect 12190 9070 12250 9090
rect 12300 9230 12360 9250
rect 12300 9190 12310 9230
rect 12350 9190 12360 9230
rect 12300 9130 12360 9190
rect 12300 9090 12310 9130
rect 12350 9090 12360 9130
rect 12300 9070 12360 9090
rect 12410 9230 12470 9250
rect 12410 9190 12420 9230
rect 12460 9190 12470 9230
rect 12410 9130 12470 9190
rect 12410 9090 12420 9130
rect 12460 9090 12470 9130
rect 12410 9070 12470 9090
rect 12520 9230 12580 9250
rect 12520 9190 12530 9230
rect 12570 9190 12580 9230
rect 12520 9130 12580 9190
rect 12520 9090 12530 9130
rect 12570 9090 12580 9130
rect 12520 9070 12580 9090
rect 12630 9230 12690 9250
rect 12630 9190 12640 9230
rect 12680 9190 12690 9230
rect 12630 9130 12690 9190
rect 12630 9090 12640 9130
rect 12680 9090 12690 9130
rect 12630 9070 12690 9090
rect 12740 9230 12800 9250
rect 12740 9190 12750 9230
rect 12790 9190 12800 9230
rect 12740 9130 12800 9190
rect 12740 9090 12750 9130
rect 12790 9090 12800 9130
rect 12740 9070 12800 9090
rect 12850 9230 12910 9250
rect 12850 9190 12860 9230
rect 12900 9190 12910 9230
rect 12850 9130 12910 9190
rect 12850 9090 12860 9130
rect 12900 9090 12910 9130
rect 12850 9070 12910 9090
rect 12960 9230 13100 9250
rect 12960 9190 12970 9230
rect 13010 9190 13050 9230
rect 13090 9190 13100 9230
rect 12960 9130 13100 9190
rect 12960 9090 12970 9130
rect 13010 9090 13050 9130
rect 13090 9090 13100 9130
rect 12960 9070 13100 9090
rect 13460 9230 13600 9250
rect 13460 9190 13470 9230
rect 13510 9190 13550 9230
rect 13590 9190 13600 9230
rect 13460 9130 13600 9190
rect 13460 9090 13470 9130
rect 13510 9090 13550 9130
rect 13590 9090 13600 9130
rect 13460 9070 13600 9090
rect 13650 9230 13710 9250
rect 13650 9190 13660 9230
rect 13700 9190 13710 9230
rect 13650 9130 13710 9190
rect 13650 9090 13660 9130
rect 13700 9090 13710 9130
rect 13650 9070 13710 9090
rect 13760 9230 13820 9250
rect 13760 9190 13770 9230
rect 13810 9190 13820 9230
rect 13760 9130 13820 9190
rect 13760 9090 13770 9130
rect 13810 9090 13820 9130
rect 13760 9070 13820 9090
rect 13870 9230 13930 9250
rect 13870 9190 13880 9230
rect 13920 9190 13930 9230
rect 13870 9130 13930 9190
rect 13870 9090 13880 9130
rect 13920 9090 13930 9130
rect 13870 9070 13930 9090
rect 13980 9230 14040 9250
rect 13980 9190 13990 9230
rect 14030 9190 14040 9230
rect 13980 9130 14040 9190
rect 13980 9090 13990 9130
rect 14030 9090 14040 9130
rect 13980 9070 14040 9090
rect 14090 9230 14150 9250
rect 14090 9190 14100 9230
rect 14140 9190 14150 9230
rect 14090 9130 14150 9190
rect 14090 9090 14100 9130
rect 14140 9090 14150 9130
rect 14090 9070 14150 9090
rect 14200 9230 14260 9250
rect 14200 9190 14210 9230
rect 14250 9190 14260 9230
rect 14200 9130 14260 9190
rect 14200 9090 14210 9130
rect 14250 9090 14260 9130
rect 14200 9070 14260 9090
rect 14310 9230 14370 9250
rect 14310 9190 14320 9230
rect 14360 9190 14370 9230
rect 14310 9130 14370 9190
rect 14310 9090 14320 9130
rect 14360 9090 14370 9130
rect 14310 9070 14370 9090
rect 14420 9230 14480 9250
rect 14420 9190 14430 9230
rect 14470 9190 14480 9230
rect 14420 9130 14480 9190
rect 14420 9090 14430 9130
rect 14470 9090 14480 9130
rect 14420 9070 14480 9090
rect 14530 9230 14590 9250
rect 14530 9190 14540 9230
rect 14580 9190 14590 9230
rect 14530 9130 14590 9190
rect 14530 9090 14540 9130
rect 14580 9090 14590 9130
rect 14530 9070 14590 9090
rect 14640 9230 14700 9250
rect 14640 9190 14650 9230
rect 14690 9190 14700 9230
rect 14640 9130 14700 9190
rect 14640 9090 14650 9130
rect 14690 9090 14700 9130
rect 14640 9070 14700 9090
rect 14750 9230 14810 9250
rect 14750 9190 14760 9230
rect 14800 9190 14810 9230
rect 14750 9130 14810 9190
rect 14750 9090 14760 9130
rect 14800 9090 14810 9130
rect 14750 9070 14810 9090
rect 14860 9230 15000 9250
rect 14860 9190 14870 9230
rect 14910 9190 14950 9230
rect 14990 9190 15000 9230
rect 14860 9130 15000 9190
rect 14860 9090 14870 9130
rect 14910 9090 14950 9130
rect 14990 9090 15000 9130
rect 14860 9070 15000 9090
rect 11630 9010 11710 9030
rect 11630 8970 11650 9010
rect 11690 8970 11710 9010
rect 11630 8950 11710 8970
rect 12950 9010 13030 9030
rect 12950 8970 12970 9010
rect 13010 8970 13030 9010
rect 12950 8950 13030 8970
rect 13530 9010 13610 9030
rect 13530 8970 13550 9010
rect 13590 8970 13610 9010
rect 13530 8950 13610 8970
rect 14850 9010 14930 9030
rect 14850 8970 14870 9010
rect 14910 8970 14930 9010
rect 14850 8950 14930 8970
<< viali >>
rect 13260 19030 13300 19070
rect 13260 18950 13300 18990
rect 13260 18870 13300 18910
rect 9590 18595 9630 18600
rect 10700 18597 10740 18610
rect 8810 18589 8850 18590
rect 8810 18555 8850 18589
rect 8810 18550 8850 18555
rect 8776 18035 8882 18432
rect 8776 16650 8882 17047
rect 9590 18561 9630 18595
rect 9590 18560 9630 18561
rect 9590 18041 9628 18438
rect 9590 15080 9628 15477
rect 10700 18570 10740 18597
rect 10700 18050 10740 18440
rect 10370 16310 10410 16700
rect 11660 18392 11666 18414
rect 11666 18392 11694 18414
rect 11660 18380 11694 18392
rect 11760 18380 11794 18414
rect 11860 18380 11894 18414
rect 11960 18392 11992 18414
rect 11992 18392 11994 18414
rect 12060 18392 12082 18414
rect 12082 18392 12094 18414
rect 12160 18392 12172 18414
rect 12172 18392 12194 18414
rect 11960 18380 11994 18392
rect 12060 18380 12094 18392
rect 12160 18380 12194 18392
rect 11660 18302 11666 18314
rect 11666 18302 11694 18314
rect 11660 18280 11694 18302
rect 11760 18280 11794 18314
rect 11860 18280 11894 18314
rect 11960 18302 11992 18314
rect 11992 18302 11994 18314
rect 12060 18302 12082 18314
rect 12082 18302 12094 18314
rect 12160 18302 12172 18314
rect 12172 18302 12194 18314
rect 11960 18280 11994 18302
rect 12060 18280 12094 18302
rect 12160 18280 12194 18302
rect 11660 18212 11666 18214
rect 11666 18212 11694 18214
rect 11660 18180 11694 18212
rect 11760 18180 11794 18214
rect 11860 18180 11894 18214
rect 11960 18212 11992 18214
rect 11992 18212 11994 18214
rect 12060 18212 12082 18214
rect 12082 18212 12094 18214
rect 12160 18212 12172 18214
rect 12172 18212 12194 18214
rect 11960 18180 11994 18212
rect 12060 18180 12094 18212
rect 12160 18180 12194 18212
rect 11660 18080 11694 18114
rect 11760 18080 11794 18114
rect 11860 18080 11894 18114
rect 11960 18080 11994 18114
rect 12060 18080 12094 18114
rect 12160 18080 12194 18114
rect 11660 17980 11694 18014
rect 11760 17980 11794 18014
rect 11860 17980 11894 18014
rect 11960 17980 11994 18014
rect 12060 17980 12094 18014
rect 12160 17980 12194 18014
rect 11660 17886 11694 17914
rect 11660 17880 11666 17886
rect 11666 17880 11694 17886
rect 11760 17880 11794 17914
rect 11860 17880 11894 17914
rect 11960 17886 11994 17914
rect 12060 17886 12094 17914
rect 12160 17886 12194 17914
rect 11960 17880 11992 17886
rect 11992 17880 11994 17886
rect 12060 17880 12082 17886
rect 12082 17880 12094 17886
rect 12160 17880 12172 17886
rect 12172 17880 12194 17886
rect 13020 18392 13026 18414
rect 13026 18392 13054 18414
rect 13020 18380 13054 18392
rect 13120 18380 13154 18414
rect 13220 18380 13254 18414
rect 13320 18392 13352 18414
rect 13352 18392 13354 18414
rect 13420 18392 13442 18414
rect 13442 18392 13454 18414
rect 13520 18392 13532 18414
rect 13532 18392 13554 18414
rect 13320 18380 13354 18392
rect 13420 18380 13454 18392
rect 13520 18380 13554 18392
rect 13020 18302 13026 18314
rect 13026 18302 13054 18314
rect 13020 18280 13054 18302
rect 13120 18280 13154 18314
rect 13220 18280 13254 18314
rect 13320 18302 13352 18314
rect 13352 18302 13354 18314
rect 13420 18302 13442 18314
rect 13442 18302 13454 18314
rect 13520 18302 13532 18314
rect 13532 18302 13554 18314
rect 13320 18280 13354 18302
rect 13420 18280 13454 18302
rect 13520 18280 13554 18302
rect 13020 18212 13026 18214
rect 13026 18212 13054 18214
rect 13020 18180 13054 18212
rect 13120 18180 13154 18214
rect 13220 18180 13254 18214
rect 13320 18212 13352 18214
rect 13352 18212 13354 18214
rect 13420 18212 13442 18214
rect 13442 18212 13454 18214
rect 13520 18212 13532 18214
rect 13532 18212 13554 18214
rect 13320 18180 13354 18212
rect 13420 18180 13454 18212
rect 13520 18180 13554 18212
rect 13020 18080 13054 18114
rect 13120 18080 13154 18114
rect 13220 18080 13254 18114
rect 13320 18080 13354 18114
rect 13420 18080 13454 18114
rect 13520 18080 13554 18114
rect 13020 17980 13054 18014
rect 13120 17980 13154 18014
rect 13220 17980 13254 18014
rect 13320 17980 13354 18014
rect 13420 17980 13454 18014
rect 13520 17980 13554 18014
rect 13020 17886 13054 17914
rect 13020 17880 13026 17886
rect 13026 17880 13054 17886
rect 13120 17880 13154 17914
rect 13220 17880 13254 17914
rect 13320 17886 13354 17914
rect 13420 17886 13454 17914
rect 13520 17886 13554 17914
rect 13320 17880 13352 17886
rect 13352 17880 13354 17886
rect 13420 17880 13442 17886
rect 13442 17880 13454 17886
rect 13520 17880 13532 17886
rect 13532 17880 13554 17886
rect 14380 18392 14386 18414
rect 14386 18392 14414 18414
rect 14380 18380 14414 18392
rect 14480 18380 14514 18414
rect 14580 18380 14614 18414
rect 14680 18392 14712 18414
rect 14712 18392 14714 18414
rect 14780 18392 14802 18414
rect 14802 18392 14814 18414
rect 14880 18392 14892 18414
rect 14892 18392 14914 18414
rect 14680 18380 14714 18392
rect 14780 18380 14814 18392
rect 14880 18380 14914 18392
rect 14380 18302 14386 18314
rect 14386 18302 14414 18314
rect 14380 18280 14414 18302
rect 14480 18280 14514 18314
rect 14580 18280 14614 18314
rect 14680 18302 14712 18314
rect 14712 18302 14714 18314
rect 14780 18302 14802 18314
rect 14802 18302 14814 18314
rect 14880 18302 14892 18314
rect 14892 18302 14914 18314
rect 14680 18280 14714 18302
rect 14780 18280 14814 18302
rect 14880 18280 14914 18302
rect 14380 18212 14386 18214
rect 14386 18212 14414 18214
rect 14380 18180 14414 18212
rect 14480 18180 14514 18214
rect 14580 18180 14614 18214
rect 14680 18212 14712 18214
rect 14712 18212 14714 18214
rect 14780 18212 14802 18214
rect 14802 18212 14814 18214
rect 14880 18212 14892 18214
rect 14892 18212 14914 18214
rect 14680 18180 14714 18212
rect 14780 18180 14814 18212
rect 14880 18180 14914 18212
rect 14380 18080 14414 18114
rect 14480 18080 14514 18114
rect 14580 18080 14614 18114
rect 14680 18080 14714 18114
rect 14780 18080 14814 18114
rect 14880 18080 14914 18114
rect 14380 17980 14414 18014
rect 14480 17980 14514 18014
rect 14580 17980 14614 18014
rect 14680 17980 14714 18014
rect 14780 17980 14814 18014
rect 14880 17980 14914 18014
rect 14380 17886 14414 17914
rect 14380 17880 14386 17886
rect 14386 17880 14414 17886
rect 14480 17880 14514 17914
rect 14580 17880 14614 17914
rect 14680 17886 14714 17914
rect 14780 17886 14814 17914
rect 14880 17886 14914 17914
rect 14680 17880 14712 17886
rect 14712 17880 14714 17886
rect 14780 17880 14802 17886
rect 14802 17880 14814 17886
rect 14880 17880 14892 17886
rect 14892 17880 14914 17886
rect 15690 18597 15730 18610
rect 15690 18570 15730 18597
rect 16800 18595 16840 18610
rect 11660 17032 11666 17054
rect 11666 17032 11694 17054
rect 11660 17020 11694 17032
rect 11760 17020 11794 17054
rect 11860 17020 11894 17054
rect 11960 17032 11992 17054
rect 11992 17032 11994 17054
rect 12060 17032 12082 17054
rect 12082 17032 12094 17054
rect 12160 17032 12172 17054
rect 12172 17032 12194 17054
rect 11960 17020 11994 17032
rect 12060 17020 12094 17032
rect 12160 17020 12194 17032
rect 11660 16942 11666 16954
rect 11666 16942 11694 16954
rect 11660 16920 11694 16942
rect 11760 16920 11794 16954
rect 11860 16920 11894 16954
rect 11960 16942 11992 16954
rect 11992 16942 11994 16954
rect 12060 16942 12082 16954
rect 12082 16942 12094 16954
rect 12160 16942 12172 16954
rect 12172 16942 12194 16954
rect 11960 16920 11994 16942
rect 12060 16920 12094 16942
rect 12160 16920 12194 16942
rect 11660 16852 11666 16854
rect 11666 16852 11694 16854
rect 11660 16820 11694 16852
rect 11760 16820 11794 16854
rect 11860 16820 11894 16854
rect 11960 16852 11992 16854
rect 11992 16852 11994 16854
rect 12060 16852 12082 16854
rect 12082 16852 12094 16854
rect 12160 16852 12172 16854
rect 12172 16852 12194 16854
rect 11960 16820 11994 16852
rect 12060 16820 12094 16852
rect 12160 16820 12194 16852
rect 11660 16720 11694 16754
rect 11760 16720 11794 16754
rect 11860 16720 11894 16754
rect 11960 16720 11994 16754
rect 12060 16720 12094 16754
rect 12160 16720 12194 16754
rect 11660 16620 11694 16654
rect 11760 16620 11794 16654
rect 11860 16620 11894 16654
rect 11960 16620 11994 16654
rect 12060 16620 12094 16654
rect 12160 16620 12194 16654
rect 11660 16526 11694 16554
rect 11660 16520 11666 16526
rect 11666 16520 11694 16526
rect 11760 16520 11794 16554
rect 11860 16520 11894 16554
rect 11960 16526 11994 16554
rect 12060 16526 12094 16554
rect 12160 16526 12194 16554
rect 11960 16520 11992 16526
rect 11992 16520 11994 16526
rect 12060 16520 12082 16526
rect 12082 16520 12094 16526
rect 12160 16520 12172 16526
rect 12172 16520 12194 16526
rect 13020 17032 13026 17054
rect 13026 17032 13054 17054
rect 13020 17020 13054 17032
rect 13120 17020 13154 17054
rect 13220 17020 13254 17054
rect 13320 17032 13352 17054
rect 13352 17032 13354 17054
rect 13420 17032 13442 17054
rect 13442 17032 13454 17054
rect 13520 17032 13532 17054
rect 13532 17032 13554 17054
rect 13320 17020 13354 17032
rect 13420 17020 13454 17032
rect 13520 17020 13554 17032
rect 13020 16942 13026 16954
rect 13026 16942 13054 16954
rect 13020 16920 13054 16942
rect 13120 16920 13154 16954
rect 13220 16920 13254 16954
rect 13320 16942 13352 16954
rect 13352 16942 13354 16954
rect 13420 16942 13442 16954
rect 13442 16942 13454 16954
rect 13520 16942 13532 16954
rect 13532 16942 13554 16954
rect 13320 16920 13354 16942
rect 13420 16920 13454 16942
rect 13520 16920 13554 16942
rect 13020 16852 13026 16854
rect 13026 16852 13054 16854
rect 13020 16820 13054 16852
rect 13120 16820 13154 16854
rect 13220 16820 13254 16854
rect 13320 16852 13352 16854
rect 13352 16852 13354 16854
rect 13420 16852 13442 16854
rect 13442 16852 13454 16854
rect 13520 16852 13532 16854
rect 13532 16852 13554 16854
rect 13320 16820 13354 16852
rect 13420 16820 13454 16852
rect 13520 16820 13554 16852
rect 13020 16720 13054 16754
rect 13120 16720 13154 16754
rect 13220 16720 13254 16754
rect 13320 16720 13354 16754
rect 13420 16720 13454 16754
rect 13520 16720 13554 16754
rect 13020 16620 13054 16654
rect 13120 16620 13154 16654
rect 13220 16620 13254 16654
rect 13320 16620 13354 16654
rect 13420 16620 13454 16654
rect 13520 16620 13554 16654
rect 13020 16526 13054 16554
rect 13020 16520 13026 16526
rect 13026 16520 13054 16526
rect 13120 16520 13154 16554
rect 13220 16520 13254 16554
rect 13320 16526 13354 16554
rect 13420 16526 13454 16554
rect 13520 16526 13554 16554
rect 13320 16520 13352 16526
rect 13352 16520 13354 16526
rect 13420 16520 13442 16526
rect 13442 16520 13454 16526
rect 13520 16520 13532 16526
rect 13532 16520 13554 16526
rect 14380 17032 14386 17054
rect 14386 17032 14414 17054
rect 14380 17020 14414 17032
rect 14480 17020 14514 17054
rect 14580 17020 14614 17054
rect 14680 17032 14712 17054
rect 14712 17032 14714 17054
rect 14780 17032 14802 17054
rect 14802 17032 14814 17054
rect 14880 17032 14892 17054
rect 14892 17032 14914 17054
rect 14680 17020 14714 17032
rect 14780 17020 14814 17032
rect 14880 17020 14914 17032
rect 14380 16942 14386 16954
rect 14386 16942 14414 16954
rect 14380 16920 14414 16942
rect 14480 16920 14514 16954
rect 14580 16920 14614 16954
rect 14680 16942 14712 16954
rect 14712 16942 14714 16954
rect 14780 16942 14802 16954
rect 14802 16942 14814 16954
rect 14880 16942 14892 16954
rect 14892 16942 14914 16954
rect 14680 16920 14714 16942
rect 14780 16920 14814 16942
rect 14880 16920 14914 16942
rect 14380 16852 14386 16854
rect 14386 16852 14414 16854
rect 14380 16820 14414 16852
rect 14480 16820 14514 16854
rect 14580 16820 14614 16854
rect 14680 16852 14712 16854
rect 14712 16852 14714 16854
rect 14780 16852 14802 16854
rect 14802 16852 14814 16854
rect 14880 16852 14892 16854
rect 14892 16852 14914 16854
rect 14680 16820 14714 16852
rect 14780 16820 14814 16852
rect 14880 16820 14914 16852
rect 14380 16720 14414 16754
rect 14480 16720 14514 16754
rect 14580 16720 14614 16754
rect 14680 16720 14714 16754
rect 14780 16720 14814 16754
rect 14880 16720 14914 16754
rect 14380 16620 14414 16654
rect 14480 16620 14514 16654
rect 14580 16620 14614 16654
rect 14680 16620 14714 16654
rect 14780 16620 14814 16654
rect 14880 16620 14914 16654
rect 14380 16526 14414 16554
rect 14380 16520 14386 16526
rect 14386 16520 14414 16526
rect 14480 16520 14514 16554
rect 14580 16520 14614 16554
rect 14680 16526 14714 16554
rect 14780 16526 14814 16554
rect 14880 16526 14914 16554
rect 14680 16520 14712 16526
rect 14712 16520 14714 16526
rect 14780 16520 14802 16526
rect 14802 16520 14814 16526
rect 14880 16520 14892 16526
rect 14892 16520 14914 16526
rect 15690 18050 15730 18440
rect 16020 16310 16060 16700
rect 16800 18570 16840 18595
rect 17590 18589 17630 18590
rect 11660 15672 11666 15694
rect 11666 15672 11694 15694
rect 11660 15660 11694 15672
rect 11760 15660 11794 15694
rect 11860 15660 11894 15694
rect 11960 15672 11992 15694
rect 11992 15672 11994 15694
rect 12060 15672 12082 15694
rect 12082 15672 12094 15694
rect 12160 15672 12172 15694
rect 12172 15672 12194 15694
rect 11960 15660 11994 15672
rect 12060 15660 12094 15672
rect 12160 15660 12194 15672
rect 11660 15582 11666 15594
rect 11666 15582 11694 15594
rect 11660 15560 11694 15582
rect 11760 15560 11794 15594
rect 11860 15560 11894 15594
rect 11960 15582 11992 15594
rect 11992 15582 11994 15594
rect 12060 15582 12082 15594
rect 12082 15582 12094 15594
rect 12160 15582 12172 15594
rect 12172 15582 12194 15594
rect 11960 15560 11994 15582
rect 12060 15560 12094 15582
rect 12160 15560 12194 15582
rect 11660 15492 11666 15494
rect 11666 15492 11694 15494
rect 11660 15460 11694 15492
rect 11760 15460 11794 15494
rect 11860 15460 11894 15494
rect 11960 15492 11992 15494
rect 11992 15492 11994 15494
rect 12060 15492 12082 15494
rect 12082 15492 12094 15494
rect 12160 15492 12172 15494
rect 12172 15492 12194 15494
rect 11960 15460 11994 15492
rect 12060 15460 12094 15492
rect 12160 15460 12194 15492
rect 11660 15360 11694 15394
rect 11760 15360 11794 15394
rect 11860 15360 11894 15394
rect 11960 15360 11994 15394
rect 12060 15360 12094 15394
rect 12160 15360 12194 15394
rect 11660 15260 11694 15294
rect 11760 15260 11794 15294
rect 11860 15260 11894 15294
rect 11960 15260 11994 15294
rect 12060 15260 12094 15294
rect 12160 15260 12194 15294
rect 11660 15166 11694 15194
rect 11660 15160 11666 15166
rect 11666 15160 11694 15166
rect 11760 15160 11794 15194
rect 11860 15160 11894 15194
rect 11960 15166 11994 15194
rect 12060 15166 12094 15194
rect 12160 15166 12194 15194
rect 11960 15160 11992 15166
rect 11992 15160 11994 15166
rect 12060 15160 12082 15166
rect 12082 15160 12094 15166
rect 12160 15160 12172 15166
rect 12172 15160 12194 15166
rect 13020 15672 13026 15694
rect 13026 15672 13054 15694
rect 13020 15660 13054 15672
rect 13120 15660 13154 15694
rect 13220 15660 13254 15694
rect 13320 15672 13352 15694
rect 13352 15672 13354 15694
rect 13420 15672 13442 15694
rect 13442 15672 13454 15694
rect 13520 15672 13532 15694
rect 13532 15672 13554 15694
rect 13320 15660 13354 15672
rect 13420 15660 13454 15672
rect 13520 15660 13554 15672
rect 13020 15582 13026 15594
rect 13026 15582 13054 15594
rect 13020 15560 13054 15582
rect 13120 15560 13154 15594
rect 13220 15560 13254 15594
rect 13320 15582 13352 15594
rect 13352 15582 13354 15594
rect 13420 15582 13442 15594
rect 13442 15582 13454 15594
rect 13520 15582 13532 15594
rect 13532 15582 13554 15594
rect 13320 15560 13354 15582
rect 13420 15560 13454 15582
rect 13520 15560 13554 15582
rect 13020 15492 13026 15494
rect 13026 15492 13054 15494
rect 13020 15460 13054 15492
rect 13120 15460 13154 15494
rect 13220 15460 13254 15494
rect 13320 15492 13352 15494
rect 13352 15492 13354 15494
rect 13420 15492 13442 15494
rect 13442 15492 13454 15494
rect 13520 15492 13532 15494
rect 13532 15492 13554 15494
rect 13320 15460 13354 15492
rect 13420 15460 13454 15492
rect 13520 15460 13554 15492
rect 13020 15360 13054 15394
rect 13120 15360 13154 15394
rect 13220 15360 13254 15394
rect 13320 15360 13354 15394
rect 13420 15360 13454 15394
rect 13520 15360 13554 15394
rect 13020 15260 13054 15294
rect 13120 15260 13154 15294
rect 13220 15260 13254 15294
rect 13320 15260 13354 15294
rect 13420 15260 13454 15294
rect 13520 15260 13554 15294
rect 13020 15166 13054 15194
rect 13020 15160 13026 15166
rect 13026 15160 13054 15166
rect 13120 15160 13154 15194
rect 13220 15160 13254 15194
rect 13320 15166 13354 15194
rect 13420 15166 13454 15194
rect 13520 15166 13554 15194
rect 13320 15160 13352 15166
rect 13352 15160 13354 15166
rect 13420 15160 13442 15166
rect 13442 15160 13454 15166
rect 13520 15160 13532 15166
rect 13532 15160 13554 15166
rect 14380 15672 14386 15694
rect 14386 15672 14414 15694
rect 14380 15660 14414 15672
rect 14480 15660 14514 15694
rect 14580 15660 14614 15694
rect 14680 15672 14712 15694
rect 14712 15672 14714 15694
rect 14780 15672 14802 15694
rect 14802 15672 14814 15694
rect 14880 15672 14892 15694
rect 14892 15672 14914 15694
rect 14680 15660 14714 15672
rect 14780 15660 14814 15672
rect 14880 15660 14914 15672
rect 14380 15582 14386 15594
rect 14386 15582 14414 15594
rect 14380 15560 14414 15582
rect 14480 15560 14514 15594
rect 14580 15560 14614 15594
rect 14680 15582 14712 15594
rect 14712 15582 14714 15594
rect 14780 15582 14802 15594
rect 14802 15582 14814 15594
rect 14880 15582 14892 15594
rect 14892 15582 14914 15594
rect 14680 15560 14714 15582
rect 14780 15560 14814 15582
rect 14880 15560 14914 15582
rect 14380 15492 14386 15494
rect 14386 15492 14414 15494
rect 14380 15460 14414 15492
rect 14480 15460 14514 15494
rect 14580 15460 14614 15494
rect 14680 15492 14712 15494
rect 14712 15492 14714 15494
rect 14780 15492 14802 15494
rect 14802 15492 14814 15494
rect 14880 15492 14892 15494
rect 14892 15492 14914 15494
rect 14680 15460 14714 15492
rect 14780 15460 14814 15492
rect 14880 15460 14914 15492
rect 14380 15360 14414 15394
rect 14480 15360 14514 15394
rect 14580 15360 14614 15394
rect 14680 15360 14714 15394
rect 14780 15360 14814 15394
rect 14880 15360 14914 15394
rect 14380 15260 14414 15294
rect 14480 15260 14514 15294
rect 14580 15260 14614 15294
rect 14680 15260 14714 15294
rect 14780 15260 14814 15294
rect 14880 15260 14914 15294
rect 14380 15166 14414 15194
rect 14380 15160 14386 15166
rect 14386 15160 14414 15166
rect 14480 15160 14514 15194
rect 14580 15160 14614 15194
rect 14680 15166 14714 15194
rect 14780 15166 14814 15194
rect 14880 15166 14914 15194
rect 14680 15160 14712 15166
rect 14712 15160 14714 15166
rect 14780 15160 14802 15166
rect 14802 15160 14814 15166
rect 14880 15160 14892 15166
rect 14892 15160 14914 15166
rect 16800 18041 16838 18438
rect 16800 15970 16838 16367
rect 17590 18555 17630 18589
rect 17590 18550 17630 18555
rect 17556 18035 17662 18432
rect 17556 16650 17662 17047
rect 11560 14350 11960 14402
rect 14599 14360 14996 14398
rect 11100 13760 11140 13800
rect 15490 13800 15530 13840
rect 15490 13720 15530 13760
rect 11180 13590 11220 13630
rect 11340 13590 11380 13630
rect 11500 13590 11540 13630
rect 11660 13590 11700 13630
rect 11820 13590 11860 13630
rect 11980 13590 12020 13630
rect 12140 13590 12180 13630
rect 12300 13590 12340 13630
rect 12460 13590 12500 13630
rect 12620 13590 12660 13630
rect 12780 13590 12820 13630
rect 12940 13590 12980 13630
rect 13100 13590 13140 13630
rect 13260 13590 13300 13630
rect 13420 13590 13460 13630
rect 13580 13590 13620 13630
rect 13740 13590 13780 13630
rect 13900 13590 13940 13630
rect 14060 13590 14100 13630
rect 14220 13590 14260 13630
rect 14380 13590 14420 13630
rect 14540 13590 14580 13630
rect 14700 13590 14740 13630
rect 14860 13590 14900 13630
rect 15020 13590 15060 13630
rect 15180 13590 15220 13630
rect 11920 13320 11960 13360
rect 14600 13320 14640 13360
rect 10760 12720 10800 12760
rect 10940 12680 10980 12720
rect 11180 12680 11220 12720
rect 11420 12680 11460 12720
rect 11660 12680 11700 12720
rect 12300 12680 12340 12720
rect 12540 12680 12580 12720
rect 12780 12680 12820 12720
rect 13080 12710 13120 12750
rect 15760 13200 15800 13240
rect 15760 13100 15800 13140
rect 15760 13000 15800 13040
rect 15760 12900 15800 12940
rect 15760 12800 15800 12840
rect 13440 12710 13480 12750
rect 13740 12680 13780 12720
rect 13980 12680 14020 12720
rect 14220 12680 14260 12720
rect 14860 12680 14900 12720
rect 15100 12680 15140 12720
rect 15340 12680 15380 12720
rect 15580 12680 15620 12720
rect 11443 12308 11477 12342
rect 11803 12308 11837 12342
rect 11923 12308 11957 12342
rect 12283 12308 12317 12342
rect 12403 12308 12437 12342
rect 12820 12280 12860 12320
rect 11380 12190 11420 12230
rect 11500 12190 11540 12230
rect 11620 12190 11660 12230
rect 11740 12190 11780 12230
rect 11860 12190 11900 12230
rect 11980 12190 12020 12230
rect 12100 12190 12140 12230
rect 12220 12190 12260 12230
rect 12340 12190 12380 12230
rect 12460 12190 12500 12230
rect 12580 12190 12620 12230
rect 12820 12200 12860 12240
rect 11544 12078 11578 12112
rect 11702 12078 11736 12112
rect 12026 12078 12060 12112
rect 12180 12078 12214 12112
rect 12504 12078 12538 12112
rect 12820 12120 12860 12160
rect 13700 12280 13740 12320
rect 14123 12308 14157 12342
rect 14243 12308 14277 12342
rect 14603 12308 14637 12342
rect 14723 12308 14757 12342
rect 15083 12308 15117 12342
rect 13700 12200 13740 12240
rect 13940 12190 13980 12230
rect 14060 12190 14100 12230
rect 14180 12190 14220 12230
rect 14300 12190 14340 12230
rect 14420 12190 14460 12230
rect 14540 12190 14580 12230
rect 14660 12190 14700 12230
rect 14780 12190 14820 12230
rect 14900 12190 14940 12230
rect 15020 12190 15060 12230
rect 15140 12190 15180 12230
rect 13700 12120 13740 12160
rect 14022 12078 14056 12112
rect 14346 12078 14380 12112
rect 14500 12078 14534 12112
rect 14824 12078 14858 12112
rect 14982 12078 15016 12112
rect 10720 11480 10760 11520
rect 10900 11470 10940 11510
rect 11380 11470 11420 11510
rect 11620 11470 11660 11510
rect 12100 11470 12140 11510
rect 12340 11470 12380 11510
rect 12760 11470 12800 11510
rect 13760 11470 13800 11510
rect 14180 11470 14220 11510
rect 14420 11470 14460 11510
rect 14900 11470 14940 11510
rect 15140 11470 15180 11510
rect 15620 11470 15660 11510
rect 15800 11480 15840 11520
rect 10540 11350 10580 11390
rect 10540 11250 10580 11290
rect 10660 11350 10700 11390
rect 10660 11250 10700 11290
rect 10780 11350 10820 11390
rect 10780 11250 10820 11290
rect 10900 11350 10940 11390
rect 10900 11250 10940 11290
rect 11020 11350 11060 11390
rect 11020 11250 11060 11290
rect 11140 11350 11180 11390
rect 11140 11250 11180 11290
rect 11260 11350 11300 11390
rect 11260 11250 11300 11290
rect 11380 11350 11420 11390
rect 11380 11250 11420 11290
rect 11500 11350 11540 11390
rect 11500 11250 11540 11290
rect 11620 11350 11660 11390
rect 11620 11250 11660 11290
rect 11740 11350 11780 11390
rect 11740 11250 11780 11290
rect 11860 11350 11900 11390
rect 11860 11250 11900 11290
rect 11980 11350 12020 11390
rect 11980 11250 12020 11290
rect 12100 11350 12140 11390
rect 12100 11250 12140 11290
rect 12220 11350 12260 11390
rect 12220 11250 12260 11290
rect 12340 11350 12380 11390
rect 12340 11250 12380 11290
rect 12460 11350 12500 11390
rect 12460 11250 12500 11290
rect 12580 11350 12620 11390
rect 12580 11250 12620 11290
rect 12700 11350 12740 11390
rect 12700 11250 12740 11290
rect 12820 11350 12860 11390
rect 12820 11250 12860 11290
rect 12940 11350 12980 11390
rect 12940 11250 12980 11290
rect 13580 11350 13620 11390
rect 13580 11250 13620 11290
rect 13700 11350 13740 11390
rect 13700 11250 13740 11290
rect 13820 11350 13860 11390
rect 13820 11250 13860 11290
rect 13940 11350 13980 11390
rect 13940 11250 13980 11290
rect 14060 11350 14100 11390
rect 14060 11250 14100 11290
rect 14180 11350 14220 11390
rect 14180 11250 14220 11290
rect 14300 11350 14340 11390
rect 14300 11250 14340 11290
rect 14420 11350 14460 11390
rect 14420 11250 14460 11290
rect 14540 11350 14580 11390
rect 14540 11250 14580 11290
rect 14660 11350 14700 11390
rect 14660 11250 14700 11290
rect 14780 11350 14820 11390
rect 14780 11250 14820 11290
rect 14900 11350 14940 11390
rect 14900 11250 14940 11290
rect 15020 11350 15060 11390
rect 15020 11250 15060 11290
rect 15140 11350 15180 11390
rect 15140 11250 15180 11290
rect 15260 11350 15300 11390
rect 15260 11250 15300 11290
rect 15380 11350 15420 11390
rect 15380 11250 15420 11290
rect 15500 11350 15540 11390
rect 15500 11250 15540 11290
rect 15620 11350 15660 11390
rect 15620 11250 15660 11290
rect 15740 11350 15780 11390
rect 15740 11250 15780 11290
rect 15860 11350 15900 11390
rect 15860 11250 15900 11290
rect 15980 11350 16020 11390
rect 15980 11250 16020 11290
rect 10540 11130 10580 11170
rect 12940 11130 12980 11170
rect 13580 11130 13620 11170
rect 15980 11130 16020 11170
rect 11910 10310 11950 10350
rect 12090 10310 12130 10350
rect 12270 10310 12310 10350
rect 12450 10310 12490 10350
rect 12630 10310 12670 10350
rect 12810 10310 12850 10350
rect 12990 10310 13030 10350
rect 13170 10310 13210 10350
rect 13350 10310 13390 10350
rect 13530 10310 13570 10350
rect 13710 10310 13750 10350
rect 13890 10310 13930 10350
rect 14070 10310 14110 10350
rect 14250 10310 14290 10350
rect 14430 10310 14470 10350
rect 14610 10310 14650 10350
rect 11640 10190 11680 10230
rect 11640 10090 11680 10130
rect 11640 9990 11680 10030
rect 11640 9890 11680 9930
rect 11640 9790 11680 9830
rect 11640 9690 11680 9730
rect 11820 10190 11860 10230
rect 11820 10090 11860 10130
rect 11820 9990 11860 10030
rect 11820 9890 11860 9930
rect 11820 9790 11860 9830
rect 11820 9690 11860 9730
rect 12000 10190 12040 10230
rect 12000 10090 12040 10130
rect 12000 9990 12040 10030
rect 12000 9890 12040 9930
rect 12000 9790 12040 9830
rect 12000 9690 12040 9730
rect 12180 10190 12220 10230
rect 12180 10090 12220 10130
rect 12180 9990 12220 10030
rect 12180 9890 12220 9930
rect 12180 9790 12220 9830
rect 12180 9690 12220 9730
rect 12360 10190 12400 10230
rect 12360 10090 12400 10130
rect 12360 9990 12400 10030
rect 12360 9890 12400 9930
rect 12360 9790 12400 9830
rect 12360 9690 12400 9730
rect 12540 10190 12580 10230
rect 12540 10090 12580 10130
rect 12540 9990 12580 10030
rect 12540 9890 12580 9930
rect 12540 9790 12580 9830
rect 12540 9690 12580 9730
rect 12720 10190 12760 10230
rect 12720 10090 12760 10130
rect 12720 9990 12760 10030
rect 12720 9890 12760 9930
rect 12720 9790 12760 9830
rect 12720 9690 12760 9730
rect 12900 10190 12940 10230
rect 12900 10090 12940 10130
rect 12900 9990 12940 10030
rect 12900 9890 12940 9930
rect 12900 9790 12940 9830
rect 12900 9690 12940 9730
rect 13080 10190 13120 10230
rect 13080 10090 13120 10130
rect 13080 9990 13120 10030
rect 13080 9890 13120 9930
rect 13080 9790 13120 9830
rect 13080 9690 13120 9730
rect 13260 10190 13300 10230
rect 13260 10090 13300 10130
rect 13260 9990 13300 10030
rect 13260 9890 13300 9930
rect 13260 9790 13300 9830
rect 13260 9690 13300 9730
rect 13440 10190 13480 10230
rect 13440 10090 13480 10130
rect 13440 9990 13480 10030
rect 13440 9890 13480 9930
rect 13440 9790 13480 9830
rect 13440 9690 13480 9730
rect 13620 10190 13660 10230
rect 13620 10090 13660 10130
rect 13620 9990 13660 10030
rect 13620 9890 13660 9930
rect 13620 9790 13660 9830
rect 13620 9690 13660 9730
rect 13800 10190 13840 10230
rect 13800 10090 13840 10130
rect 13800 9990 13840 10030
rect 13800 9890 13840 9930
rect 13800 9790 13840 9830
rect 13800 9690 13840 9730
rect 13980 10190 14020 10230
rect 13980 10090 14020 10130
rect 13980 9990 14020 10030
rect 13980 9890 14020 9930
rect 13980 9790 14020 9830
rect 13980 9690 14020 9730
rect 14160 10190 14200 10230
rect 14160 10090 14200 10130
rect 14160 9990 14200 10030
rect 14160 9890 14200 9930
rect 14160 9790 14200 9830
rect 14160 9690 14200 9730
rect 14340 10190 14380 10230
rect 14340 10090 14380 10130
rect 14340 9990 14380 10030
rect 14340 9890 14380 9930
rect 14340 9790 14380 9830
rect 14340 9690 14380 9730
rect 14520 10190 14560 10230
rect 14520 10090 14560 10130
rect 14520 9990 14560 10030
rect 14520 9890 14560 9930
rect 14520 9790 14560 9830
rect 14520 9690 14560 9730
rect 14700 10190 14740 10230
rect 14700 10090 14740 10130
rect 14700 9990 14740 10030
rect 14700 9890 14740 9930
rect 14700 9790 14740 9830
rect 14700 9690 14740 9730
rect 14880 10190 14920 10230
rect 14880 10090 14920 10130
rect 15610 10110 15650 10150
rect 15730 10110 15770 10150
rect 15850 10110 15890 10150
rect 14880 9990 14920 10030
rect 14880 9890 14920 9930
rect 15510 9990 15550 10030
rect 15510 9890 15550 9930
rect 15620 9990 15660 10030
rect 15620 9890 15660 9930
rect 15730 9990 15770 10030
rect 15730 9890 15770 9930
rect 15840 9990 15880 10030
rect 15840 9890 15880 9930
rect 15950 9990 15990 10030
rect 15950 9890 15990 9930
rect 14880 9790 14920 9830
rect 15510 9770 15550 9810
rect 15730 9770 15770 9810
rect 15950 9770 15990 9810
rect 14880 9690 14920 9730
rect 11640 9570 11680 9610
rect 12000 9570 12040 9610
rect 12360 9570 12400 9610
rect 12720 9570 12760 9610
rect 13080 9570 13120 9610
rect 13440 9570 13480 9610
rect 13800 9570 13840 9610
rect 14160 9570 14200 9610
rect 14520 9570 14560 9610
rect 14880 9570 14920 9610
rect 11818 9308 11852 9342
rect 11928 9308 11962 9342
rect 12038 9308 12072 9342
rect 12148 9308 12182 9342
rect 12258 9308 12292 9342
rect 12368 9308 12402 9342
rect 12478 9308 12512 9342
rect 12588 9308 12622 9342
rect 12698 9308 12732 9342
rect 12808 9308 12842 9342
rect 13718 9308 13752 9342
rect 13828 9308 13862 9342
rect 13938 9308 13972 9342
rect 14048 9308 14082 9342
rect 14158 9308 14192 9342
rect 14268 9308 14302 9342
rect 14378 9308 14412 9342
rect 14488 9308 14522 9342
rect 14598 9308 14632 9342
rect 14708 9308 14742 9342
rect 11570 9190 11610 9230
rect 11650 9190 11690 9230
rect 11570 9090 11610 9130
rect 11650 9090 11690 9130
rect 11760 9190 11800 9230
rect 11760 9090 11800 9130
rect 11870 9190 11910 9230
rect 11870 9090 11910 9130
rect 11980 9190 12020 9230
rect 11980 9090 12020 9130
rect 12090 9190 12130 9230
rect 12090 9090 12130 9130
rect 12200 9190 12240 9230
rect 12200 9090 12240 9130
rect 12310 9190 12350 9230
rect 12310 9090 12350 9130
rect 12420 9190 12460 9230
rect 12420 9090 12460 9130
rect 12530 9190 12570 9230
rect 12530 9090 12570 9130
rect 12640 9190 12680 9230
rect 12640 9090 12680 9130
rect 12750 9190 12790 9230
rect 12750 9090 12790 9130
rect 12860 9190 12900 9230
rect 12860 9090 12900 9130
rect 12970 9190 13010 9230
rect 13050 9190 13090 9230
rect 12970 9090 13010 9130
rect 13050 9090 13090 9130
rect 13470 9190 13510 9230
rect 13550 9190 13590 9230
rect 13470 9090 13510 9130
rect 13550 9090 13590 9130
rect 13660 9190 13700 9230
rect 13660 9090 13700 9130
rect 13770 9190 13810 9230
rect 13770 9090 13810 9130
rect 13880 9190 13920 9230
rect 13880 9090 13920 9130
rect 13990 9190 14030 9230
rect 13990 9090 14030 9130
rect 14100 9190 14140 9230
rect 14100 9090 14140 9130
rect 14210 9190 14250 9230
rect 14210 9090 14250 9130
rect 14320 9190 14360 9230
rect 14320 9090 14360 9130
rect 14430 9190 14470 9230
rect 14430 9090 14470 9130
rect 14540 9190 14580 9230
rect 14540 9090 14580 9130
rect 14650 9190 14690 9230
rect 14650 9090 14690 9130
rect 14760 9190 14800 9230
rect 14760 9090 14800 9130
rect 14870 9190 14910 9230
rect 14950 9190 14990 9230
rect 14870 9090 14910 9130
rect 14950 9090 14990 9130
rect 11650 8970 11690 9010
rect 12970 8970 13010 9010
rect 13550 8970 13590 9010
rect 14870 8970 14910 9010
<< metal1 >>
rect 9170 19190 9250 19200
rect 9170 19130 9180 19190
rect 9240 19130 9250 19190
rect 8790 19080 8870 19090
rect 8790 19020 8800 19080
rect 8860 19020 8870 19080
rect 8790 19000 8870 19020
rect 8790 18940 8800 19000
rect 8860 18940 8870 19000
rect 8790 18920 8870 18940
rect 8790 18860 8800 18920
rect 8860 18860 8870 18920
rect 8790 18590 8870 18860
rect 8790 18550 8810 18590
rect 8850 18550 8870 18590
rect 8790 18530 8870 18550
rect 9170 18450 9250 19130
rect 8770 18432 8888 18444
rect 8770 18035 8776 18432
rect 8882 18035 8888 18432
rect 8770 18023 8888 18035
rect 9170 18390 9180 18450
rect 9240 18390 9250 18450
rect 9170 18370 9250 18390
rect 9170 18310 9180 18370
rect 9240 18310 9250 18370
rect 9170 18280 9250 18310
rect 9170 18220 9180 18280
rect 9240 18220 9250 18280
rect 9170 18190 9250 18220
rect 9170 18130 9180 18190
rect 9240 18130 9250 18190
rect 9170 18110 9250 18130
rect 9170 18050 9180 18110
rect 9240 18050 9250 18110
rect 9170 18030 9250 18050
rect 9570 19080 9650 19090
rect 9570 19020 9580 19080
rect 9640 19020 9650 19080
rect 9570 19000 9650 19020
rect 9570 18940 9580 19000
rect 9640 18940 9650 19000
rect 9570 18920 9650 18940
rect 9570 18860 9580 18920
rect 9640 18860 9650 18920
rect 9570 18600 9650 18860
rect 9570 18560 9590 18600
rect 9630 18560 9650 18600
rect 9570 18438 9650 18560
rect 9570 18041 9590 18438
rect 9628 18041 9650 18438
rect 9570 18020 9650 18041
rect 10680 19080 10760 19090
rect 10680 19020 10690 19080
rect 10750 19020 10760 19080
rect 10680 19000 10760 19020
rect 10680 18940 10690 19000
rect 10750 18940 10760 19000
rect 10680 18920 10760 18940
rect 10680 18860 10690 18920
rect 10750 18860 10760 18920
rect 10680 18610 10760 18860
rect 10680 18570 10700 18610
rect 10740 18570 10760 18610
rect 10680 18440 10760 18570
rect 10680 18050 10700 18440
rect 10740 18050 10760 18440
rect 10680 18030 10760 18050
rect 8770 17047 8888 17059
rect 8770 16650 8776 17047
rect 8882 16650 8888 17047
rect 8770 16638 8888 16650
rect 10350 16700 10430 16720
rect 8790 11180 8870 16638
rect 10350 16310 10370 16700
rect 10410 16310 10430 16700
rect 9570 15477 9650 15500
rect 9570 15080 9590 15477
rect 9628 15080 9650 15477
rect 8790 11120 8800 11180
rect 8860 11120 8870 11180
rect 8790 9360 8870 11120
rect 9460 13810 9540 13820
rect 9460 13750 9470 13810
rect 9530 13750 9540 13810
rect 9460 10690 9540 13750
rect 9570 12120 9650 15080
rect 10350 14720 10430 16310
rect 10350 14660 10360 14720
rect 10420 14660 10430 14720
rect 10350 14650 10430 14660
rect 9570 12060 9580 12120
rect 9640 12060 9650 12120
rect 9570 10800 9650 12060
rect 9570 10740 9580 10800
rect 9640 10740 9650 10800
rect 9570 10730 9650 10740
rect 9680 14090 9760 14100
rect 9680 14030 9690 14090
rect 9750 14030 9760 14090
rect 9680 12350 9760 14030
rect 9680 12290 9690 12350
rect 9750 12290 9760 12350
rect 9460 10630 9470 10690
rect 9530 10630 9540 10690
rect 9460 10620 9540 10630
rect 8790 9300 8800 9360
rect 8860 9300 8870 9360
rect 8790 9290 8870 9300
rect 9680 8910 9760 12290
rect 10620 13980 10700 13990
rect 10620 13920 10630 13980
rect 10690 13920 10700 13980
rect 10620 11650 10700 13920
rect 11030 13980 11110 19200
rect 18190 19190 18270 19200
rect 18190 19130 18200 19190
rect 18260 19130 18270 19190
rect 13240 19080 13320 19090
rect 13240 19020 13250 19080
rect 13310 19020 13320 19080
rect 13240 19000 13320 19020
rect 13240 18940 13250 19000
rect 13310 18940 13320 19000
rect 13240 18920 13320 18940
rect 13240 18860 13250 18920
rect 13310 18860 13320 18920
rect 13240 18850 13320 18860
rect 15670 19080 15750 19090
rect 15670 19020 15680 19080
rect 15740 19020 15750 19080
rect 15670 19000 15750 19020
rect 15670 18940 15680 19000
rect 15740 18940 15750 19000
rect 15670 18920 15750 18940
rect 15670 18860 15680 18920
rect 15740 18860 15750 18920
rect 15670 18610 15750 18860
rect 15670 18570 15690 18610
rect 15730 18570 15750 18610
rect 11570 18414 14990 18490
rect 11570 18380 11660 18414
rect 11694 18380 11760 18414
rect 11794 18380 11860 18414
rect 11894 18380 11960 18414
rect 11994 18380 12060 18414
rect 12094 18380 12160 18414
rect 12194 18380 13020 18414
rect 13054 18380 13120 18414
rect 13154 18380 13220 18414
rect 13254 18380 13320 18414
rect 13354 18380 13420 18414
rect 13454 18380 13520 18414
rect 13554 18380 14380 18414
rect 14414 18380 14480 18414
rect 14514 18380 14580 18414
rect 14614 18380 14680 18414
rect 14714 18380 14780 18414
rect 14814 18380 14880 18414
rect 14914 18380 14990 18414
rect 11570 18314 14990 18380
rect 11570 18280 11660 18314
rect 11694 18280 11760 18314
rect 11794 18280 11860 18314
rect 11894 18280 11960 18314
rect 11994 18280 12060 18314
rect 12094 18280 12160 18314
rect 12194 18280 13020 18314
rect 13054 18280 13120 18314
rect 13154 18280 13220 18314
rect 13254 18280 13320 18314
rect 13354 18280 13420 18314
rect 13454 18280 13520 18314
rect 13554 18280 14380 18314
rect 14414 18280 14480 18314
rect 14514 18280 14580 18314
rect 14614 18280 14680 18314
rect 14714 18280 14780 18314
rect 14814 18280 14880 18314
rect 14914 18280 14990 18314
rect 11570 18214 14990 18280
rect 11570 18180 11660 18214
rect 11694 18180 11760 18214
rect 11794 18180 11860 18214
rect 11894 18180 11960 18214
rect 11994 18180 12060 18214
rect 12094 18180 12160 18214
rect 12194 18180 13020 18214
rect 13054 18180 13120 18214
rect 13154 18180 13220 18214
rect 13254 18180 13320 18214
rect 13354 18180 13420 18214
rect 13454 18180 13520 18214
rect 13554 18180 14380 18214
rect 14414 18180 14480 18214
rect 14514 18180 14580 18214
rect 14614 18180 14680 18214
rect 14714 18180 14780 18214
rect 14814 18180 14880 18214
rect 14914 18180 14990 18214
rect 11570 18114 14990 18180
rect 11570 18080 11660 18114
rect 11694 18080 11760 18114
rect 11794 18080 11860 18114
rect 11894 18080 11960 18114
rect 11994 18080 12060 18114
rect 12094 18080 12160 18114
rect 12194 18080 13020 18114
rect 13054 18080 13120 18114
rect 13154 18080 13220 18114
rect 13254 18080 13320 18114
rect 13354 18080 13420 18114
rect 13454 18080 13520 18114
rect 13554 18080 14380 18114
rect 14414 18080 14480 18114
rect 14514 18080 14580 18114
rect 14614 18080 14680 18114
rect 14714 18080 14780 18114
rect 14814 18080 14880 18114
rect 14914 18080 14990 18114
rect 11570 18014 14990 18080
rect 15670 18440 15750 18570
rect 15670 18050 15690 18440
rect 15730 18050 15750 18440
rect 15670 18030 15750 18050
rect 16780 19080 16860 19090
rect 16780 19020 16790 19080
rect 16850 19020 16860 19080
rect 16780 19000 16860 19020
rect 16780 18940 16790 19000
rect 16850 18940 16860 19000
rect 16780 18920 16860 18940
rect 16780 18860 16790 18920
rect 16850 18860 16860 18920
rect 16780 18610 16860 18860
rect 16780 18570 16800 18610
rect 16840 18570 16860 18610
rect 16780 18438 16860 18570
rect 17570 19080 17650 19090
rect 17570 19020 17580 19080
rect 17640 19020 17650 19080
rect 17570 19000 17650 19020
rect 17570 18940 17580 19000
rect 17640 18940 17650 19000
rect 17570 18920 17650 18940
rect 17570 18860 17580 18920
rect 17640 18860 17650 18920
rect 17570 18590 17650 18860
rect 18190 18850 18270 19130
rect 18190 18790 18200 18850
rect 18260 18790 18270 18850
rect 18190 18780 18270 18790
rect 17570 18550 17590 18590
rect 17630 18550 17650 18590
rect 17570 18530 17650 18550
rect 17950 18450 18030 18460
rect 16780 18041 16800 18438
rect 16838 18041 16860 18438
rect 16780 18030 16860 18041
rect 17550 18432 17668 18444
rect 17550 18035 17556 18432
rect 17662 18035 17668 18432
rect 16794 18029 16844 18030
rect 17550 18023 17668 18035
rect 17950 18390 17960 18450
rect 18020 18390 18030 18450
rect 17950 18370 18030 18390
rect 17950 18310 17960 18370
rect 18020 18310 18030 18370
rect 17950 18280 18030 18310
rect 17950 18220 17960 18280
rect 18020 18220 18030 18280
rect 17950 18190 18030 18220
rect 17950 18130 17960 18190
rect 18020 18130 18030 18190
rect 17950 18110 18030 18130
rect 17950 18050 17960 18110
rect 18020 18050 18030 18110
rect 18640 18150 18740 18170
rect 18640 18090 18660 18150
rect 18720 18090 18740 18150
rect 18640 18070 18740 18090
rect 11570 17980 11660 18014
rect 11694 17980 11760 18014
rect 11794 17980 11860 18014
rect 11894 17980 11960 18014
rect 11994 17980 12060 18014
rect 12094 17980 12160 18014
rect 12194 17980 13020 18014
rect 13054 17980 13120 18014
rect 13154 17980 13220 18014
rect 13254 17980 13320 18014
rect 13354 17980 13420 18014
rect 13454 17980 13520 18014
rect 13554 17980 14380 18014
rect 14414 17980 14480 18014
rect 14514 17980 14580 18014
rect 14614 17980 14680 18014
rect 14714 17980 14780 18014
rect 14814 17980 14880 18014
rect 14914 17980 14990 18014
rect 11570 17914 14990 17980
rect 11570 17880 11660 17914
rect 11694 17880 11760 17914
rect 11794 17880 11860 17914
rect 11894 17880 11960 17914
rect 11994 17880 12060 17914
rect 12094 17880 12160 17914
rect 12194 17880 13020 17914
rect 13054 17880 13120 17914
rect 13154 17880 13220 17914
rect 13254 17880 13320 17914
rect 13354 17880 13420 17914
rect 13454 17880 13520 17914
rect 13554 17880 14380 17914
rect 14414 17880 14480 17914
rect 14514 17880 14580 17914
rect 14614 17880 14680 17914
rect 14714 17880 14780 17914
rect 14814 17880 14880 17914
rect 14914 17880 14990 17914
rect 11570 17790 14990 17880
rect 11570 17054 12270 17790
rect 11570 17020 11660 17054
rect 11694 17020 11760 17054
rect 11794 17020 11860 17054
rect 11894 17020 11960 17054
rect 11994 17020 12060 17054
rect 12094 17020 12160 17054
rect 12194 17020 12270 17054
rect 11570 16954 12270 17020
rect 11570 16920 11660 16954
rect 11694 16920 11760 16954
rect 11794 16920 11860 16954
rect 11894 16920 11960 16954
rect 11994 16920 12060 16954
rect 12094 16920 12160 16954
rect 12194 16920 12270 16954
rect 11570 16854 12270 16920
rect 11570 16820 11660 16854
rect 11694 16820 11760 16854
rect 11794 16820 11860 16854
rect 11894 16820 11960 16854
rect 11994 16820 12060 16854
rect 12094 16820 12160 16854
rect 12194 16820 12270 16854
rect 11140 16810 11220 16820
rect 11140 16750 11150 16810
rect 11210 16750 11220 16810
rect 11140 14410 11220 16750
rect 11570 16810 12270 16820
rect 11570 16750 11580 16810
rect 11640 16754 12270 16810
rect 11640 16750 11660 16754
rect 11570 16720 11660 16750
rect 11694 16720 11760 16754
rect 11794 16720 11860 16754
rect 11894 16720 11960 16754
rect 11994 16720 12060 16754
rect 12094 16720 12160 16754
rect 12194 16720 12270 16754
rect 11570 16654 12270 16720
rect 11570 16620 11660 16654
rect 11694 16620 11760 16654
rect 11794 16620 11860 16654
rect 11894 16620 11960 16654
rect 11994 16620 12060 16654
rect 12094 16620 12160 16654
rect 12194 16620 12270 16654
rect 11570 16554 12270 16620
rect 11570 16520 11660 16554
rect 11694 16520 11760 16554
rect 11794 16520 11860 16554
rect 11894 16520 11960 16554
rect 11994 16520 12060 16554
rect 12094 16520 12160 16554
rect 12194 16520 12270 16554
rect 11570 15770 12270 16520
rect 12930 17054 13630 17130
rect 12930 17020 13020 17054
rect 13054 17020 13120 17054
rect 13154 17020 13220 17054
rect 13254 17020 13320 17054
rect 13354 17020 13420 17054
rect 13454 17020 13520 17054
rect 13554 17020 13630 17054
rect 12930 16954 13630 17020
rect 12930 16920 13020 16954
rect 13054 16920 13120 16954
rect 13154 16920 13220 16954
rect 13254 16920 13320 16954
rect 13354 16920 13420 16954
rect 13454 16920 13520 16954
rect 13554 16920 13630 16954
rect 12930 16854 13630 16920
rect 12930 16820 13020 16854
rect 13054 16820 13120 16854
rect 13154 16820 13220 16854
rect 13254 16820 13320 16854
rect 13354 16820 13420 16854
rect 13454 16820 13520 16854
rect 13554 16820 13630 16854
rect 12930 16810 13630 16820
rect 12930 16754 13250 16810
rect 13310 16754 13630 16810
rect 12930 16720 13020 16754
rect 13054 16720 13120 16754
rect 13154 16720 13220 16754
rect 13310 16750 13320 16754
rect 13254 16720 13320 16750
rect 13354 16720 13420 16754
rect 13454 16720 13520 16754
rect 13554 16720 13630 16754
rect 12930 16654 13630 16720
rect 12930 16620 13020 16654
rect 13054 16620 13120 16654
rect 13154 16620 13220 16654
rect 13254 16620 13320 16654
rect 13354 16620 13420 16654
rect 13454 16620 13520 16654
rect 13554 16620 13630 16654
rect 12930 16554 13630 16620
rect 12930 16520 13020 16554
rect 13054 16520 13120 16554
rect 13154 16520 13220 16554
rect 13254 16520 13320 16554
rect 13354 16520 13420 16554
rect 13454 16520 13520 16554
rect 13554 16520 13630 16554
rect 12930 16430 13630 16520
rect 14290 17054 14990 17790
rect 14290 17020 14380 17054
rect 14414 17020 14480 17054
rect 14514 17020 14580 17054
rect 14614 17020 14680 17054
rect 14714 17020 14780 17054
rect 14814 17020 14880 17054
rect 14914 17020 14990 17054
rect 14290 16954 14990 17020
rect 14290 16920 14380 16954
rect 14414 16920 14480 16954
rect 14514 16920 14580 16954
rect 14614 16920 14680 16954
rect 14714 16920 14780 16954
rect 14814 16920 14880 16954
rect 14914 16920 14990 16954
rect 14290 16854 14990 16920
rect 14290 16820 14380 16854
rect 14414 16820 14480 16854
rect 14514 16820 14580 16854
rect 14614 16820 14680 16854
rect 14714 16820 14780 16854
rect 14814 16820 14880 16854
rect 14914 16820 14990 16854
rect 17550 17047 17668 17059
rect 14290 16754 14990 16820
rect 14290 16720 14380 16754
rect 14414 16720 14480 16754
rect 14514 16720 14580 16754
rect 14614 16720 14680 16754
rect 14714 16720 14780 16754
rect 14814 16720 14880 16754
rect 14914 16720 14990 16754
rect 14290 16654 14990 16720
rect 14290 16620 14380 16654
rect 14414 16620 14480 16654
rect 14514 16620 14580 16654
rect 14614 16620 14680 16654
rect 14714 16620 14780 16654
rect 14814 16620 14880 16654
rect 14914 16620 14990 16654
rect 14290 16554 14990 16620
rect 14290 16520 14380 16554
rect 14414 16520 14480 16554
rect 14514 16520 14580 16554
rect 14614 16520 14680 16554
rect 14714 16520 14780 16554
rect 14814 16520 14880 16554
rect 14914 16520 14990 16554
rect 14290 15770 14990 16520
rect 11570 15694 14990 15770
rect 11570 15660 11660 15694
rect 11694 15660 11760 15694
rect 11794 15660 11860 15694
rect 11894 15660 11960 15694
rect 11994 15660 12060 15694
rect 12094 15660 12160 15694
rect 12194 15660 13020 15694
rect 13054 15660 13120 15694
rect 13154 15660 13220 15694
rect 13254 15660 13320 15694
rect 13354 15660 13420 15694
rect 13454 15660 13520 15694
rect 13554 15660 14380 15694
rect 14414 15660 14480 15694
rect 14514 15660 14580 15694
rect 14614 15660 14680 15694
rect 14714 15660 14780 15694
rect 14814 15660 14880 15694
rect 14914 15660 14990 15694
rect 11570 15594 14990 15660
rect 11570 15560 11660 15594
rect 11694 15560 11760 15594
rect 11794 15560 11860 15594
rect 11894 15560 11960 15594
rect 11994 15560 12060 15594
rect 12094 15560 12160 15594
rect 12194 15560 13020 15594
rect 13054 15560 13120 15594
rect 13154 15560 13220 15594
rect 13254 15560 13320 15594
rect 13354 15560 13420 15594
rect 13454 15560 13520 15594
rect 13554 15560 14380 15594
rect 14414 15560 14480 15594
rect 14514 15560 14580 15594
rect 14614 15560 14680 15594
rect 14714 15560 14780 15594
rect 14814 15560 14880 15594
rect 14914 15560 14990 15594
rect 11570 15494 14990 15560
rect 11570 15460 11660 15494
rect 11694 15460 11760 15494
rect 11794 15460 11860 15494
rect 11894 15460 11960 15494
rect 11994 15460 12060 15494
rect 12094 15460 12160 15494
rect 12194 15460 13020 15494
rect 13054 15460 13120 15494
rect 13154 15460 13220 15494
rect 13254 15460 13320 15494
rect 13354 15460 13420 15494
rect 13454 15460 13520 15494
rect 13554 15460 14380 15494
rect 14414 15460 14480 15494
rect 14514 15460 14580 15494
rect 14614 15460 14680 15494
rect 14714 15460 14780 15494
rect 14814 15460 14880 15494
rect 14914 15460 14990 15494
rect 11570 15394 14990 15460
rect 11570 15360 11660 15394
rect 11694 15360 11760 15394
rect 11794 15360 11860 15394
rect 11894 15360 11960 15394
rect 11994 15360 12060 15394
rect 12094 15360 12160 15394
rect 12194 15360 13020 15394
rect 13054 15360 13120 15394
rect 13154 15360 13220 15394
rect 13254 15360 13320 15394
rect 13354 15360 13420 15394
rect 13454 15360 13520 15394
rect 13554 15360 14380 15394
rect 14414 15360 14480 15394
rect 14514 15360 14580 15394
rect 14614 15360 14680 15394
rect 14714 15360 14780 15394
rect 14814 15360 14880 15394
rect 14914 15360 14990 15394
rect 11570 15294 14990 15360
rect 11570 15260 11660 15294
rect 11694 15260 11760 15294
rect 11794 15260 11860 15294
rect 11894 15260 11960 15294
rect 11994 15260 12060 15294
rect 12094 15260 12160 15294
rect 12194 15260 13020 15294
rect 13054 15260 13120 15294
rect 13154 15260 13220 15294
rect 13254 15260 13320 15294
rect 13354 15260 13420 15294
rect 13454 15260 13520 15294
rect 13554 15260 14380 15294
rect 14414 15260 14480 15294
rect 14514 15260 14580 15294
rect 14614 15260 14680 15294
rect 14714 15260 14780 15294
rect 14814 15260 14880 15294
rect 14914 15260 14990 15294
rect 11570 15194 14990 15260
rect 11570 15160 11660 15194
rect 11694 15160 11760 15194
rect 11794 15160 11860 15194
rect 11894 15160 11960 15194
rect 11994 15160 12060 15194
rect 12094 15160 12160 15194
rect 12194 15160 13020 15194
rect 13054 15160 13120 15194
rect 13154 15160 13220 15194
rect 13254 15160 13320 15194
rect 13354 15160 13420 15194
rect 13454 15160 13520 15194
rect 13554 15160 14380 15194
rect 14414 15160 14480 15194
rect 14514 15160 14580 15194
rect 14614 15160 14680 15194
rect 14714 15160 14780 15194
rect 14814 15160 14880 15194
rect 14914 15160 14990 15194
rect 11570 15070 14990 15160
rect 15340 16810 15420 16820
rect 15340 16750 15350 16810
rect 15410 16750 15420 16810
rect 15340 14800 15420 16750
rect 15340 14740 15350 14800
rect 15410 14740 15420 14800
rect 15340 14730 15420 14740
rect 16000 16700 16080 16720
rect 16000 16310 16020 16700
rect 16060 16310 16080 16700
rect 17550 16650 17556 17047
rect 17662 16650 17668 17047
rect 17550 16638 17668 16650
rect 16000 14800 16080 16310
rect 16780 16367 16860 16390
rect 16780 15970 16800 16367
rect 16838 15970 16860 16367
rect 16350 15350 16590 15370
rect 16350 15290 16360 15350
rect 16420 15290 16440 15350
rect 16500 15290 16520 15350
rect 16580 15290 16590 15350
rect 16000 14740 16010 14800
rect 16070 14740 16080 14800
rect 16000 14730 16080 14740
rect 16240 14800 16320 14810
rect 16240 14740 16250 14800
rect 16310 14740 16320 14800
rect 16240 14730 16320 14740
rect 14580 14720 15020 14730
rect 14580 14660 14590 14720
rect 14650 14660 14680 14720
rect 14740 14660 14770 14720
rect 14830 14660 14860 14720
rect 14920 14660 14950 14720
rect 15010 14660 15020 14720
rect 11140 14350 11150 14410
rect 11210 14350 11220 14410
rect 11140 14340 11220 14350
rect 11540 14402 11980 14420
rect 11540 14350 11560 14402
rect 11960 14350 11980 14402
rect 11540 14340 11980 14350
rect 14580 14402 15020 14660
rect 14580 14398 14600 14402
rect 14580 14360 14599 14398
rect 14580 14350 14600 14360
rect 15000 14350 15020 14402
rect 14580 14340 15020 14350
rect 16150 14410 16230 14420
rect 16150 14350 16160 14410
rect 16220 14350 16230 14410
rect 16150 14340 16230 14350
rect 11030 13920 11040 13980
rect 11100 13920 11110 13980
rect 11030 13910 11110 13920
rect 15470 13850 15550 13860
rect 11080 13810 11160 13820
rect 11080 13750 11090 13810
rect 11150 13750 11160 13810
rect 11080 13740 11160 13750
rect 15470 13790 15480 13850
rect 15540 13790 15550 13850
rect 15470 13770 15550 13790
rect 15470 13710 15480 13770
rect 15540 13710 15550 13770
rect 15470 13700 15550 13710
rect 11160 13640 11240 13650
rect 11160 13580 11170 13640
rect 11230 13580 11240 13640
rect 11160 13570 11240 13580
rect 11320 13640 11400 13650
rect 11320 13580 11330 13640
rect 11390 13580 11400 13640
rect 11320 13570 11400 13580
rect 11480 13640 11560 13650
rect 11480 13580 11490 13640
rect 11550 13580 11560 13640
rect 11480 13570 11560 13580
rect 11640 13640 11720 13650
rect 11640 13580 11650 13640
rect 11710 13580 11720 13640
rect 11640 13570 11720 13580
rect 11800 13640 11880 13650
rect 11800 13580 11810 13640
rect 11870 13580 11880 13640
rect 11800 13570 11880 13580
rect 11960 13640 12040 13650
rect 11960 13580 11970 13640
rect 12030 13580 12040 13640
rect 11960 13570 12040 13580
rect 12120 13640 12200 13650
rect 12120 13580 12130 13640
rect 12190 13580 12200 13640
rect 12120 13570 12200 13580
rect 12280 13640 12360 13650
rect 12280 13580 12290 13640
rect 12350 13580 12360 13640
rect 12280 13570 12360 13580
rect 12440 13640 12520 13650
rect 12440 13580 12450 13640
rect 12510 13580 12520 13640
rect 12440 13570 12520 13580
rect 12600 13640 12680 13650
rect 12600 13580 12610 13640
rect 12670 13580 12680 13640
rect 12600 13570 12680 13580
rect 12760 13640 12840 13650
rect 12760 13580 12770 13640
rect 12830 13580 12840 13640
rect 12760 13570 12840 13580
rect 12920 13640 13000 13650
rect 12920 13580 12930 13640
rect 12990 13580 13000 13640
rect 12920 13570 13000 13580
rect 13080 13640 13160 13650
rect 13080 13580 13090 13640
rect 13150 13580 13160 13640
rect 13080 13570 13160 13580
rect 13240 13640 13320 13650
rect 13240 13580 13250 13640
rect 13310 13580 13320 13640
rect 13240 13570 13320 13580
rect 13400 13640 13480 13650
rect 13400 13580 13410 13640
rect 13470 13580 13480 13640
rect 13400 13570 13480 13580
rect 13560 13640 13640 13650
rect 13560 13580 13570 13640
rect 13630 13580 13640 13640
rect 13560 13570 13640 13580
rect 13720 13640 13800 13650
rect 13720 13580 13730 13640
rect 13790 13580 13800 13640
rect 13720 13570 13800 13580
rect 13880 13640 13960 13650
rect 13880 13580 13890 13640
rect 13950 13580 13960 13640
rect 13880 13570 13960 13580
rect 14040 13640 14120 13650
rect 14040 13580 14050 13640
rect 14110 13580 14120 13640
rect 14040 13570 14120 13580
rect 14200 13640 14280 13650
rect 14200 13580 14210 13640
rect 14270 13580 14280 13640
rect 14200 13570 14280 13580
rect 14360 13640 14440 13650
rect 14360 13580 14370 13640
rect 14430 13580 14440 13640
rect 14360 13570 14440 13580
rect 14520 13640 14600 13650
rect 14520 13580 14530 13640
rect 14590 13580 14600 13640
rect 14520 13570 14600 13580
rect 14680 13640 14760 13650
rect 14680 13580 14690 13640
rect 14750 13580 14760 13640
rect 14680 13570 14760 13580
rect 14840 13640 14920 13650
rect 14840 13580 14850 13640
rect 14910 13580 14920 13640
rect 14840 13570 14920 13580
rect 15000 13640 15080 13650
rect 15000 13580 15010 13640
rect 15070 13580 15080 13640
rect 15000 13570 15080 13580
rect 15160 13640 15240 13650
rect 15160 13580 15170 13640
rect 15230 13580 15240 13640
rect 15160 13570 15240 13580
rect 11900 13530 11980 13540
rect 11900 13470 11910 13530
rect 11970 13470 11980 13530
rect 11900 13450 11980 13470
rect 11900 13390 11910 13450
rect 11970 13390 11980 13450
rect 11900 13370 11980 13390
rect 11900 13310 11910 13370
rect 11970 13310 11980 13370
rect 11900 13300 11980 13310
rect 13160 13530 13400 13540
rect 13160 13470 13170 13530
rect 13230 13470 13250 13530
rect 13310 13470 13330 13530
rect 13390 13470 13400 13530
rect 13160 13450 13400 13470
rect 13160 13390 13170 13450
rect 13230 13390 13250 13450
rect 13310 13390 13330 13450
rect 13390 13390 13400 13450
rect 13160 13370 13400 13390
rect 13160 13310 13170 13370
rect 13230 13310 13250 13370
rect 13310 13310 13330 13370
rect 13390 13310 13400 13370
rect 10740 12760 10820 12780
rect 10740 12720 10760 12760
rect 10800 12720 10820 12760
rect 13070 12750 13130 12770
rect 10740 12460 10820 12720
rect 10920 12730 11000 12740
rect 10920 12670 10930 12730
rect 10990 12670 11000 12730
rect 10920 12650 11000 12670
rect 10920 12590 10930 12650
rect 10990 12590 11000 12650
rect 10920 12570 11000 12590
rect 10920 12510 10930 12570
rect 10990 12510 11000 12570
rect 10920 12500 11000 12510
rect 11160 12730 11240 12740
rect 11160 12670 11170 12730
rect 11230 12670 11240 12730
rect 11160 12650 11240 12670
rect 11160 12590 11170 12650
rect 11230 12590 11240 12650
rect 11160 12570 11240 12590
rect 11160 12510 11170 12570
rect 11230 12510 11240 12570
rect 11160 12500 11240 12510
rect 11400 12730 11480 12740
rect 11400 12670 11410 12730
rect 11470 12670 11480 12730
rect 11400 12650 11480 12670
rect 11400 12590 11410 12650
rect 11470 12590 11480 12650
rect 11400 12570 11480 12590
rect 11400 12510 11410 12570
rect 11470 12510 11480 12570
rect 11400 12500 11480 12510
rect 11640 12730 11720 12740
rect 11640 12670 11650 12730
rect 11710 12670 11720 12730
rect 11640 12650 11720 12670
rect 11640 12590 11650 12650
rect 11710 12590 11720 12650
rect 11640 12570 11720 12590
rect 11640 12510 11650 12570
rect 11710 12510 11720 12570
rect 11640 12500 11720 12510
rect 12280 12730 12360 12740
rect 12280 12670 12290 12730
rect 12350 12670 12360 12730
rect 12280 12650 12360 12670
rect 12280 12590 12290 12650
rect 12350 12590 12360 12650
rect 12280 12570 12360 12590
rect 12280 12510 12290 12570
rect 12350 12510 12360 12570
rect 12280 12500 12360 12510
rect 12520 12730 12600 12740
rect 12520 12670 12530 12730
rect 12590 12670 12600 12730
rect 12520 12650 12600 12670
rect 12520 12590 12530 12650
rect 12590 12590 12600 12650
rect 12520 12570 12600 12590
rect 12520 12510 12530 12570
rect 12590 12510 12600 12570
rect 12520 12500 12600 12510
rect 12760 12730 12840 12740
rect 12760 12670 12770 12730
rect 12830 12670 12840 12730
rect 12760 12650 12840 12670
rect 12760 12590 12770 12650
rect 12830 12590 12840 12650
rect 12760 12570 12840 12590
rect 12760 12510 12770 12570
rect 12830 12510 12840 12570
rect 12760 12500 12840 12510
rect 13070 12710 13080 12750
rect 13120 12710 13130 12750
rect 10740 12400 10750 12460
rect 10810 12400 10820 12460
rect 10740 12390 10820 12400
rect 11490 12460 11570 12470
rect 11490 12400 11500 12460
rect 11560 12400 11570 12460
rect 11490 12390 11570 12400
rect 11710 12460 11790 12470
rect 11710 12400 11720 12460
rect 11780 12400 11790 12460
rect 11710 12390 11790 12400
rect 11970 12460 12050 12470
rect 11970 12400 11980 12460
rect 12040 12400 12050 12460
rect 11970 12390 12050 12400
rect 12190 12460 12270 12470
rect 12190 12400 12200 12460
rect 12260 12400 12270 12460
rect 12190 12390 12270 12400
rect 12450 12460 12530 12470
rect 12450 12400 12460 12460
rect 12520 12400 12530 12460
rect 12450 12390 12530 12400
rect 11431 12350 11489 12360
rect 11431 12298 11433 12350
rect 11485 12298 11489 12350
rect 11431 12290 11489 12298
rect 11520 12250 11550 12390
rect 11730 12250 11760 12390
rect 11791 12350 11849 12360
rect 11791 12298 11793 12350
rect 11845 12298 11849 12350
rect 11791 12290 11849 12298
rect 11911 12350 11969 12360
rect 11911 12298 11913 12350
rect 11965 12298 11969 12350
rect 11911 12290 11969 12298
rect 12000 12250 12030 12390
rect 12210 12250 12240 12390
rect 12271 12350 12329 12360
rect 12271 12298 12273 12350
rect 12325 12298 12329 12350
rect 12271 12290 12329 12298
rect 12391 12350 12449 12360
rect 12391 12298 12393 12350
rect 12445 12298 12449 12350
rect 12391 12290 12449 12298
rect 12480 12250 12510 12390
rect 12800 12330 12880 12340
rect 12800 12270 12810 12330
rect 12870 12270 12880 12330
rect 12800 12250 12880 12270
rect 11370 12230 11430 12250
rect 11370 12190 11380 12230
rect 11420 12190 11430 12230
rect 11370 11920 11430 12190
rect 11490 12230 11550 12250
rect 11490 12190 11500 12230
rect 11540 12190 11550 12230
rect 11490 12170 11550 12190
rect 11610 12230 11670 12250
rect 11610 12190 11620 12230
rect 11660 12190 11670 12230
rect 11610 12170 11670 12190
rect 11730 12230 11790 12250
rect 11730 12190 11740 12230
rect 11780 12190 11790 12230
rect 11730 12170 11790 12190
rect 11850 12230 11910 12250
rect 11850 12190 11860 12230
rect 11900 12190 11910 12230
rect 11850 12170 11910 12190
rect 11970 12230 12030 12250
rect 11970 12190 11980 12230
rect 12020 12190 12030 12230
rect 11970 12170 12030 12190
rect 12090 12230 12150 12250
rect 12090 12190 12100 12230
rect 12140 12190 12150 12230
rect 12090 12170 12150 12190
rect 12210 12230 12270 12250
rect 12210 12190 12220 12230
rect 12260 12190 12270 12230
rect 12210 12170 12270 12190
rect 12330 12230 12390 12250
rect 12330 12190 12340 12230
rect 12380 12190 12390 12230
rect 12330 12170 12390 12190
rect 12450 12230 12510 12250
rect 12450 12190 12460 12230
rect 12500 12190 12510 12230
rect 12450 12170 12510 12190
rect 12570 12230 12630 12250
rect 12570 12190 12580 12230
rect 12620 12190 12630 12230
rect 12570 12170 12630 12190
rect 12800 12190 12810 12250
rect 12870 12190 12880 12250
rect 12800 12170 12880 12190
rect 11532 12122 11590 12130
rect 11532 12070 11536 12122
rect 11588 12070 11590 12122
rect 11532 12060 11590 12070
rect 11620 12030 11660 12170
rect 11690 12122 11748 12130
rect 11690 12070 11694 12122
rect 11746 12070 11748 12122
rect 11690 12060 11748 12070
rect 11600 12020 11680 12030
rect 11600 11960 11610 12020
rect 11670 11960 11680 12020
rect 11360 11910 11440 11920
rect 11360 11850 11370 11910
rect 11430 11850 11440 11910
rect 10620 11640 10780 11650
rect 10620 11580 10630 11640
rect 10690 11580 10710 11640
rect 10770 11580 10780 11640
rect 10620 11570 10780 11580
rect 11120 11640 11200 11650
rect 11120 11580 11130 11640
rect 11190 11580 11200 11640
rect 11120 11570 11200 11580
rect 11360 11640 11440 11850
rect 11360 11580 11370 11640
rect 11430 11580 11440 11640
rect 11360 11570 11440 11580
rect 10710 11520 10770 11570
rect 10710 11480 10720 11520
rect 10760 11480 10770 11520
rect 10710 11460 10770 11480
rect 10880 11520 10960 11530
rect 10880 11460 10890 11520
rect 10950 11460 10960 11520
rect 10880 11450 10960 11460
rect 10530 11390 10590 11410
rect 10530 11350 10540 11390
rect 10580 11350 10590 11390
rect 10530 11290 10590 11350
rect 10530 11250 10540 11290
rect 10580 11250 10590 11290
rect 10530 11170 10590 11250
rect 10650 11390 10710 11410
rect 10650 11350 10660 11390
rect 10700 11350 10710 11390
rect 10650 11290 10710 11350
rect 10650 11250 10660 11290
rect 10700 11250 10710 11290
rect 10650 11190 10710 11250
rect 10770 11390 10830 11410
rect 10770 11350 10780 11390
rect 10820 11350 10830 11390
rect 10770 11290 10830 11350
rect 10770 11250 10780 11290
rect 10820 11250 10830 11290
rect 10530 11130 10540 11170
rect 10580 11130 10590 11170
rect 10530 11080 10590 11130
rect 10640 11180 10720 11190
rect 10640 11120 10650 11180
rect 10710 11120 10720 11180
rect 10640 11110 10720 11120
rect 10770 11080 10830 11250
rect 10890 11390 10950 11450
rect 10890 11350 10900 11390
rect 10940 11350 10950 11390
rect 10890 11290 10950 11350
rect 10890 11250 10900 11290
rect 10940 11250 10950 11290
rect 10890 11230 10950 11250
rect 11010 11390 11070 11410
rect 11010 11350 11020 11390
rect 11060 11350 11070 11390
rect 11010 11290 11070 11350
rect 11010 11250 11020 11290
rect 11060 11250 11070 11290
rect 11010 11080 11070 11250
rect 11130 11390 11190 11570
rect 11370 11510 11430 11570
rect 11370 11470 11380 11510
rect 11420 11470 11430 11510
rect 11370 11450 11430 11470
rect 11600 11520 11680 11960
rect 11860 11920 11900 12170
rect 12014 12122 12072 12130
rect 12014 12070 12018 12122
rect 12070 12070 12072 12122
rect 12014 12060 12072 12070
rect 12100 12030 12140 12170
rect 12168 12122 12226 12130
rect 12168 12070 12172 12122
rect 12224 12070 12226 12122
rect 12168 12060 12226 12070
rect 12080 12020 12160 12030
rect 12080 11960 12090 12020
rect 12150 11960 12160 12020
rect 12080 11950 12160 11960
rect 12340 11920 12380 12170
rect 12492 12122 12550 12130
rect 12492 12070 12496 12122
rect 12548 12070 12550 12122
rect 12492 12060 12550 12070
rect 12580 12030 12620 12170
rect 12800 12110 12810 12170
rect 12870 12110 12880 12170
rect 12800 12100 12880 12110
rect 12560 12020 12640 12030
rect 12560 11960 12570 12020
rect 12630 11960 12640 12020
rect 12560 11950 12640 11960
rect 11840 11910 11920 11920
rect 11840 11850 11850 11910
rect 11910 11850 11920 11910
rect 11840 11840 11920 11850
rect 12320 11910 12400 11920
rect 12320 11850 12330 11910
rect 12390 11850 12400 11910
rect 12320 11840 12400 11850
rect 11840 11640 11920 11650
rect 11840 11580 11850 11640
rect 11910 11580 11920 11640
rect 11840 11570 11920 11580
rect 12080 11640 12160 11650
rect 12080 11580 12090 11640
rect 12150 11580 12160 11640
rect 12080 11570 12160 11580
rect 12560 11640 12640 11650
rect 12560 11580 12570 11640
rect 12630 11580 12640 11640
rect 12560 11570 12640 11580
rect 12740 11640 12820 11650
rect 12740 11580 12750 11640
rect 12810 11580 12820 11640
rect 12740 11570 12820 11580
rect 11600 11460 11610 11520
rect 11670 11460 11680 11520
rect 11600 11450 11680 11460
rect 11130 11350 11140 11390
rect 11180 11350 11190 11390
rect 11130 11290 11190 11350
rect 11130 11250 11140 11290
rect 11180 11250 11190 11290
rect 11130 11230 11190 11250
rect 11250 11390 11310 11410
rect 11250 11350 11260 11390
rect 11300 11350 11310 11390
rect 11250 11290 11310 11350
rect 11250 11250 11260 11290
rect 11300 11250 11310 11290
rect 11250 11080 11310 11250
rect 11370 11390 11430 11410
rect 11370 11350 11380 11390
rect 11420 11350 11430 11390
rect 11370 11290 11430 11350
rect 11370 11250 11380 11290
rect 11420 11250 11430 11290
rect 11370 11190 11430 11250
rect 11490 11390 11550 11410
rect 11490 11350 11500 11390
rect 11540 11350 11550 11390
rect 11490 11290 11550 11350
rect 11490 11250 11500 11290
rect 11540 11250 11550 11290
rect 11360 11180 11440 11190
rect 11360 11120 11370 11180
rect 11430 11120 11440 11180
rect 11360 11110 11440 11120
rect 11490 11080 11550 11250
rect 11610 11390 11670 11450
rect 11610 11350 11620 11390
rect 11660 11350 11670 11390
rect 11610 11290 11670 11350
rect 11610 11250 11620 11290
rect 11660 11250 11670 11290
rect 11610 11230 11670 11250
rect 11730 11390 11790 11410
rect 11730 11350 11740 11390
rect 11780 11350 11790 11390
rect 11730 11290 11790 11350
rect 11730 11250 11740 11290
rect 11780 11250 11790 11290
rect 11730 11080 11790 11250
rect 11850 11390 11910 11570
rect 12090 11510 12150 11570
rect 12090 11470 12100 11510
rect 12140 11470 12150 11510
rect 12090 11450 12150 11470
rect 12320 11520 12400 11530
rect 12320 11460 12330 11520
rect 12390 11460 12400 11520
rect 12320 11450 12400 11460
rect 11850 11350 11860 11390
rect 11900 11350 11910 11390
rect 11850 11290 11910 11350
rect 11850 11250 11860 11290
rect 11900 11250 11910 11290
rect 11850 11230 11910 11250
rect 11970 11390 12030 11410
rect 11970 11350 11980 11390
rect 12020 11350 12030 11390
rect 11970 11290 12030 11350
rect 11970 11250 11980 11290
rect 12020 11250 12030 11290
rect 11970 11080 12030 11250
rect 12090 11390 12150 11410
rect 12090 11350 12100 11390
rect 12140 11350 12150 11390
rect 12090 11290 12150 11350
rect 12090 11250 12100 11290
rect 12140 11250 12150 11290
rect 12090 11190 12150 11250
rect 12210 11390 12270 11410
rect 12210 11350 12220 11390
rect 12260 11350 12270 11390
rect 12210 11290 12270 11350
rect 12210 11250 12220 11290
rect 12260 11250 12270 11290
rect 12080 11180 12160 11190
rect 12080 11120 12090 11180
rect 12150 11120 12160 11180
rect 12080 11110 12160 11120
rect 12210 11080 12270 11250
rect 12330 11390 12390 11450
rect 12330 11350 12340 11390
rect 12380 11350 12390 11390
rect 12330 11290 12390 11350
rect 12330 11250 12340 11290
rect 12380 11250 12390 11290
rect 12330 11230 12390 11250
rect 12450 11390 12510 11410
rect 12450 11350 12460 11390
rect 12500 11350 12510 11390
rect 12450 11290 12510 11350
rect 12450 11250 12460 11290
rect 12500 11250 12510 11290
rect 12450 11080 12510 11250
rect 12570 11390 12630 11570
rect 12750 11510 12810 11570
rect 12750 11470 12760 11510
rect 12800 11470 12810 11510
rect 12750 11450 12810 11470
rect 12570 11350 12580 11390
rect 12620 11350 12630 11390
rect 12570 11290 12630 11350
rect 12570 11250 12580 11290
rect 12620 11250 12630 11290
rect 12570 11230 12630 11250
rect 12690 11390 12750 11410
rect 12690 11350 12700 11390
rect 12740 11350 12750 11390
rect 12690 11290 12750 11350
rect 12690 11250 12700 11290
rect 12740 11250 12750 11290
rect 12690 11080 12750 11250
rect 12810 11390 12870 11410
rect 12810 11350 12820 11390
rect 12860 11350 12870 11390
rect 12810 11290 12870 11350
rect 12810 11250 12820 11290
rect 12860 11250 12870 11290
rect 12810 11190 12870 11250
rect 12930 11390 12990 11410
rect 12930 11350 12940 11390
rect 12980 11350 12990 11390
rect 12930 11290 12990 11350
rect 12930 11250 12940 11290
rect 12980 11250 12990 11290
rect 12800 11180 12880 11190
rect 12800 11120 12810 11180
rect 12870 11120 12880 11180
rect 12800 11110 12880 11120
rect 12930 11170 12990 11250
rect 13070 11190 13130 12710
rect 13160 12330 13400 13310
rect 14580 13530 14660 13540
rect 14580 13470 14590 13530
rect 14650 13470 14660 13530
rect 14580 13450 14660 13470
rect 14580 13390 14590 13450
rect 14650 13390 14660 13450
rect 14580 13370 14660 13390
rect 14580 13310 14590 13370
rect 14650 13310 14660 13370
rect 14580 13300 14660 13310
rect 15750 13240 15810 13260
rect 15750 13200 15760 13240
rect 15800 13200 15810 13240
rect 15750 13140 15810 13200
rect 15750 13100 15760 13140
rect 15800 13100 15810 13140
rect 15750 13040 15810 13100
rect 15750 13000 15760 13040
rect 15800 13000 15810 13040
rect 15750 12940 15810 13000
rect 15750 12900 15760 12940
rect 15800 12900 15810 12940
rect 15750 12840 15810 12900
rect 15750 12800 15760 12840
rect 15800 12800 15810 12840
rect 13160 12270 13170 12330
rect 13230 12270 13250 12330
rect 13310 12270 13330 12330
rect 13390 12270 13400 12330
rect 13160 12250 13400 12270
rect 13160 12190 13170 12250
rect 13230 12190 13250 12250
rect 13310 12190 13330 12250
rect 13390 12190 13400 12250
rect 13160 12170 13400 12190
rect 13160 12110 13170 12170
rect 13230 12110 13250 12170
rect 13310 12110 13330 12170
rect 13390 12110 13400 12170
rect 13160 12100 13400 12110
rect 13430 12750 13490 12770
rect 13430 12710 13440 12750
rect 13480 12710 13490 12750
rect 13430 11190 13490 12710
rect 13720 12730 13800 12740
rect 13720 12670 13730 12730
rect 13790 12670 13800 12730
rect 13720 12650 13800 12670
rect 13720 12590 13730 12650
rect 13790 12590 13800 12650
rect 13720 12570 13800 12590
rect 13720 12510 13730 12570
rect 13790 12510 13800 12570
rect 13720 12500 13800 12510
rect 13960 12730 14040 12740
rect 13960 12670 13970 12730
rect 14030 12670 14040 12730
rect 13960 12650 14040 12670
rect 13960 12590 13970 12650
rect 14030 12590 14040 12650
rect 13960 12570 14040 12590
rect 13960 12510 13970 12570
rect 14030 12510 14040 12570
rect 13960 12500 14040 12510
rect 14200 12730 14280 12740
rect 14200 12670 14210 12730
rect 14270 12670 14280 12730
rect 14200 12650 14280 12670
rect 14200 12590 14210 12650
rect 14270 12590 14280 12650
rect 14200 12570 14280 12590
rect 14200 12510 14210 12570
rect 14270 12510 14280 12570
rect 14200 12500 14280 12510
rect 14840 12730 14920 12740
rect 14840 12670 14850 12730
rect 14910 12670 14920 12730
rect 14840 12650 14920 12670
rect 14840 12590 14850 12650
rect 14910 12590 14920 12650
rect 14840 12570 14920 12590
rect 14840 12510 14850 12570
rect 14910 12510 14920 12570
rect 14840 12500 14920 12510
rect 15080 12730 15160 12740
rect 15080 12670 15090 12730
rect 15150 12670 15160 12730
rect 15080 12650 15160 12670
rect 15080 12590 15090 12650
rect 15150 12590 15160 12650
rect 15080 12570 15160 12590
rect 15080 12510 15090 12570
rect 15150 12510 15160 12570
rect 15080 12500 15160 12510
rect 15320 12730 15400 12740
rect 15320 12670 15330 12730
rect 15390 12670 15400 12730
rect 15320 12650 15400 12670
rect 15320 12590 15330 12650
rect 15390 12590 15400 12650
rect 15320 12570 15400 12590
rect 15320 12510 15330 12570
rect 15390 12510 15400 12570
rect 15320 12500 15400 12510
rect 15560 12730 15640 12740
rect 15560 12670 15570 12730
rect 15630 12670 15640 12730
rect 15560 12650 15640 12670
rect 15560 12590 15570 12650
rect 15630 12590 15640 12650
rect 15560 12570 15640 12590
rect 15560 12510 15570 12570
rect 15630 12510 15640 12570
rect 15560 12500 15640 12510
rect 15750 12470 15810 12800
rect 14030 12460 14110 12470
rect 14030 12400 14040 12460
rect 14100 12400 14110 12460
rect 14030 12390 14110 12400
rect 14290 12460 14370 12470
rect 14290 12400 14300 12460
rect 14360 12400 14370 12460
rect 14290 12390 14370 12400
rect 14510 12460 14590 12470
rect 14510 12400 14520 12460
rect 14580 12400 14590 12460
rect 14510 12390 14590 12400
rect 14770 12460 14850 12470
rect 14770 12400 14780 12460
rect 14840 12400 14850 12460
rect 14770 12390 14850 12400
rect 14990 12460 15070 12470
rect 14990 12400 15000 12460
rect 15060 12400 15070 12460
rect 14990 12390 15070 12400
rect 15740 12460 15820 12470
rect 15740 12400 15750 12460
rect 15810 12400 15820 12460
rect 15740 12390 15820 12400
rect 13680 12330 13760 12340
rect 13680 12270 13690 12330
rect 13750 12270 13760 12330
rect 13680 12250 13760 12270
rect 14050 12250 14080 12390
rect 14111 12350 14169 12360
rect 14111 12298 14115 12350
rect 14167 12298 14169 12350
rect 14111 12290 14169 12298
rect 14231 12350 14289 12360
rect 14231 12298 14235 12350
rect 14287 12298 14289 12350
rect 14231 12290 14289 12298
rect 14320 12250 14350 12390
rect 14530 12250 14560 12390
rect 14591 12350 14649 12360
rect 14591 12298 14595 12350
rect 14647 12298 14649 12350
rect 14591 12290 14649 12298
rect 14711 12350 14769 12360
rect 14711 12298 14715 12350
rect 14767 12298 14769 12350
rect 14711 12290 14769 12298
rect 14800 12250 14830 12390
rect 15010 12250 15040 12390
rect 16170 12360 16210 14340
rect 15071 12350 15129 12360
rect 15071 12298 15075 12350
rect 15127 12298 15129 12350
rect 15071 12290 15129 12298
rect 16150 12350 16230 12360
rect 16150 12290 16160 12350
rect 16220 12290 16230 12350
rect 16150 12280 16230 12290
rect 13680 12190 13690 12250
rect 13750 12190 13760 12250
rect 13680 12170 13760 12190
rect 13930 12230 13990 12250
rect 13930 12190 13940 12230
rect 13980 12190 13990 12230
rect 13930 12170 13990 12190
rect 14050 12230 14110 12250
rect 14050 12190 14060 12230
rect 14100 12190 14110 12230
rect 14050 12170 14110 12190
rect 14170 12230 14230 12250
rect 14170 12190 14180 12230
rect 14220 12190 14230 12230
rect 14170 12170 14230 12190
rect 14290 12230 14350 12250
rect 14290 12190 14300 12230
rect 14340 12190 14350 12230
rect 14290 12170 14350 12190
rect 14410 12230 14470 12250
rect 14410 12190 14420 12230
rect 14460 12190 14470 12230
rect 14410 12170 14470 12190
rect 14530 12230 14590 12250
rect 14530 12190 14540 12230
rect 14580 12190 14590 12230
rect 14530 12170 14590 12190
rect 14650 12230 14710 12250
rect 14650 12190 14660 12230
rect 14700 12190 14710 12230
rect 14650 12170 14710 12190
rect 14770 12230 14830 12250
rect 14770 12190 14780 12230
rect 14820 12190 14830 12230
rect 14770 12170 14830 12190
rect 14890 12230 14950 12250
rect 14890 12190 14900 12230
rect 14940 12190 14950 12230
rect 14890 12170 14950 12190
rect 15010 12230 15070 12250
rect 15010 12190 15020 12230
rect 15060 12190 15070 12230
rect 15010 12170 15070 12190
rect 15130 12230 15190 12250
rect 15130 12190 15140 12230
rect 15180 12190 15190 12230
rect 13680 12110 13690 12170
rect 13750 12110 13760 12170
rect 13680 12100 13760 12110
rect 13940 12030 13980 12170
rect 14010 12122 14068 12130
rect 14010 12070 14012 12122
rect 14064 12070 14068 12122
rect 14010 12060 14068 12070
rect 13920 12020 14000 12030
rect 13920 11960 13930 12020
rect 13990 11960 14000 12020
rect 13920 11950 14000 11960
rect 14180 11920 14220 12170
rect 14334 12122 14392 12130
rect 14334 12070 14336 12122
rect 14388 12070 14392 12122
rect 14334 12060 14392 12070
rect 14420 12030 14460 12170
rect 14488 12122 14546 12130
rect 14488 12070 14490 12122
rect 14542 12070 14546 12122
rect 14488 12060 14546 12070
rect 14400 12020 14480 12030
rect 14400 11960 14410 12020
rect 14470 11960 14480 12020
rect 14400 11950 14480 11960
rect 14660 11920 14700 12170
rect 14812 12122 14870 12130
rect 14812 12070 14814 12122
rect 14866 12070 14870 12122
rect 14812 12060 14870 12070
rect 14900 12030 14940 12170
rect 14970 12122 15028 12130
rect 14970 12070 14972 12122
rect 15024 12070 15028 12122
rect 14970 12060 15028 12070
rect 14880 12020 14960 12030
rect 14880 11960 14890 12020
rect 14950 11960 14960 12020
rect 14160 11910 14240 11920
rect 14160 11850 14170 11910
rect 14230 11850 14240 11910
rect 14160 11840 14240 11850
rect 14640 11910 14720 11920
rect 14640 11850 14650 11910
rect 14710 11850 14720 11910
rect 14640 11840 14720 11850
rect 13740 11800 13820 11810
rect 13740 11740 13750 11800
rect 13810 11740 13820 11800
rect 13740 11720 13820 11740
rect 13740 11660 13750 11720
rect 13810 11660 13820 11720
rect 13740 11640 13820 11660
rect 13740 11580 13750 11640
rect 13810 11580 13820 11640
rect 13740 11570 13820 11580
rect 13920 11800 14000 11810
rect 13920 11740 13930 11800
rect 13990 11740 14000 11800
rect 13920 11720 14000 11740
rect 13920 11660 13930 11720
rect 13990 11660 14000 11720
rect 13920 11640 14000 11660
rect 13920 11580 13930 11640
rect 13990 11580 14000 11640
rect 13920 11570 14000 11580
rect 14160 11800 14240 11810
rect 14160 11740 14170 11800
rect 14230 11740 14240 11800
rect 14160 11720 14240 11740
rect 14160 11660 14170 11720
rect 14230 11660 14240 11720
rect 14160 11640 14240 11660
rect 14160 11580 14170 11640
rect 14230 11580 14240 11640
rect 14160 11570 14240 11580
rect 14400 11800 14480 11810
rect 14400 11740 14410 11800
rect 14470 11740 14480 11800
rect 14400 11720 14480 11740
rect 14400 11660 14410 11720
rect 14470 11660 14480 11720
rect 14400 11640 14480 11660
rect 14400 11580 14410 11640
rect 14470 11580 14480 11640
rect 14400 11570 14480 11580
rect 14640 11800 14720 11810
rect 14640 11740 14650 11800
rect 14710 11740 14720 11800
rect 14640 11720 14720 11740
rect 14640 11660 14650 11720
rect 14710 11660 14720 11720
rect 14640 11640 14720 11660
rect 14640 11580 14650 11640
rect 14710 11580 14720 11640
rect 14640 11570 14720 11580
rect 13750 11510 13810 11570
rect 13750 11470 13760 11510
rect 13800 11470 13810 11510
rect 13750 11450 13810 11470
rect 13570 11390 13630 11410
rect 13570 11350 13580 11390
rect 13620 11350 13630 11390
rect 13570 11290 13630 11350
rect 13570 11250 13580 11290
rect 13620 11250 13630 11290
rect 12930 11130 12940 11170
rect 12980 11130 12990 11170
rect 12930 11080 12990 11130
rect 13060 11180 13140 11190
rect 13060 11120 13070 11180
rect 13130 11120 13140 11180
rect 13060 11110 13140 11120
rect 13420 11180 13500 11190
rect 13420 11120 13430 11180
rect 13490 11120 13500 11180
rect 10520 11070 10600 11080
rect 10520 11010 10530 11070
rect 10590 11010 10600 11070
rect 10520 10990 10600 11010
rect 10520 10930 10530 10990
rect 10590 10930 10600 10990
rect 10520 10910 10600 10930
rect 10520 10850 10530 10910
rect 10590 10850 10600 10910
rect 10520 10840 10600 10850
rect 10760 11070 10840 11080
rect 10760 11010 10770 11070
rect 10830 11010 10840 11070
rect 10760 10990 10840 11010
rect 10760 10930 10770 10990
rect 10830 10930 10840 10990
rect 10760 10910 10840 10930
rect 10760 10850 10770 10910
rect 10830 10850 10840 10910
rect 10760 10840 10840 10850
rect 11000 11070 11080 11080
rect 11000 11010 11010 11070
rect 11070 11010 11080 11070
rect 11000 10990 11080 11010
rect 11000 10930 11010 10990
rect 11070 10930 11080 10990
rect 11000 10910 11080 10930
rect 11000 10850 11010 10910
rect 11070 10850 11080 10910
rect 11000 10840 11080 10850
rect 11240 11070 11320 11080
rect 11240 11010 11250 11070
rect 11310 11010 11320 11070
rect 11240 10990 11320 11010
rect 11240 10930 11250 10990
rect 11310 10930 11320 10990
rect 11240 10910 11320 10930
rect 11240 10850 11250 10910
rect 11310 10850 11320 10910
rect 11240 10840 11320 10850
rect 11480 11070 11560 11080
rect 11480 11010 11490 11070
rect 11550 11010 11560 11070
rect 11480 10990 11560 11010
rect 11480 10930 11490 10990
rect 11550 10930 11560 10990
rect 11480 10910 11560 10930
rect 11480 10850 11490 10910
rect 11550 10850 11560 10910
rect 11480 10840 11560 10850
rect 11720 11070 11800 11080
rect 11720 11010 11730 11070
rect 11790 11010 11800 11070
rect 11720 10990 11800 11010
rect 11720 10930 11730 10990
rect 11790 10930 11800 10990
rect 11720 10910 11800 10930
rect 11720 10850 11730 10910
rect 11790 10850 11800 10910
rect 11720 10840 11800 10850
rect 11960 11070 12040 11080
rect 11960 11010 11970 11070
rect 12030 11010 12040 11070
rect 11960 10990 12040 11010
rect 11960 10930 11970 10990
rect 12030 10930 12040 10990
rect 11960 10910 12040 10930
rect 11960 10850 11970 10910
rect 12030 10850 12040 10910
rect 11960 10840 12040 10850
rect 12200 11070 12280 11080
rect 12200 11010 12210 11070
rect 12270 11010 12280 11070
rect 12200 10990 12280 11010
rect 12200 10930 12210 10990
rect 12270 10930 12280 10990
rect 12200 10910 12280 10930
rect 12200 10850 12210 10910
rect 12270 10850 12280 10910
rect 12200 10840 12280 10850
rect 12440 11070 12520 11080
rect 12440 11010 12450 11070
rect 12510 11010 12520 11070
rect 12440 10990 12520 11010
rect 12440 10930 12450 10990
rect 12510 10930 12520 10990
rect 12440 10910 12520 10930
rect 12440 10850 12450 10910
rect 12510 10850 12520 10910
rect 12440 10840 12520 10850
rect 12680 11070 12760 11080
rect 12680 11010 12690 11070
rect 12750 11010 12760 11070
rect 12680 10990 12760 11010
rect 12680 10930 12690 10990
rect 12750 10930 12760 10990
rect 12680 10910 12760 10930
rect 12680 10850 12690 10910
rect 12750 10850 12760 10910
rect 12680 10840 12760 10850
rect 12920 11070 13000 11080
rect 12920 11010 12930 11070
rect 12990 11010 13000 11070
rect 12920 10990 13000 11010
rect 12920 10930 12930 10990
rect 12990 10930 13000 10990
rect 12920 10910 13000 10930
rect 12920 10850 12930 10910
rect 12990 10850 13000 10910
rect 12920 10840 13000 10850
rect 11800 10800 11880 10810
rect 11800 10740 11810 10800
rect 11870 10740 11880 10800
rect 11800 10730 11880 10740
rect 13240 10800 13320 10810
rect 13240 10740 13250 10800
rect 13310 10740 13320 10800
rect 13240 10730 13320 10740
rect 11630 10230 11690 10250
rect 11630 10190 11640 10230
rect 11680 10190 11690 10230
rect 11630 10130 11690 10190
rect 11630 10090 11640 10130
rect 11680 10090 11690 10130
rect 11630 10030 11690 10090
rect 11630 9990 11640 10030
rect 11680 9990 11690 10030
rect 11630 9930 11690 9990
rect 11630 9890 11640 9930
rect 11680 9890 11690 9930
rect 11630 9830 11690 9890
rect 11630 9790 11640 9830
rect 11680 9790 11690 9830
rect 11630 9730 11690 9790
rect 11630 9690 11640 9730
rect 11680 9690 11690 9730
rect 11630 9670 11690 9690
rect 11810 10230 11870 10730
rect 12160 10690 12240 10700
rect 12160 10630 12170 10690
rect 12230 10630 12240 10690
rect 12160 10620 12240 10630
rect 11900 10360 11970 10370
rect 11960 10300 11970 10360
rect 11900 10290 11970 10300
rect 12070 10360 12150 10370
rect 12070 10300 12080 10360
rect 12140 10300 12150 10360
rect 12070 10290 12150 10300
rect 12180 10250 12220 10620
rect 12520 10580 12600 10590
rect 12520 10520 12530 10580
rect 12590 10520 12600 10580
rect 12520 10510 12600 10520
rect 12250 10360 12330 10370
rect 12250 10300 12260 10360
rect 12320 10300 12330 10360
rect 12250 10290 12330 10300
rect 12430 10360 12510 10370
rect 12430 10300 12440 10360
rect 12500 10300 12510 10360
rect 12430 10290 12510 10300
rect 12540 10250 12580 10510
rect 12880 10470 12960 10480
rect 12880 10410 12890 10470
rect 12950 10410 12960 10470
rect 12880 10400 12960 10410
rect 12610 10360 12690 10370
rect 12610 10300 12620 10360
rect 12680 10300 12690 10360
rect 12610 10290 12690 10300
rect 12790 10360 12870 10370
rect 12790 10300 12800 10360
rect 12860 10300 12870 10360
rect 12790 10290 12870 10300
rect 12900 10250 12940 10400
rect 12970 10360 13050 10370
rect 12970 10300 12980 10360
rect 13040 10300 13050 10360
rect 12970 10290 13050 10300
rect 13150 10360 13220 10370
rect 13150 10300 13160 10360
rect 13150 10290 13220 10300
rect 11810 10190 11820 10230
rect 11860 10190 11870 10230
rect 11810 10130 11870 10190
rect 11810 10090 11820 10130
rect 11860 10090 11870 10130
rect 11810 10030 11870 10090
rect 11810 9990 11820 10030
rect 11860 9990 11870 10030
rect 11810 9930 11870 9990
rect 11810 9890 11820 9930
rect 11860 9890 11870 9930
rect 11810 9830 11870 9890
rect 11810 9790 11820 9830
rect 11860 9790 11870 9830
rect 11810 9730 11870 9790
rect 11810 9690 11820 9730
rect 11860 9690 11870 9730
rect 11810 9670 11870 9690
rect 11990 10230 12050 10250
rect 11990 10190 12000 10230
rect 12040 10190 12050 10230
rect 11990 10130 12050 10190
rect 11990 10090 12000 10130
rect 12040 10090 12050 10130
rect 11990 10030 12050 10090
rect 11990 9990 12000 10030
rect 12040 9990 12050 10030
rect 11990 9930 12050 9990
rect 11990 9890 12000 9930
rect 12040 9890 12050 9930
rect 11990 9830 12050 9890
rect 11990 9790 12000 9830
rect 12040 9790 12050 9830
rect 11990 9730 12050 9790
rect 11990 9690 12000 9730
rect 12040 9690 12050 9730
rect 11990 9670 12050 9690
rect 12170 10230 12230 10250
rect 12170 10190 12180 10230
rect 12220 10190 12230 10230
rect 12170 10130 12230 10190
rect 12170 10090 12180 10130
rect 12220 10090 12230 10130
rect 12170 10030 12230 10090
rect 12170 9990 12180 10030
rect 12220 9990 12230 10030
rect 12170 9930 12230 9990
rect 12170 9890 12180 9930
rect 12220 9890 12230 9930
rect 12170 9830 12230 9890
rect 12170 9790 12180 9830
rect 12220 9790 12230 9830
rect 12170 9730 12230 9790
rect 12170 9690 12180 9730
rect 12220 9690 12230 9730
rect 12170 9670 12230 9690
rect 12350 10230 12410 10250
rect 12350 10190 12360 10230
rect 12400 10190 12410 10230
rect 12350 10130 12410 10190
rect 12350 10090 12360 10130
rect 12400 10090 12410 10130
rect 12350 10030 12410 10090
rect 12350 9990 12360 10030
rect 12400 9990 12410 10030
rect 12350 9930 12410 9990
rect 12350 9890 12360 9930
rect 12400 9890 12410 9930
rect 12350 9830 12410 9890
rect 12350 9790 12360 9830
rect 12400 9790 12410 9830
rect 12350 9730 12410 9790
rect 12350 9690 12360 9730
rect 12400 9690 12410 9730
rect 12350 9670 12410 9690
rect 12530 10230 12590 10250
rect 12530 10190 12540 10230
rect 12580 10190 12590 10230
rect 12530 10130 12590 10190
rect 12530 10090 12540 10130
rect 12580 10090 12590 10130
rect 12530 10030 12590 10090
rect 12530 9990 12540 10030
rect 12580 9990 12590 10030
rect 12530 9930 12590 9990
rect 12530 9890 12540 9930
rect 12580 9890 12590 9930
rect 12530 9830 12590 9890
rect 12530 9790 12540 9830
rect 12580 9790 12590 9830
rect 12530 9730 12590 9790
rect 12530 9690 12540 9730
rect 12580 9690 12590 9730
rect 12530 9670 12590 9690
rect 12710 10230 12770 10250
rect 12710 10190 12720 10230
rect 12760 10190 12770 10230
rect 12710 10130 12770 10190
rect 12710 10090 12720 10130
rect 12760 10090 12770 10130
rect 12710 10030 12770 10090
rect 12710 9990 12720 10030
rect 12760 9990 12770 10030
rect 12710 9930 12770 9990
rect 12710 9890 12720 9930
rect 12760 9890 12770 9930
rect 12710 9830 12770 9890
rect 12710 9790 12720 9830
rect 12760 9790 12770 9830
rect 12710 9730 12770 9790
rect 12710 9690 12720 9730
rect 12760 9690 12770 9730
rect 12710 9670 12770 9690
rect 12890 10230 12950 10250
rect 12890 10190 12900 10230
rect 12940 10190 12950 10230
rect 12890 10130 12950 10190
rect 12890 10090 12900 10130
rect 12940 10090 12950 10130
rect 12890 10030 12950 10090
rect 12890 9990 12900 10030
rect 12940 9990 12950 10030
rect 12890 9930 12950 9990
rect 12890 9890 12900 9930
rect 12940 9890 12950 9930
rect 12890 9830 12950 9890
rect 12890 9790 12900 9830
rect 12940 9790 12950 9830
rect 12890 9730 12950 9790
rect 12890 9690 12900 9730
rect 12940 9690 12950 9730
rect 12890 9670 12950 9690
rect 13070 10230 13130 10250
rect 13070 10190 13080 10230
rect 13120 10190 13130 10230
rect 13070 10130 13130 10190
rect 13070 10090 13080 10130
rect 13120 10090 13130 10130
rect 13070 10030 13130 10090
rect 13070 9990 13080 10030
rect 13120 9990 13130 10030
rect 13070 9930 13130 9990
rect 13070 9890 13080 9930
rect 13120 9890 13130 9930
rect 13070 9830 13130 9890
rect 13070 9790 13080 9830
rect 13120 9790 13130 9830
rect 13070 9730 13130 9790
rect 13070 9690 13080 9730
rect 13120 9690 13130 9730
rect 13070 9670 13130 9690
rect 13250 10230 13310 10730
rect 13420 10370 13500 11120
rect 13570 11170 13630 11250
rect 13690 11390 13750 11410
rect 13690 11350 13700 11390
rect 13740 11350 13750 11390
rect 13690 11290 13750 11350
rect 13690 11250 13700 11290
rect 13740 11250 13750 11290
rect 13690 11190 13750 11250
rect 13810 11390 13870 11410
rect 13810 11350 13820 11390
rect 13860 11350 13870 11390
rect 13810 11290 13870 11350
rect 13810 11250 13820 11290
rect 13860 11250 13870 11290
rect 13570 11130 13580 11170
rect 13620 11130 13630 11170
rect 13570 11080 13630 11130
rect 13680 11180 13760 11190
rect 13680 11120 13690 11180
rect 13750 11120 13760 11180
rect 13680 11110 13760 11120
rect 13810 11080 13870 11250
rect 13930 11390 13990 11570
rect 14160 11520 14240 11530
rect 14160 11460 14170 11520
rect 14230 11460 14240 11520
rect 14160 11450 14240 11460
rect 14410 11510 14470 11570
rect 14410 11470 14420 11510
rect 14460 11470 14470 11510
rect 14410 11450 14470 11470
rect 13930 11350 13940 11390
rect 13980 11350 13990 11390
rect 13930 11290 13990 11350
rect 13930 11250 13940 11290
rect 13980 11250 13990 11290
rect 13930 11230 13990 11250
rect 14050 11390 14110 11410
rect 14050 11350 14060 11390
rect 14100 11350 14110 11390
rect 14050 11290 14110 11350
rect 14050 11250 14060 11290
rect 14100 11250 14110 11290
rect 14050 11080 14110 11250
rect 14170 11390 14230 11450
rect 14170 11350 14180 11390
rect 14220 11350 14230 11390
rect 14170 11290 14230 11350
rect 14170 11250 14180 11290
rect 14220 11250 14230 11290
rect 14170 11230 14230 11250
rect 14290 11390 14350 11410
rect 14290 11350 14300 11390
rect 14340 11350 14350 11390
rect 14290 11290 14350 11350
rect 14290 11250 14300 11290
rect 14340 11250 14350 11290
rect 14290 11080 14350 11250
rect 14410 11390 14470 11410
rect 14410 11350 14420 11390
rect 14460 11350 14470 11390
rect 14410 11290 14470 11350
rect 14410 11250 14420 11290
rect 14460 11250 14470 11290
rect 14410 11190 14470 11250
rect 14530 11390 14590 11410
rect 14530 11350 14540 11390
rect 14580 11350 14590 11390
rect 14530 11290 14590 11350
rect 14530 11250 14540 11290
rect 14580 11250 14590 11290
rect 14400 11180 14480 11190
rect 14400 11120 14410 11180
rect 14470 11120 14480 11180
rect 14400 11110 14480 11120
rect 14530 11080 14590 11250
rect 14650 11390 14710 11570
rect 14880 11520 14960 11960
rect 15130 11920 15190 12190
rect 15120 11910 15200 11920
rect 15120 11850 15130 11910
rect 15190 11850 15200 11910
rect 15120 11800 15200 11850
rect 15120 11740 15130 11800
rect 15190 11740 15200 11800
rect 15120 11720 15200 11740
rect 15120 11660 15130 11720
rect 15190 11660 15200 11720
rect 15120 11640 15200 11660
rect 15120 11580 15130 11640
rect 15190 11580 15200 11640
rect 15120 11570 15200 11580
rect 15360 11800 15440 11810
rect 15360 11740 15370 11800
rect 15430 11740 15440 11800
rect 15360 11720 15440 11740
rect 15360 11660 15370 11720
rect 15430 11660 15440 11720
rect 15360 11640 15440 11660
rect 15360 11580 15370 11640
rect 15430 11580 15440 11640
rect 15360 11570 15440 11580
rect 15780 11800 15860 11810
rect 15780 11740 15790 11800
rect 15850 11740 15860 11800
rect 15780 11720 15860 11740
rect 15780 11660 15790 11720
rect 15850 11660 15860 11720
rect 15780 11640 15860 11660
rect 15780 11580 15790 11640
rect 15850 11580 15860 11640
rect 15780 11570 15860 11580
rect 14880 11460 14890 11520
rect 14950 11460 14960 11520
rect 14880 11450 14960 11460
rect 15130 11510 15190 11570
rect 15130 11470 15140 11510
rect 15180 11470 15190 11510
rect 15130 11450 15190 11470
rect 14650 11350 14660 11390
rect 14700 11350 14710 11390
rect 14650 11290 14710 11350
rect 14650 11250 14660 11290
rect 14700 11250 14710 11290
rect 14650 11230 14710 11250
rect 14770 11390 14830 11410
rect 14770 11350 14780 11390
rect 14820 11350 14830 11390
rect 14770 11290 14830 11350
rect 14770 11250 14780 11290
rect 14820 11250 14830 11290
rect 14770 11080 14830 11250
rect 14890 11390 14950 11450
rect 14890 11350 14900 11390
rect 14940 11350 14950 11390
rect 14890 11290 14950 11350
rect 14890 11250 14900 11290
rect 14940 11250 14950 11290
rect 14890 11230 14950 11250
rect 15010 11390 15070 11410
rect 15010 11350 15020 11390
rect 15060 11350 15070 11390
rect 15010 11290 15070 11350
rect 15010 11250 15020 11290
rect 15060 11250 15070 11290
rect 15010 11080 15070 11250
rect 15130 11390 15190 11410
rect 15130 11350 15140 11390
rect 15180 11350 15190 11390
rect 15130 11290 15190 11350
rect 15130 11250 15140 11290
rect 15180 11250 15190 11290
rect 15130 11190 15190 11250
rect 15250 11390 15310 11410
rect 15250 11350 15260 11390
rect 15300 11350 15310 11390
rect 15250 11290 15310 11350
rect 15250 11250 15260 11290
rect 15300 11250 15310 11290
rect 15120 11180 15200 11190
rect 15120 11120 15130 11180
rect 15190 11120 15200 11180
rect 15120 11110 15200 11120
rect 15250 11080 15310 11250
rect 15370 11390 15430 11570
rect 15600 11520 15680 11530
rect 15600 11460 15610 11520
rect 15670 11460 15680 11520
rect 15790 11520 15850 11570
rect 15790 11480 15800 11520
rect 15840 11480 15850 11520
rect 15790 11460 15850 11480
rect 15600 11450 15680 11460
rect 15370 11350 15380 11390
rect 15420 11350 15430 11390
rect 15370 11290 15430 11350
rect 15370 11250 15380 11290
rect 15420 11250 15430 11290
rect 15370 11230 15430 11250
rect 15490 11390 15550 11410
rect 15490 11350 15500 11390
rect 15540 11350 15550 11390
rect 15490 11290 15550 11350
rect 15490 11250 15500 11290
rect 15540 11250 15550 11290
rect 15490 11080 15550 11250
rect 15610 11390 15670 11450
rect 15610 11350 15620 11390
rect 15660 11350 15670 11390
rect 15610 11290 15670 11350
rect 15610 11250 15620 11290
rect 15660 11250 15670 11290
rect 15610 11230 15670 11250
rect 15730 11390 15790 11410
rect 15730 11350 15740 11390
rect 15780 11350 15790 11390
rect 15730 11290 15790 11350
rect 15730 11250 15740 11290
rect 15780 11250 15790 11290
rect 15730 11080 15790 11250
rect 15850 11390 15910 11410
rect 15850 11350 15860 11390
rect 15900 11350 15910 11390
rect 15850 11290 15910 11350
rect 15850 11250 15860 11290
rect 15900 11250 15910 11290
rect 15850 11190 15910 11250
rect 15970 11390 16030 11410
rect 15970 11350 15980 11390
rect 16020 11350 16030 11390
rect 15970 11290 16030 11350
rect 15970 11250 15980 11290
rect 16020 11250 16030 11290
rect 15840 11180 15920 11190
rect 15840 11120 15850 11180
rect 15910 11120 15920 11180
rect 13560 11070 13640 11080
rect 13560 11010 13570 11070
rect 13630 11010 13640 11070
rect 13560 10990 13640 11010
rect 13560 10930 13570 10990
rect 13630 10930 13640 10990
rect 13560 10910 13640 10930
rect 13560 10850 13570 10910
rect 13630 10850 13640 10910
rect 13560 10840 13640 10850
rect 13800 11070 13880 11080
rect 13800 11010 13810 11070
rect 13870 11010 13880 11070
rect 13800 10990 13880 11010
rect 13800 10930 13810 10990
rect 13870 10930 13880 10990
rect 13800 10910 13880 10930
rect 13800 10850 13810 10910
rect 13870 10850 13880 10910
rect 13800 10840 13880 10850
rect 14040 11070 14120 11080
rect 14040 11010 14050 11070
rect 14110 11010 14120 11070
rect 14040 10990 14120 11010
rect 14040 10930 14050 10990
rect 14110 10930 14120 10990
rect 14040 10910 14120 10930
rect 14040 10850 14050 10910
rect 14110 10850 14120 10910
rect 14040 10840 14120 10850
rect 14280 11070 14360 11080
rect 14280 11010 14290 11070
rect 14350 11010 14360 11070
rect 14280 10990 14360 11010
rect 14280 10930 14290 10990
rect 14350 10930 14360 10990
rect 14280 10910 14360 10930
rect 14280 10850 14290 10910
rect 14350 10850 14360 10910
rect 14280 10840 14360 10850
rect 14520 11070 14600 11080
rect 14520 11010 14530 11070
rect 14590 11010 14600 11070
rect 14520 10990 14600 11010
rect 14520 10930 14530 10990
rect 14590 10930 14600 10990
rect 14520 10910 14600 10930
rect 14520 10850 14530 10910
rect 14590 10850 14600 10910
rect 14520 10840 14600 10850
rect 14760 11070 14840 11080
rect 14760 11010 14770 11070
rect 14830 11010 14840 11070
rect 14760 10990 14840 11010
rect 14760 10930 14770 10990
rect 14830 10930 14840 10990
rect 14760 10910 14840 10930
rect 14760 10850 14770 10910
rect 14830 10850 14840 10910
rect 14760 10840 14840 10850
rect 15000 11070 15080 11080
rect 15000 11010 15010 11070
rect 15070 11010 15080 11070
rect 15000 10990 15080 11010
rect 15000 10930 15010 10990
rect 15070 10930 15080 10990
rect 15000 10910 15080 10930
rect 15000 10850 15010 10910
rect 15070 10850 15080 10910
rect 15000 10840 15080 10850
rect 15240 11070 15320 11080
rect 15240 11010 15250 11070
rect 15310 11010 15320 11070
rect 15240 10990 15320 11010
rect 15240 10930 15250 10990
rect 15310 10930 15320 10990
rect 15240 10910 15320 10930
rect 15240 10850 15250 10910
rect 15310 10850 15320 10910
rect 15240 10840 15320 10850
rect 15480 11070 15560 11080
rect 15480 11010 15490 11070
rect 15550 11010 15560 11070
rect 15480 10990 15560 11010
rect 15480 10930 15490 10990
rect 15550 10930 15560 10990
rect 15480 10910 15560 10930
rect 15480 10850 15490 10910
rect 15550 10850 15560 10910
rect 15480 10840 15560 10850
rect 15720 11070 15800 11080
rect 15720 11010 15730 11070
rect 15790 11010 15800 11070
rect 15720 10990 15800 11010
rect 15720 10930 15730 10990
rect 15790 10930 15800 10990
rect 15720 10910 15800 10930
rect 15720 10850 15730 10910
rect 15790 10850 15800 10910
rect 15720 10840 15800 10850
rect 14680 10800 14760 10810
rect 14680 10740 14690 10800
rect 14750 10740 14760 10800
rect 14680 10730 14760 10740
rect 14320 10690 14400 10700
rect 14320 10630 14330 10690
rect 14390 10630 14400 10690
rect 14320 10620 14400 10630
rect 13960 10580 14040 10590
rect 13960 10520 13970 10580
rect 14030 10520 14040 10580
rect 13960 10510 14040 10520
rect 13600 10470 13680 10480
rect 13600 10410 13610 10470
rect 13670 10410 13680 10470
rect 13600 10400 13680 10410
rect 13340 10360 13590 10370
rect 13400 10300 13430 10360
rect 13490 10300 13520 10360
rect 13580 10300 13590 10360
rect 13340 10290 13590 10300
rect 13620 10250 13660 10400
rect 13690 10360 13770 10370
rect 13690 10300 13700 10360
rect 13760 10300 13770 10360
rect 13690 10290 13770 10300
rect 13870 10360 13950 10370
rect 13870 10300 13880 10360
rect 13940 10300 13950 10360
rect 13870 10290 13950 10300
rect 13980 10250 14020 10510
rect 14050 10360 14130 10370
rect 14050 10300 14060 10360
rect 14120 10300 14130 10360
rect 14050 10290 14130 10300
rect 14230 10360 14310 10370
rect 14230 10300 14240 10360
rect 14300 10300 14310 10360
rect 14230 10290 14310 10300
rect 14340 10250 14380 10620
rect 14410 10360 14490 10370
rect 14410 10300 14420 10360
rect 14480 10300 14490 10360
rect 14410 10290 14490 10300
rect 14590 10360 14660 10370
rect 14590 10300 14600 10360
rect 14590 10290 14660 10300
rect 13250 10190 13260 10230
rect 13300 10190 13310 10230
rect 13250 10130 13310 10190
rect 13250 10090 13260 10130
rect 13300 10090 13310 10130
rect 13250 10030 13310 10090
rect 13250 9990 13260 10030
rect 13300 9990 13310 10030
rect 13250 9930 13310 9990
rect 13250 9890 13260 9930
rect 13300 9890 13310 9930
rect 13250 9830 13310 9890
rect 13250 9790 13260 9830
rect 13300 9790 13310 9830
rect 13250 9730 13310 9790
rect 13250 9690 13260 9730
rect 13300 9690 13310 9730
rect 13250 9670 13310 9690
rect 13430 10230 13490 10250
rect 13430 10190 13440 10230
rect 13480 10190 13490 10230
rect 13430 10130 13490 10190
rect 13430 10090 13440 10130
rect 13480 10090 13490 10130
rect 13430 10030 13490 10090
rect 13430 9990 13440 10030
rect 13480 9990 13490 10030
rect 13430 9930 13490 9990
rect 13430 9890 13440 9930
rect 13480 9890 13490 9930
rect 13430 9830 13490 9890
rect 13430 9790 13440 9830
rect 13480 9790 13490 9830
rect 13430 9730 13490 9790
rect 13430 9690 13440 9730
rect 13480 9690 13490 9730
rect 13430 9670 13490 9690
rect 13610 10230 13670 10250
rect 13610 10190 13620 10230
rect 13660 10190 13670 10230
rect 13610 10130 13670 10190
rect 13610 10090 13620 10130
rect 13660 10090 13670 10130
rect 13610 10030 13670 10090
rect 13610 9990 13620 10030
rect 13660 9990 13670 10030
rect 13610 9930 13670 9990
rect 13610 9890 13620 9930
rect 13660 9890 13670 9930
rect 13610 9830 13670 9890
rect 13610 9790 13620 9830
rect 13660 9790 13670 9830
rect 13610 9730 13670 9790
rect 13610 9690 13620 9730
rect 13660 9690 13670 9730
rect 13610 9670 13670 9690
rect 13790 10230 13850 10250
rect 13790 10190 13800 10230
rect 13840 10190 13850 10230
rect 13790 10130 13850 10190
rect 13790 10090 13800 10130
rect 13840 10090 13850 10130
rect 13790 10030 13850 10090
rect 13790 9990 13800 10030
rect 13840 9990 13850 10030
rect 13790 9930 13850 9990
rect 13790 9890 13800 9930
rect 13840 9890 13850 9930
rect 13790 9830 13850 9890
rect 13790 9790 13800 9830
rect 13840 9790 13850 9830
rect 13790 9730 13850 9790
rect 13790 9690 13800 9730
rect 13840 9690 13850 9730
rect 13790 9670 13850 9690
rect 13970 10230 14030 10250
rect 13970 10190 13980 10230
rect 14020 10190 14030 10230
rect 13970 10130 14030 10190
rect 13970 10090 13980 10130
rect 14020 10090 14030 10130
rect 13970 10030 14030 10090
rect 13970 9990 13980 10030
rect 14020 9990 14030 10030
rect 13970 9930 14030 9990
rect 13970 9890 13980 9930
rect 14020 9890 14030 9930
rect 13970 9830 14030 9890
rect 13970 9790 13980 9830
rect 14020 9790 14030 9830
rect 13970 9730 14030 9790
rect 13970 9690 13980 9730
rect 14020 9690 14030 9730
rect 13970 9670 14030 9690
rect 14150 10230 14210 10250
rect 14150 10190 14160 10230
rect 14200 10190 14210 10230
rect 14150 10130 14210 10190
rect 14150 10090 14160 10130
rect 14200 10090 14210 10130
rect 14150 10030 14210 10090
rect 14150 9990 14160 10030
rect 14200 9990 14210 10030
rect 14150 9930 14210 9990
rect 14150 9890 14160 9930
rect 14200 9890 14210 9930
rect 14150 9830 14210 9890
rect 14150 9790 14160 9830
rect 14200 9790 14210 9830
rect 14150 9730 14210 9790
rect 14150 9690 14160 9730
rect 14200 9690 14210 9730
rect 14150 9670 14210 9690
rect 14330 10230 14390 10250
rect 14330 10190 14340 10230
rect 14380 10190 14390 10230
rect 14330 10130 14390 10190
rect 14330 10090 14340 10130
rect 14380 10090 14390 10130
rect 14330 10030 14390 10090
rect 14330 9990 14340 10030
rect 14380 9990 14390 10030
rect 14330 9930 14390 9990
rect 14330 9890 14340 9930
rect 14380 9890 14390 9930
rect 14330 9830 14390 9890
rect 14330 9790 14340 9830
rect 14380 9790 14390 9830
rect 14330 9730 14390 9790
rect 14330 9690 14340 9730
rect 14380 9690 14390 9730
rect 14330 9670 14390 9690
rect 14510 10230 14570 10250
rect 14510 10190 14520 10230
rect 14560 10190 14570 10230
rect 14510 10130 14570 10190
rect 14510 10090 14520 10130
rect 14560 10090 14570 10130
rect 14510 10030 14570 10090
rect 14510 9990 14520 10030
rect 14560 9990 14570 10030
rect 14510 9930 14570 9990
rect 14510 9890 14520 9930
rect 14560 9890 14570 9930
rect 14510 9830 14570 9890
rect 14510 9790 14520 9830
rect 14560 9790 14570 9830
rect 14510 9730 14570 9790
rect 14510 9690 14520 9730
rect 14560 9690 14570 9730
rect 14510 9670 14570 9690
rect 14690 10230 14750 10730
rect 15710 10690 15790 10700
rect 15710 10630 15720 10690
rect 15780 10630 15790 10690
rect 15240 10580 15320 10590
rect 15240 10520 15250 10580
rect 15310 10520 15320 10580
rect 15240 10510 15320 10520
rect 14690 10190 14700 10230
rect 14740 10190 14750 10230
rect 14690 10130 14750 10190
rect 14690 10090 14700 10130
rect 14740 10090 14750 10130
rect 14690 10030 14750 10090
rect 14690 9990 14700 10030
rect 14740 9990 14750 10030
rect 14690 9930 14750 9990
rect 14690 9890 14700 9930
rect 14740 9890 14750 9930
rect 14690 9830 14750 9890
rect 14690 9790 14700 9830
rect 14740 9790 14750 9830
rect 14690 9730 14750 9790
rect 14690 9690 14700 9730
rect 14740 9690 14750 9730
rect 14690 9670 14750 9690
rect 14870 10230 14930 10250
rect 14870 10190 14880 10230
rect 14920 10190 14930 10230
rect 14870 10130 14930 10190
rect 14870 10090 14880 10130
rect 14920 10090 14930 10130
rect 14870 10030 14930 10090
rect 14870 9990 14880 10030
rect 14920 9990 14930 10030
rect 14870 9930 14930 9990
rect 14870 9890 14880 9930
rect 14920 9890 14930 9930
rect 14870 9830 14930 9890
rect 15260 9830 15300 10510
rect 15590 10160 15670 10170
rect 15590 10100 15600 10160
rect 15660 10100 15670 10160
rect 15590 10090 15670 10100
rect 15710 10150 15790 10630
rect 15840 10170 15920 11120
rect 15970 11170 16030 11250
rect 15970 11130 15980 11170
rect 16020 11130 16030 11170
rect 15970 11080 16030 11130
rect 15960 11070 16040 11080
rect 15960 11010 15970 11070
rect 16030 11010 16040 11070
rect 15960 10990 16040 11010
rect 15960 10930 15970 10990
rect 16030 10930 16040 10990
rect 15960 10910 16040 10930
rect 15960 10850 15970 10910
rect 16030 10850 16040 10910
rect 15960 10840 16040 10850
rect 16170 10480 16210 12280
rect 16260 12130 16300 14730
rect 16240 12120 16320 12130
rect 16240 12060 16250 12120
rect 16310 12060 16320 12120
rect 16240 12050 16320 12060
rect 16260 10590 16300 12050
rect 16350 11800 16590 15290
rect 16780 14090 16860 15970
rect 16780 14030 16790 14090
rect 16850 14030 16860 14090
rect 16780 14020 16860 14030
rect 16350 11740 16360 11800
rect 16420 11740 16440 11800
rect 16500 11740 16520 11800
rect 16580 11740 16590 11800
rect 16350 11720 16590 11740
rect 16350 11660 16360 11720
rect 16420 11660 16440 11720
rect 16500 11660 16520 11720
rect 16580 11660 16590 11720
rect 16350 11640 16590 11660
rect 16350 11580 16360 11640
rect 16420 11580 16440 11640
rect 16500 11580 16520 11640
rect 16580 11580 16590 11640
rect 16350 11570 16590 11580
rect 17570 11180 17650 16638
rect 17950 16050 18030 18050
rect 17950 15990 17960 16050
rect 18020 15990 18030 16050
rect 17950 15980 18030 15990
rect 18120 17450 18200 17460
rect 18120 17390 18130 17450
rect 18190 17390 18200 17450
rect 18120 13040 18200 17390
rect 18650 13980 18730 18070
rect 18780 16750 18880 16770
rect 18780 16690 18800 16750
rect 18860 16690 18880 16750
rect 18780 16670 18880 16690
rect 18780 15350 18880 15370
rect 18780 15290 18800 15350
rect 18860 15290 18880 15350
rect 18780 15270 18880 15290
rect 18650 13920 18660 13980
rect 18720 13920 18730 13980
rect 18650 13910 18730 13920
rect 17570 11120 17580 11180
rect 17640 11120 17650 11180
rect 17570 11110 17650 11120
rect 16240 10580 16320 10590
rect 16240 10520 16250 10580
rect 16310 10520 16320 10580
rect 16240 10510 16320 10520
rect 16150 10470 16230 10480
rect 16150 10410 16160 10470
rect 16220 10410 16230 10470
rect 16150 10400 16230 10410
rect 15710 10110 15730 10150
rect 15770 10110 15790 10150
rect 15710 10090 15790 10110
rect 15830 10160 15910 10170
rect 15830 10100 15840 10160
rect 15900 10100 15910 10160
rect 15830 10090 15910 10100
rect 15500 10030 15560 10050
rect 15500 9990 15510 10030
rect 15550 9990 15560 10030
rect 15500 9930 15560 9990
rect 15500 9890 15510 9930
rect 15550 9890 15560 9930
rect 15500 9830 15560 9890
rect 15610 10030 15670 10090
rect 15610 9990 15620 10030
rect 15660 9990 15670 10030
rect 15610 9930 15670 9990
rect 15610 9890 15620 9930
rect 15660 9890 15670 9930
rect 15610 9870 15670 9890
rect 15720 10030 15780 10050
rect 15720 9990 15730 10030
rect 15770 9990 15780 10030
rect 15720 9930 15780 9990
rect 15720 9890 15730 9930
rect 15770 9890 15780 9930
rect 15720 9830 15780 9890
rect 15830 10030 15890 10090
rect 15830 9990 15840 10030
rect 15880 9990 15890 10030
rect 15830 9930 15890 9990
rect 15830 9890 15840 9930
rect 15880 9890 15890 9930
rect 15830 9870 15890 9890
rect 15940 10030 16000 10050
rect 15940 9990 15950 10030
rect 15990 9990 16000 10030
rect 15940 9930 16000 9990
rect 15940 9890 15950 9930
rect 15990 9890 16000 9930
rect 15940 9830 16000 9890
rect 14870 9790 14880 9830
rect 14920 9790 14930 9830
rect 14870 9730 14930 9790
rect 15240 9820 15320 9830
rect 15240 9760 15250 9820
rect 15310 9760 15320 9820
rect 15240 9750 15320 9760
rect 15490 9810 15570 9830
rect 15490 9770 15510 9810
rect 15550 9770 15570 9810
rect 15490 9750 15570 9770
rect 15710 9820 15790 9830
rect 15710 9760 15720 9820
rect 15780 9760 15790 9820
rect 15710 9750 15790 9760
rect 15930 9810 16010 9830
rect 15930 9770 15950 9810
rect 15990 9770 16010 9810
rect 15930 9750 16010 9770
rect 14870 9690 14880 9730
rect 14920 9690 14930 9730
rect 14870 9670 14930 9690
rect 15500 9630 15560 9750
rect 15940 9630 16000 9750
rect 11620 9620 11700 9630
rect 11620 9560 11630 9620
rect 11690 9560 11700 9620
rect 11620 9540 11700 9560
rect 11620 9480 11630 9540
rect 11690 9480 11700 9540
rect 11620 9460 11700 9480
rect 11620 9400 11630 9460
rect 11690 9400 11700 9460
rect 11620 9390 11700 9400
rect 11980 9620 12060 9630
rect 11980 9560 11990 9620
rect 12050 9560 12060 9620
rect 11980 9540 12060 9560
rect 11980 9480 11990 9540
rect 12050 9480 12060 9540
rect 11980 9460 12060 9480
rect 11980 9400 11990 9460
rect 12050 9400 12060 9460
rect 11980 9390 12060 9400
rect 12340 9620 12420 9630
rect 12340 9560 12350 9620
rect 12410 9560 12420 9620
rect 12340 9540 12420 9560
rect 12340 9480 12350 9540
rect 12410 9480 12420 9540
rect 12340 9460 12420 9480
rect 12340 9400 12350 9460
rect 12410 9400 12420 9460
rect 12340 9390 12420 9400
rect 12700 9620 12780 9630
rect 12700 9560 12710 9620
rect 12770 9560 12780 9620
rect 12700 9540 12780 9560
rect 12700 9480 12710 9540
rect 12770 9480 12780 9540
rect 12700 9460 12780 9480
rect 12700 9400 12710 9460
rect 12770 9400 12780 9460
rect 12700 9390 12780 9400
rect 13060 9620 13140 9630
rect 13060 9560 13070 9620
rect 13130 9560 13140 9620
rect 13060 9540 13140 9560
rect 13060 9480 13070 9540
rect 13130 9480 13140 9540
rect 13060 9460 13140 9480
rect 13060 9400 13070 9460
rect 13130 9400 13140 9460
rect 13060 9390 13140 9400
rect 13420 9620 13500 9630
rect 13420 9560 13430 9620
rect 13490 9560 13500 9620
rect 13420 9540 13500 9560
rect 13420 9480 13430 9540
rect 13490 9480 13500 9540
rect 13420 9460 13500 9480
rect 13420 9400 13430 9460
rect 13490 9400 13500 9460
rect 13420 9390 13500 9400
rect 13780 9620 13860 9630
rect 13780 9560 13790 9620
rect 13850 9560 13860 9620
rect 13780 9540 13860 9560
rect 13780 9480 13790 9540
rect 13850 9480 13860 9540
rect 13780 9460 13860 9480
rect 13780 9400 13790 9460
rect 13850 9400 13860 9460
rect 13780 9390 13860 9400
rect 14140 9620 14220 9630
rect 14140 9560 14150 9620
rect 14210 9560 14220 9620
rect 14140 9540 14220 9560
rect 14140 9480 14150 9540
rect 14210 9480 14220 9540
rect 14140 9460 14220 9480
rect 14140 9400 14150 9460
rect 14210 9400 14220 9460
rect 14140 9390 14220 9400
rect 14500 9620 14580 9630
rect 14500 9560 14510 9620
rect 14570 9560 14580 9620
rect 14500 9540 14580 9560
rect 14500 9480 14510 9540
rect 14570 9480 14580 9540
rect 14500 9460 14580 9480
rect 14500 9400 14510 9460
rect 14570 9400 14580 9460
rect 14500 9390 14580 9400
rect 14860 9620 14940 9630
rect 14860 9560 14870 9620
rect 14930 9560 14940 9620
rect 14860 9540 14940 9560
rect 14860 9480 14870 9540
rect 14930 9480 14940 9540
rect 14860 9460 14940 9480
rect 14860 9400 14870 9460
rect 14930 9400 14940 9460
rect 14860 9390 14940 9400
rect 15490 9620 15570 9630
rect 15490 9560 15500 9620
rect 15560 9560 15570 9620
rect 15490 9540 15570 9560
rect 15490 9480 15500 9540
rect 15560 9480 15570 9540
rect 15490 9460 15570 9480
rect 15490 9400 15500 9460
rect 15560 9400 15570 9460
rect 15490 9390 15570 9400
rect 15930 9620 16010 9630
rect 15930 9560 15940 9620
rect 16000 9560 16010 9620
rect 15930 9540 16010 9560
rect 15930 9480 15940 9540
rect 16000 9480 16010 9540
rect 15930 9460 16010 9480
rect 15930 9400 15940 9460
rect 16000 9400 16010 9460
rect 15930 9390 16010 9400
rect 11806 9350 11864 9360
rect 11806 9298 11808 9350
rect 11860 9298 11864 9350
rect 11806 9290 11864 9298
rect 11916 9350 11974 9360
rect 11916 9298 11918 9350
rect 11970 9298 11974 9350
rect 11916 9290 11974 9298
rect 12026 9350 12084 9360
rect 12026 9298 12028 9350
rect 12080 9298 12084 9350
rect 12026 9290 12084 9298
rect 12136 9350 12194 9360
rect 12136 9298 12138 9350
rect 12190 9298 12194 9350
rect 12136 9290 12194 9298
rect 12246 9350 12304 9360
rect 12246 9298 12248 9350
rect 12300 9298 12304 9350
rect 12246 9290 12304 9298
rect 12356 9350 12414 9360
rect 12356 9298 12358 9350
rect 12410 9298 12414 9350
rect 12356 9290 12414 9298
rect 12466 9350 12524 9360
rect 12466 9298 12468 9350
rect 12520 9298 12524 9350
rect 12466 9290 12524 9298
rect 12576 9350 12634 9360
rect 12576 9298 12578 9350
rect 12630 9298 12634 9350
rect 12576 9290 12634 9298
rect 12686 9350 12744 9360
rect 12686 9298 12688 9350
rect 12740 9298 12744 9350
rect 12686 9290 12744 9298
rect 12796 9350 12854 9360
rect 12796 9298 12798 9350
rect 12850 9298 12854 9350
rect 12796 9290 12854 9298
rect 13706 9350 13764 9360
rect 13706 9298 13708 9350
rect 13760 9298 13764 9350
rect 13706 9290 13764 9298
rect 13816 9350 13874 9360
rect 13816 9298 13818 9350
rect 13870 9298 13874 9350
rect 13816 9290 13874 9298
rect 13926 9350 13984 9360
rect 13926 9298 13928 9350
rect 13980 9298 13984 9350
rect 13926 9290 13984 9298
rect 14036 9350 14094 9360
rect 14036 9298 14038 9350
rect 14090 9298 14094 9350
rect 14036 9290 14094 9298
rect 14146 9350 14204 9360
rect 14146 9298 14148 9350
rect 14200 9298 14204 9350
rect 14146 9290 14204 9298
rect 14256 9350 14314 9360
rect 14256 9298 14258 9350
rect 14310 9298 14314 9350
rect 14256 9290 14314 9298
rect 14366 9350 14424 9360
rect 14366 9298 14368 9350
rect 14420 9298 14424 9350
rect 14366 9290 14424 9298
rect 14476 9350 14534 9360
rect 14476 9298 14478 9350
rect 14530 9298 14534 9350
rect 14476 9290 14534 9298
rect 14586 9350 14644 9360
rect 14586 9298 14588 9350
rect 14640 9298 14644 9350
rect 14586 9290 14644 9298
rect 14696 9350 14754 9360
rect 14696 9298 14698 9350
rect 14750 9298 14754 9350
rect 14696 9290 14754 9298
rect 11560 9230 11700 9250
rect 11560 9190 11570 9230
rect 11610 9190 11650 9230
rect 11690 9190 11700 9230
rect 11560 9130 11700 9190
rect 11560 9090 11570 9130
rect 11610 9090 11650 9130
rect 11690 9090 11700 9130
rect 11560 9070 11700 9090
rect 11640 9030 11700 9070
rect 11750 9230 11810 9250
rect 11750 9190 11760 9230
rect 11800 9190 11810 9230
rect 11750 9130 11810 9190
rect 11750 9090 11760 9130
rect 11800 9090 11810 9130
rect 11630 9020 11710 9030
rect 11630 8960 11640 9020
rect 11700 8960 11710 9020
rect 11630 8950 11710 8960
rect 11750 8920 11810 9090
rect 11860 9230 11920 9250
rect 11860 9190 11870 9230
rect 11910 9190 11920 9230
rect 11860 9130 11920 9190
rect 11860 9090 11870 9130
rect 11910 9090 11920 9130
rect 11860 9030 11920 9090
rect 11970 9230 12030 9250
rect 11970 9190 11980 9230
rect 12020 9190 12030 9230
rect 11970 9130 12030 9190
rect 11970 9090 11980 9130
rect 12020 9090 12030 9130
rect 11850 9020 11930 9030
rect 11850 8960 11860 9020
rect 11920 8960 11930 9020
rect 11850 8950 11930 8960
rect 11970 8920 12030 9090
rect 12080 9230 12140 9250
rect 12080 9190 12090 9230
rect 12130 9190 12140 9230
rect 12080 9130 12140 9190
rect 12080 9090 12090 9130
rect 12130 9090 12140 9130
rect 12080 9030 12140 9090
rect 12190 9230 12250 9250
rect 12190 9190 12200 9230
rect 12240 9190 12250 9230
rect 12190 9130 12250 9190
rect 12190 9090 12200 9130
rect 12240 9090 12250 9130
rect 12070 9020 12150 9030
rect 12070 8960 12080 9020
rect 12140 8960 12150 9020
rect 12070 8950 12150 8960
rect 12190 8920 12250 9090
rect 12300 9230 12360 9250
rect 12300 9190 12310 9230
rect 12350 9190 12360 9230
rect 12300 9130 12360 9190
rect 12300 9090 12310 9130
rect 12350 9090 12360 9130
rect 12300 9030 12360 9090
rect 12410 9230 12470 9250
rect 12410 9190 12420 9230
rect 12460 9190 12470 9230
rect 12410 9130 12470 9190
rect 12410 9090 12420 9130
rect 12460 9090 12470 9130
rect 12290 9020 12370 9030
rect 12290 8960 12300 9020
rect 12360 8960 12370 9020
rect 12290 8950 12370 8960
rect 12410 8920 12470 9090
rect 12520 9230 12580 9250
rect 12520 9190 12530 9230
rect 12570 9190 12580 9230
rect 12520 9130 12580 9190
rect 12520 9090 12530 9130
rect 12570 9090 12580 9130
rect 12520 9030 12580 9090
rect 12630 9230 12690 9250
rect 12630 9190 12640 9230
rect 12680 9190 12690 9230
rect 12630 9130 12690 9190
rect 12630 9090 12640 9130
rect 12680 9090 12690 9130
rect 12510 9020 12590 9030
rect 12510 8960 12520 9020
rect 12580 8960 12590 9020
rect 12510 8950 12590 8960
rect 12630 8920 12690 9090
rect 12740 9230 12800 9250
rect 12740 9190 12750 9230
rect 12790 9190 12800 9230
rect 12740 9130 12800 9190
rect 12740 9090 12750 9130
rect 12790 9090 12800 9130
rect 12740 9030 12800 9090
rect 12850 9230 12910 9250
rect 12850 9190 12860 9230
rect 12900 9190 12910 9230
rect 12850 9130 12910 9190
rect 12850 9090 12860 9130
rect 12900 9090 12910 9130
rect 12730 9020 12810 9030
rect 12730 8960 12740 9020
rect 12800 8960 12810 9020
rect 12730 8950 12810 8960
rect 12850 8920 12910 9090
rect 12960 9230 13100 9250
rect 12960 9190 12970 9230
rect 13010 9190 13050 9230
rect 13090 9190 13100 9230
rect 12960 9130 13100 9190
rect 12960 9090 12970 9130
rect 13010 9090 13050 9130
rect 13090 9090 13100 9130
rect 12960 9070 13100 9090
rect 13460 9230 13600 9250
rect 13460 9190 13470 9230
rect 13510 9190 13550 9230
rect 13590 9190 13600 9230
rect 13460 9130 13600 9190
rect 13460 9090 13470 9130
rect 13510 9090 13550 9130
rect 13590 9090 13600 9130
rect 13460 9070 13600 9090
rect 12960 9030 13020 9070
rect 13540 9030 13600 9070
rect 13650 9230 13710 9250
rect 13650 9190 13660 9230
rect 13700 9190 13710 9230
rect 13650 9130 13710 9190
rect 13650 9090 13660 9130
rect 13700 9090 13710 9130
rect 12950 9020 13030 9030
rect 12950 8960 12960 9020
rect 13020 8960 13030 9020
rect 12950 8950 13030 8960
rect 13530 9020 13610 9030
rect 13530 8960 13540 9020
rect 13600 8960 13610 9020
rect 13530 8950 13610 8960
rect 9680 8850 9690 8910
rect 9750 8850 9760 8910
rect 9680 8840 9760 8850
rect 11740 8910 11820 8920
rect 11740 8850 11750 8910
rect 11810 8850 11820 8910
rect 11740 8840 11820 8850
rect 11960 8910 12040 8920
rect 11960 8850 11970 8910
rect 12030 8850 12040 8910
rect 11960 8840 12040 8850
rect 12180 8910 12260 8920
rect 12180 8850 12190 8910
rect 12250 8850 12260 8910
rect 12180 8840 12260 8850
rect 12400 8910 12480 8920
rect 12400 8850 12410 8910
rect 12470 8850 12480 8910
rect 12400 8840 12480 8850
rect 12620 8910 12700 8920
rect 12620 8850 12630 8910
rect 12690 8850 12700 8910
rect 12620 8840 12700 8850
rect 12840 8910 12920 8920
rect 13650 8910 13710 9090
rect 13760 9230 13820 9250
rect 13760 9190 13770 9230
rect 13810 9190 13820 9230
rect 13760 9130 13820 9190
rect 13760 9090 13770 9130
rect 13810 9090 13820 9130
rect 13760 9030 13820 9090
rect 13870 9230 13930 9250
rect 13870 9190 13880 9230
rect 13920 9190 13930 9230
rect 13870 9130 13930 9190
rect 13870 9090 13880 9130
rect 13920 9090 13930 9130
rect 13750 9020 13830 9030
rect 13750 8960 13760 9020
rect 13820 8960 13830 9020
rect 13750 8950 13830 8960
rect 13870 8910 13930 9090
rect 13980 9230 14040 9250
rect 13980 9190 13990 9230
rect 14030 9190 14040 9230
rect 13980 9130 14040 9190
rect 13980 9090 13990 9130
rect 14030 9090 14040 9130
rect 13980 9030 14040 9090
rect 14090 9230 14150 9250
rect 14090 9190 14100 9230
rect 14140 9190 14150 9230
rect 14090 9130 14150 9190
rect 14090 9090 14100 9130
rect 14140 9090 14150 9130
rect 13970 9020 14050 9030
rect 13970 8960 13980 9020
rect 14040 8960 14050 9020
rect 13970 8950 14050 8960
rect 14090 8910 14150 9090
rect 14200 9230 14260 9250
rect 14200 9190 14210 9230
rect 14250 9190 14260 9230
rect 14200 9130 14260 9190
rect 14200 9090 14210 9130
rect 14250 9090 14260 9130
rect 14200 9030 14260 9090
rect 14310 9230 14370 9250
rect 14310 9190 14320 9230
rect 14360 9190 14370 9230
rect 14310 9130 14370 9190
rect 14310 9090 14320 9130
rect 14360 9090 14370 9130
rect 14190 9020 14270 9030
rect 14190 8960 14200 9020
rect 14260 8960 14270 9020
rect 14190 8950 14270 8960
rect 14310 8910 14370 9090
rect 14420 9230 14480 9250
rect 14420 9190 14430 9230
rect 14470 9190 14480 9230
rect 14420 9130 14480 9190
rect 14420 9090 14430 9130
rect 14470 9090 14480 9130
rect 14420 9030 14480 9090
rect 14530 9230 14590 9250
rect 14530 9190 14540 9230
rect 14580 9190 14590 9230
rect 14530 9130 14590 9190
rect 14530 9090 14540 9130
rect 14580 9090 14590 9130
rect 14410 9020 14490 9030
rect 14410 8960 14420 9020
rect 14480 8960 14490 9020
rect 14410 8950 14490 8960
rect 14530 8910 14590 9090
rect 14640 9230 14700 9250
rect 14640 9190 14650 9230
rect 14690 9190 14700 9230
rect 14640 9130 14700 9190
rect 14640 9090 14650 9130
rect 14690 9090 14700 9130
rect 14640 9030 14700 9090
rect 14750 9230 14810 9250
rect 14750 9190 14760 9230
rect 14800 9190 14810 9230
rect 14750 9130 14810 9190
rect 14750 9090 14760 9130
rect 14800 9090 14810 9130
rect 14630 9020 14710 9030
rect 14630 8960 14640 9020
rect 14700 8960 14710 9020
rect 14630 8950 14710 8960
rect 14750 8910 14810 9090
rect 14860 9230 15000 9250
rect 14860 9190 14870 9230
rect 14910 9190 14950 9230
rect 14990 9190 15000 9230
rect 14860 9130 15000 9190
rect 14860 9090 14870 9130
rect 14910 9090 14950 9130
rect 14990 9090 15000 9130
rect 14860 9070 15000 9090
rect 14860 9030 14920 9070
rect 14850 9020 14930 9030
rect 14850 8960 14860 9020
rect 14920 8960 14930 9020
rect 14850 8950 14930 8960
rect 12840 8850 12850 8910
rect 12910 8850 12920 8910
rect 12840 8840 12920 8850
rect 13640 8900 13720 8910
rect 13640 8840 13650 8900
rect 13710 8840 13720 8900
rect 13640 8820 13720 8840
rect 13640 8760 13650 8820
rect 13710 8760 13720 8820
rect 13640 8740 13720 8760
rect 13640 8680 13650 8740
rect 13710 8680 13720 8740
rect 13640 8670 13720 8680
rect 13860 8900 13940 8910
rect 13860 8840 13870 8900
rect 13930 8840 13940 8900
rect 13860 8820 13940 8840
rect 13860 8760 13870 8820
rect 13930 8760 13940 8820
rect 13860 8740 13940 8760
rect 13860 8680 13870 8740
rect 13930 8680 13940 8740
rect 13860 8670 13940 8680
rect 14080 8900 14160 8910
rect 14080 8840 14090 8900
rect 14150 8840 14160 8900
rect 14080 8820 14160 8840
rect 14080 8760 14090 8820
rect 14150 8760 14160 8820
rect 14080 8740 14160 8760
rect 14080 8680 14090 8740
rect 14150 8680 14160 8740
rect 14080 8670 14160 8680
rect 14300 8900 14380 8910
rect 14300 8840 14310 8900
rect 14370 8840 14380 8900
rect 14300 8820 14380 8840
rect 14300 8760 14310 8820
rect 14370 8760 14380 8820
rect 14300 8740 14380 8760
rect 14300 8680 14310 8740
rect 14370 8680 14380 8740
rect 14300 8670 14380 8680
rect 14520 8900 14600 8910
rect 14520 8840 14530 8900
rect 14590 8840 14600 8900
rect 14520 8820 14600 8840
rect 14520 8760 14530 8820
rect 14590 8760 14600 8820
rect 14520 8740 14600 8760
rect 14520 8680 14530 8740
rect 14590 8680 14600 8740
rect 14520 8670 14600 8680
rect 14740 8900 14820 8910
rect 14740 8840 14750 8900
rect 14810 8840 14820 8900
rect 14740 8820 14820 8840
rect 14740 8760 14750 8820
rect 14810 8760 14820 8820
rect 14740 8740 14820 8760
rect 14740 8680 14750 8740
rect 14810 8680 14820 8740
rect 14740 8670 14820 8680
<< via1 >>
rect 9180 19130 9240 19190
rect 8800 19020 8860 19080
rect 8800 18940 8860 19000
rect 8800 18860 8860 18920
rect 8790 18050 8870 18420
rect 9180 18390 9240 18450
rect 9180 18310 9240 18370
rect 9180 18220 9240 18280
rect 9180 18130 9240 18190
rect 9180 18050 9240 18110
rect 9580 19020 9640 19080
rect 9580 18940 9640 19000
rect 9580 18860 9640 18920
rect 10690 19020 10750 19080
rect 10690 18940 10750 19000
rect 10690 18860 10750 18920
rect 8800 11120 8860 11180
rect 9470 13750 9530 13810
rect 10360 14660 10420 14720
rect 9580 12060 9640 12120
rect 9580 10740 9640 10800
rect 9690 14030 9750 14090
rect 9690 12290 9750 12350
rect 9470 10630 9530 10690
rect 8800 9300 8860 9360
rect 10630 13920 10690 13980
rect 18200 19130 18260 19190
rect 13250 19070 13310 19080
rect 13250 19030 13260 19070
rect 13260 19030 13300 19070
rect 13300 19030 13310 19070
rect 13250 19020 13310 19030
rect 13250 18990 13310 19000
rect 13250 18950 13260 18990
rect 13260 18950 13300 18990
rect 13300 18950 13310 18990
rect 13250 18940 13310 18950
rect 13250 18910 13310 18920
rect 13250 18870 13260 18910
rect 13260 18870 13300 18910
rect 13300 18870 13310 18910
rect 13250 18860 13310 18870
rect 15680 19020 15740 19080
rect 15680 18940 15740 19000
rect 15680 18860 15740 18920
rect 16790 19020 16850 19080
rect 16790 18940 16850 19000
rect 16790 18860 16850 18920
rect 17580 19020 17640 19080
rect 17580 18940 17640 19000
rect 17580 18860 17640 18920
rect 18200 18790 18260 18850
rect 17570 18050 17650 18420
rect 17960 18390 18020 18450
rect 17960 18310 18020 18370
rect 17960 18220 18020 18280
rect 17960 18130 18020 18190
rect 17960 18050 18020 18110
rect 18660 18090 18720 18150
rect 11150 16750 11210 16810
rect 11580 16750 11640 16810
rect 13250 16754 13310 16810
rect 13250 16750 13254 16754
rect 13254 16750 13310 16754
rect 15350 16750 15410 16810
rect 15350 14740 15410 14800
rect 17570 16680 17650 16760
rect 16360 15290 16420 15350
rect 16440 15290 16500 15350
rect 16520 15290 16580 15350
rect 16010 14740 16070 14800
rect 16250 14740 16310 14800
rect 14590 14660 14650 14720
rect 14680 14660 14740 14720
rect 14770 14660 14830 14720
rect 14860 14660 14920 14720
rect 14950 14660 15010 14720
rect 11150 14350 11210 14410
rect 11560 14350 11960 14402
rect 14600 14398 15000 14402
rect 14600 14360 14996 14398
rect 14996 14360 15000 14398
rect 14600 14350 15000 14360
rect 16160 14350 16220 14410
rect 11040 13920 11100 13980
rect 11090 13800 11150 13810
rect 11090 13760 11100 13800
rect 11100 13760 11140 13800
rect 11140 13760 11150 13800
rect 11090 13750 11150 13760
rect 15480 13840 15540 13850
rect 15480 13800 15490 13840
rect 15490 13800 15530 13840
rect 15530 13800 15540 13840
rect 15480 13790 15540 13800
rect 15480 13760 15540 13770
rect 15480 13720 15490 13760
rect 15490 13720 15530 13760
rect 15530 13720 15540 13760
rect 15480 13710 15540 13720
rect 11170 13630 11230 13640
rect 11170 13590 11180 13630
rect 11180 13590 11220 13630
rect 11220 13590 11230 13630
rect 11170 13580 11230 13590
rect 11330 13630 11390 13640
rect 11330 13590 11340 13630
rect 11340 13590 11380 13630
rect 11380 13590 11390 13630
rect 11330 13580 11390 13590
rect 11490 13630 11550 13640
rect 11490 13590 11500 13630
rect 11500 13590 11540 13630
rect 11540 13590 11550 13630
rect 11490 13580 11550 13590
rect 11650 13630 11710 13640
rect 11650 13590 11660 13630
rect 11660 13590 11700 13630
rect 11700 13590 11710 13630
rect 11650 13580 11710 13590
rect 11810 13630 11870 13640
rect 11810 13590 11820 13630
rect 11820 13590 11860 13630
rect 11860 13590 11870 13630
rect 11810 13580 11870 13590
rect 11970 13630 12030 13640
rect 11970 13590 11980 13630
rect 11980 13590 12020 13630
rect 12020 13590 12030 13630
rect 11970 13580 12030 13590
rect 12130 13630 12190 13640
rect 12130 13590 12140 13630
rect 12140 13590 12180 13630
rect 12180 13590 12190 13630
rect 12130 13580 12190 13590
rect 12290 13630 12350 13640
rect 12290 13590 12300 13630
rect 12300 13590 12340 13630
rect 12340 13590 12350 13630
rect 12290 13580 12350 13590
rect 12450 13630 12510 13640
rect 12450 13590 12460 13630
rect 12460 13590 12500 13630
rect 12500 13590 12510 13630
rect 12450 13580 12510 13590
rect 12610 13630 12670 13640
rect 12610 13590 12620 13630
rect 12620 13590 12660 13630
rect 12660 13590 12670 13630
rect 12610 13580 12670 13590
rect 12770 13630 12830 13640
rect 12770 13590 12780 13630
rect 12780 13590 12820 13630
rect 12820 13590 12830 13630
rect 12770 13580 12830 13590
rect 12930 13630 12990 13640
rect 12930 13590 12940 13630
rect 12940 13590 12980 13630
rect 12980 13590 12990 13630
rect 12930 13580 12990 13590
rect 13090 13630 13150 13640
rect 13090 13590 13100 13630
rect 13100 13590 13140 13630
rect 13140 13590 13150 13630
rect 13090 13580 13150 13590
rect 13250 13630 13310 13640
rect 13250 13590 13260 13630
rect 13260 13590 13300 13630
rect 13300 13590 13310 13630
rect 13250 13580 13310 13590
rect 13410 13630 13470 13640
rect 13410 13590 13420 13630
rect 13420 13590 13460 13630
rect 13460 13590 13470 13630
rect 13410 13580 13470 13590
rect 13570 13630 13630 13640
rect 13570 13590 13580 13630
rect 13580 13590 13620 13630
rect 13620 13590 13630 13630
rect 13570 13580 13630 13590
rect 13730 13630 13790 13640
rect 13730 13590 13740 13630
rect 13740 13590 13780 13630
rect 13780 13590 13790 13630
rect 13730 13580 13790 13590
rect 13890 13630 13950 13640
rect 13890 13590 13900 13630
rect 13900 13590 13940 13630
rect 13940 13590 13950 13630
rect 13890 13580 13950 13590
rect 14050 13630 14110 13640
rect 14050 13590 14060 13630
rect 14060 13590 14100 13630
rect 14100 13590 14110 13630
rect 14050 13580 14110 13590
rect 14210 13630 14270 13640
rect 14210 13590 14220 13630
rect 14220 13590 14260 13630
rect 14260 13590 14270 13630
rect 14210 13580 14270 13590
rect 14370 13630 14430 13640
rect 14370 13590 14380 13630
rect 14380 13590 14420 13630
rect 14420 13590 14430 13630
rect 14370 13580 14430 13590
rect 14530 13630 14590 13640
rect 14530 13590 14540 13630
rect 14540 13590 14580 13630
rect 14580 13590 14590 13630
rect 14530 13580 14590 13590
rect 14690 13630 14750 13640
rect 14690 13590 14700 13630
rect 14700 13590 14740 13630
rect 14740 13590 14750 13630
rect 14690 13580 14750 13590
rect 14850 13630 14910 13640
rect 14850 13590 14860 13630
rect 14860 13590 14900 13630
rect 14900 13590 14910 13630
rect 14850 13580 14910 13590
rect 15010 13630 15070 13640
rect 15010 13590 15020 13630
rect 15020 13590 15060 13630
rect 15060 13590 15070 13630
rect 15010 13580 15070 13590
rect 15170 13630 15230 13640
rect 15170 13590 15180 13630
rect 15180 13590 15220 13630
rect 15220 13590 15230 13630
rect 15170 13580 15230 13590
rect 11910 13470 11970 13530
rect 11910 13390 11970 13450
rect 11910 13360 11970 13370
rect 11910 13320 11920 13360
rect 11920 13320 11960 13360
rect 11960 13320 11970 13360
rect 11910 13310 11970 13320
rect 13170 13470 13230 13530
rect 13250 13470 13310 13530
rect 13330 13470 13390 13530
rect 13170 13390 13230 13450
rect 13250 13390 13310 13450
rect 13330 13390 13390 13450
rect 13170 13310 13230 13370
rect 13250 13310 13310 13370
rect 13330 13310 13390 13370
rect 10930 12720 10990 12730
rect 10930 12680 10940 12720
rect 10940 12680 10980 12720
rect 10980 12680 10990 12720
rect 10930 12670 10990 12680
rect 10930 12590 10990 12650
rect 10930 12510 10990 12570
rect 11170 12720 11230 12730
rect 11170 12680 11180 12720
rect 11180 12680 11220 12720
rect 11220 12680 11230 12720
rect 11170 12670 11230 12680
rect 11170 12590 11230 12650
rect 11170 12510 11230 12570
rect 11410 12720 11470 12730
rect 11410 12680 11420 12720
rect 11420 12680 11460 12720
rect 11460 12680 11470 12720
rect 11410 12670 11470 12680
rect 11410 12590 11470 12650
rect 11410 12510 11470 12570
rect 11650 12720 11710 12730
rect 11650 12680 11660 12720
rect 11660 12680 11700 12720
rect 11700 12680 11710 12720
rect 11650 12670 11710 12680
rect 11650 12590 11710 12650
rect 11650 12510 11710 12570
rect 12290 12720 12350 12730
rect 12290 12680 12300 12720
rect 12300 12680 12340 12720
rect 12340 12680 12350 12720
rect 12290 12670 12350 12680
rect 12290 12590 12350 12650
rect 12290 12510 12350 12570
rect 12530 12720 12590 12730
rect 12530 12680 12540 12720
rect 12540 12680 12580 12720
rect 12580 12680 12590 12720
rect 12530 12670 12590 12680
rect 12530 12590 12590 12650
rect 12530 12510 12590 12570
rect 12770 12720 12830 12730
rect 12770 12680 12780 12720
rect 12780 12680 12820 12720
rect 12820 12680 12830 12720
rect 12770 12670 12830 12680
rect 12770 12590 12830 12650
rect 12770 12510 12830 12570
rect 10750 12400 10810 12460
rect 11500 12400 11560 12460
rect 11720 12400 11780 12460
rect 11980 12400 12040 12460
rect 12200 12400 12260 12460
rect 12460 12400 12520 12460
rect 11433 12342 11485 12350
rect 11433 12308 11443 12342
rect 11443 12308 11477 12342
rect 11477 12308 11485 12342
rect 11433 12298 11485 12308
rect 11793 12342 11845 12350
rect 11793 12308 11803 12342
rect 11803 12308 11837 12342
rect 11837 12308 11845 12342
rect 11793 12298 11845 12308
rect 11913 12342 11965 12350
rect 11913 12308 11923 12342
rect 11923 12308 11957 12342
rect 11957 12308 11965 12342
rect 11913 12298 11965 12308
rect 12273 12342 12325 12350
rect 12273 12308 12283 12342
rect 12283 12308 12317 12342
rect 12317 12308 12325 12342
rect 12273 12298 12325 12308
rect 12393 12342 12445 12350
rect 12393 12308 12403 12342
rect 12403 12308 12437 12342
rect 12437 12308 12445 12342
rect 12393 12298 12445 12308
rect 12810 12320 12870 12330
rect 12810 12280 12820 12320
rect 12820 12280 12860 12320
rect 12860 12280 12870 12320
rect 12810 12270 12870 12280
rect 12810 12240 12870 12250
rect 12810 12200 12820 12240
rect 12820 12200 12860 12240
rect 12860 12200 12870 12240
rect 12810 12190 12870 12200
rect 11536 12112 11588 12122
rect 11536 12078 11544 12112
rect 11544 12078 11578 12112
rect 11578 12078 11588 12112
rect 11536 12070 11588 12078
rect 11694 12112 11746 12122
rect 11694 12078 11702 12112
rect 11702 12078 11736 12112
rect 11736 12078 11746 12112
rect 11694 12070 11746 12078
rect 11610 11960 11670 12020
rect 11370 11850 11430 11910
rect 10630 11580 10690 11640
rect 10710 11580 10770 11640
rect 11130 11580 11190 11640
rect 11370 11580 11430 11640
rect 10890 11510 10950 11520
rect 10890 11470 10900 11510
rect 10900 11470 10940 11510
rect 10940 11470 10950 11510
rect 10890 11460 10950 11470
rect 10650 11120 10710 11180
rect 12018 12112 12070 12122
rect 12018 12078 12026 12112
rect 12026 12078 12060 12112
rect 12060 12078 12070 12112
rect 12018 12070 12070 12078
rect 12172 12112 12224 12122
rect 12172 12078 12180 12112
rect 12180 12078 12214 12112
rect 12214 12078 12224 12112
rect 12172 12070 12224 12078
rect 12090 11960 12150 12020
rect 12496 12112 12548 12122
rect 12496 12078 12504 12112
rect 12504 12078 12538 12112
rect 12538 12078 12548 12112
rect 12496 12070 12548 12078
rect 12810 12160 12870 12170
rect 12810 12120 12820 12160
rect 12820 12120 12860 12160
rect 12860 12120 12870 12160
rect 12810 12110 12870 12120
rect 12570 11960 12630 12020
rect 11850 11850 11910 11910
rect 12330 11850 12390 11910
rect 11850 11580 11910 11640
rect 12090 11580 12150 11640
rect 12570 11580 12630 11640
rect 12750 11580 12810 11640
rect 11610 11510 11670 11520
rect 11610 11470 11620 11510
rect 11620 11470 11660 11510
rect 11660 11470 11670 11510
rect 11610 11460 11670 11470
rect 11370 11120 11430 11180
rect 12330 11510 12390 11520
rect 12330 11470 12340 11510
rect 12340 11470 12380 11510
rect 12380 11470 12390 11510
rect 12330 11460 12390 11470
rect 12090 11120 12150 11180
rect 12810 11120 12870 11180
rect 14590 13470 14650 13530
rect 14590 13390 14650 13450
rect 14590 13360 14650 13370
rect 14590 13320 14600 13360
rect 14600 13320 14640 13360
rect 14640 13320 14650 13360
rect 14590 13310 14650 13320
rect 13170 12270 13230 12330
rect 13250 12270 13310 12330
rect 13330 12270 13390 12330
rect 13170 12190 13230 12250
rect 13250 12190 13310 12250
rect 13330 12190 13390 12250
rect 13170 12110 13230 12170
rect 13250 12110 13310 12170
rect 13330 12110 13390 12170
rect 13730 12720 13790 12730
rect 13730 12680 13740 12720
rect 13740 12680 13780 12720
rect 13780 12680 13790 12720
rect 13730 12670 13790 12680
rect 13730 12590 13790 12650
rect 13730 12510 13790 12570
rect 13970 12720 14030 12730
rect 13970 12680 13980 12720
rect 13980 12680 14020 12720
rect 14020 12680 14030 12720
rect 13970 12670 14030 12680
rect 13970 12590 14030 12650
rect 13970 12510 14030 12570
rect 14210 12720 14270 12730
rect 14210 12680 14220 12720
rect 14220 12680 14260 12720
rect 14260 12680 14270 12720
rect 14210 12670 14270 12680
rect 14210 12590 14270 12650
rect 14210 12510 14270 12570
rect 14850 12720 14910 12730
rect 14850 12680 14860 12720
rect 14860 12680 14900 12720
rect 14900 12680 14910 12720
rect 14850 12670 14910 12680
rect 14850 12590 14910 12650
rect 14850 12510 14910 12570
rect 15090 12720 15150 12730
rect 15090 12680 15100 12720
rect 15100 12680 15140 12720
rect 15140 12680 15150 12720
rect 15090 12670 15150 12680
rect 15090 12590 15150 12650
rect 15090 12510 15150 12570
rect 15330 12720 15390 12730
rect 15330 12680 15340 12720
rect 15340 12680 15380 12720
rect 15380 12680 15390 12720
rect 15330 12670 15390 12680
rect 15330 12590 15390 12650
rect 15330 12510 15390 12570
rect 15570 12720 15630 12730
rect 15570 12680 15580 12720
rect 15580 12680 15620 12720
rect 15620 12680 15630 12720
rect 15570 12670 15630 12680
rect 15570 12590 15630 12650
rect 15570 12510 15630 12570
rect 14040 12400 14100 12460
rect 14300 12400 14360 12460
rect 14520 12400 14580 12460
rect 14780 12400 14840 12460
rect 15000 12400 15060 12460
rect 15750 12400 15810 12460
rect 13690 12320 13750 12330
rect 13690 12280 13700 12320
rect 13700 12280 13740 12320
rect 13740 12280 13750 12320
rect 13690 12270 13750 12280
rect 14115 12342 14167 12350
rect 14115 12308 14123 12342
rect 14123 12308 14157 12342
rect 14157 12308 14167 12342
rect 14115 12298 14167 12308
rect 14235 12342 14287 12350
rect 14235 12308 14243 12342
rect 14243 12308 14277 12342
rect 14277 12308 14287 12342
rect 14235 12298 14287 12308
rect 14595 12342 14647 12350
rect 14595 12308 14603 12342
rect 14603 12308 14637 12342
rect 14637 12308 14647 12342
rect 14595 12298 14647 12308
rect 14715 12342 14767 12350
rect 14715 12308 14723 12342
rect 14723 12308 14757 12342
rect 14757 12308 14767 12342
rect 14715 12298 14767 12308
rect 15075 12342 15127 12350
rect 15075 12308 15083 12342
rect 15083 12308 15117 12342
rect 15117 12308 15127 12342
rect 15075 12298 15127 12308
rect 16160 12290 16220 12350
rect 13690 12240 13750 12250
rect 13690 12200 13700 12240
rect 13700 12200 13740 12240
rect 13740 12200 13750 12240
rect 13690 12190 13750 12200
rect 13690 12160 13750 12170
rect 13690 12120 13700 12160
rect 13700 12120 13740 12160
rect 13740 12120 13750 12160
rect 13690 12110 13750 12120
rect 14012 12112 14064 12122
rect 14012 12078 14022 12112
rect 14022 12078 14056 12112
rect 14056 12078 14064 12112
rect 14012 12070 14064 12078
rect 13930 11960 13990 12020
rect 14336 12112 14388 12122
rect 14336 12078 14346 12112
rect 14346 12078 14380 12112
rect 14380 12078 14388 12112
rect 14336 12070 14388 12078
rect 14490 12112 14542 12122
rect 14490 12078 14500 12112
rect 14500 12078 14534 12112
rect 14534 12078 14542 12112
rect 14490 12070 14542 12078
rect 14410 11960 14470 12020
rect 14814 12112 14866 12122
rect 14814 12078 14824 12112
rect 14824 12078 14858 12112
rect 14858 12078 14866 12112
rect 14814 12070 14866 12078
rect 14972 12112 15024 12122
rect 14972 12078 14982 12112
rect 14982 12078 15016 12112
rect 15016 12078 15024 12112
rect 14972 12070 15024 12078
rect 14890 11960 14950 12020
rect 14170 11850 14230 11910
rect 14650 11850 14710 11910
rect 13750 11740 13810 11800
rect 13750 11660 13810 11720
rect 13750 11580 13810 11640
rect 13930 11740 13990 11800
rect 13930 11660 13990 11720
rect 13930 11580 13990 11640
rect 14170 11740 14230 11800
rect 14170 11660 14230 11720
rect 14170 11580 14230 11640
rect 14410 11740 14470 11800
rect 14410 11660 14470 11720
rect 14410 11580 14470 11640
rect 14650 11740 14710 11800
rect 14650 11660 14710 11720
rect 14650 11580 14710 11640
rect 13070 11120 13130 11180
rect 13430 11120 13490 11180
rect 10530 11010 10590 11070
rect 10530 10930 10590 10990
rect 10530 10850 10590 10910
rect 10770 11010 10830 11070
rect 10770 10930 10830 10990
rect 10770 10850 10830 10910
rect 11010 11010 11070 11070
rect 11010 10930 11070 10990
rect 11010 10850 11070 10910
rect 11250 11010 11310 11070
rect 11250 10930 11310 10990
rect 11250 10850 11310 10910
rect 11490 11010 11550 11070
rect 11490 10930 11550 10990
rect 11490 10850 11550 10910
rect 11730 11010 11790 11070
rect 11730 10930 11790 10990
rect 11730 10850 11790 10910
rect 11970 11010 12030 11070
rect 11970 10930 12030 10990
rect 11970 10850 12030 10910
rect 12210 11010 12270 11070
rect 12210 10930 12270 10990
rect 12210 10850 12270 10910
rect 12450 11010 12510 11070
rect 12450 10930 12510 10990
rect 12450 10850 12510 10910
rect 12690 11010 12750 11070
rect 12690 10930 12750 10990
rect 12690 10850 12750 10910
rect 12930 11010 12990 11070
rect 12930 10930 12990 10990
rect 12930 10850 12990 10910
rect 11810 10740 11870 10800
rect 13250 10740 13310 10800
rect 12170 10630 12230 10690
rect 11900 10350 11960 10360
rect 11900 10310 11910 10350
rect 11910 10310 11950 10350
rect 11950 10310 11960 10350
rect 11900 10300 11960 10310
rect 12080 10350 12140 10360
rect 12080 10310 12090 10350
rect 12090 10310 12130 10350
rect 12130 10310 12140 10350
rect 12080 10300 12140 10310
rect 12530 10520 12590 10580
rect 12260 10350 12320 10360
rect 12260 10310 12270 10350
rect 12270 10310 12310 10350
rect 12310 10310 12320 10350
rect 12260 10300 12320 10310
rect 12440 10350 12500 10360
rect 12440 10310 12450 10350
rect 12450 10310 12490 10350
rect 12490 10310 12500 10350
rect 12440 10300 12500 10310
rect 12890 10410 12950 10470
rect 12620 10350 12680 10360
rect 12620 10310 12630 10350
rect 12630 10310 12670 10350
rect 12670 10310 12680 10350
rect 12620 10300 12680 10310
rect 12800 10350 12860 10360
rect 12800 10310 12810 10350
rect 12810 10310 12850 10350
rect 12850 10310 12860 10350
rect 12800 10300 12860 10310
rect 12980 10350 13040 10360
rect 12980 10310 12990 10350
rect 12990 10310 13030 10350
rect 13030 10310 13040 10350
rect 12980 10300 13040 10310
rect 13160 10350 13220 10360
rect 13160 10310 13170 10350
rect 13170 10310 13210 10350
rect 13210 10310 13220 10350
rect 13160 10300 13220 10310
rect 13690 11120 13750 11180
rect 14170 11510 14230 11520
rect 14170 11470 14180 11510
rect 14180 11470 14220 11510
rect 14220 11470 14230 11510
rect 14170 11460 14230 11470
rect 14410 11120 14470 11180
rect 15130 11850 15190 11910
rect 15130 11740 15190 11800
rect 15130 11660 15190 11720
rect 15130 11580 15190 11640
rect 15370 11740 15430 11800
rect 15370 11660 15430 11720
rect 15370 11580 15430 11640
rect 15790 11740 15850 11800
rect 15790 11660 15850 11720
rect 15790 11580 15850 11640
rect 14890 11510 14950 11520
rect 14890 11470 14900 11510
rect 14900 11470 14940 11510
rect 14940 11470 14950 11510
rect 14890 11460 14950 11470
rect 15130 11120 15190 11180
rect 15610 11510 15670 11520
rect 15610 11470 15620 11510
rect 15620 11470 15660 11510
rect 15660 11470 15670 11510
rect 15610 11460 15670 11470
rect 15850 11120 15910 11180
rect 13570 11010 13630 11070
rect 13570 10930 13630 10990
rect 13570 10850 13630 10910
rect 13810 11010 13870 11070
rect 13810 10930 13870 10990
rect 13810 10850 13870 10910
rect 14050 11010 14110 11070
rect 14050 10930 14110 10990
rect 14050 10850 14110 10910
rect 14290 11010 14350 11070
rect 14290 10930 14350 10990
rect 14290 10850 14350 10910
rect 14530 11010 14590 11070
rect 14530 10930 14590 10990
rect 14530 10850 14590 10910
rect 14770 11010 14830 11070
rect 14770 10930 14830 10990
rect 14770 10850 14830 10910
rect 15010 11010 15070 11070
rect 15010 10930 15070 10990
rect 15010 10850 15070 10910
rect 15250 11010 15310 11070
rect 15250 10930 15310 10990
rect 15250 10850 15310 10910
rect 15490 11010 15550 11070
rect 15490 10930 15550 10990
rect 15490 10850 15550 10910
rect 15730 11010 15790 11070
rect 15730 10930 15790 10990
rect 15730 10850 15790 10910
rect 14690 10740 14750 10800
rect 14330 10630 14390 10690
rect 13970 10520 14030 10580
rect 13610 10410 13670 10470
rect 13340 10350 13400 10360
rect 13340 10310 13350 10350
rect 13350 10310 13390 10350
rect 13390 10310 13400 10350
rect 13340 10300 13400 10310
rect 13430 10300 13490 10360
rect 13520 10350 13580 10360
rect 13520 10310 13530 10350
rect 13530 10310 13570 10350
rect 13570 10310 13580 10350
rect 13520 10300 13580 10310
rect 13700 10350 13760 10360
rect 13700 10310 13710 10350
rect 13710 10310 13750 10350
rect 13750 10310 13760 10350
rect 13700 10300 13760 10310
rect 13880 10350 13940 10360
rect 13880 10310 13890 10350
rect 13890 10310 13930 10350
rect 13930 10310 13940 10350
rect 13880 10300 13940 10310
rect 14060 10350 14120 10360
rect 14060 10310 14070 10350
rect 14070 10310 14110 10350
rect 14110 10310 14120 10350
rect 14060 10300 14120 10310
rect 14240 10350 14300 10360
rect 14240 10310 14250 10350
rect 14250 10310 14290 10350
rect 14290 10310 14300 10350
rect 14240 10300 14300 10310
rect 14420 10350 14480 10360
rect 14420 10310 14430 10350
rect 14430 10310 14470 10350
rect 14470 10310 14480 10350
rect 14420 10300 14480 10310
rect 14600 10350 14660 10360
rect 14600 10310 14610 10350
rect 14610 10310 14650 10350
rect 14650 10310 14660 10350
rect 14600 10300 14660 10310
rect 15720 10630 15780 10690
rect 15250 10520 15310 10580
rect 15600 10150 15660 10160
rect 15600 10110 15610 10150
rect 15610 10110 15650 10150
rect 15650 10110 15660 10150
rect 15600 10100 15660 10110
rect 15970 11010 16030 11070
rect 15970 10930 16030 10990
rect 15970 10850 16030 10910
rect 16250 12060 16310 12120
rect 16790 14030 16850 14090
rect 16360 11740 16420 11800
rect 16440 11740 16500 11800
rect 16520 11740 16580 11800
rect 16360 11660 16420 11720
rect 16440 11660 16500 11720
rect 16520 11660 16580 11720
rect 16360 11580 16420 11640
rect 16440 11580 16500 11640
rect 16520 11580 16580 11640
rect 17960 15990 18020 16050
rect 18130 17390 18190 17450
rect 18800 16690 18860 16750
rect 18800 15290 18860 15350
rect 18660 13920 18720 13980
rect 17580 11120 17640 11180
rect 16250 10520 16310 10580
rect 16160 10410 16220 10470
rect 15840 10150 15900 10160
rect 15840 10110 15850 10150
rect 15850 10110 15890 10150
rect 15890 10110 15900 10150
rect 15840 10100 15900 10110
rect 15250 9760 15310 9820
rect 15720 9810 15780 9820
rect 15720 9770 15730 9810
rect 15730 9770 15770 9810
rect 15770 9770 15780 9810
rect 15720 9760 15780 9770
rect 11630 9610 11690 9620
rect 11630 9570 11640 9610
rect 11640 9570 11680 9610
rect 11680 9570 11690 9610
rect 11630 9560 11690 9570
rect 11630 9480 11690 9540
rect 11630 9400 11690 9460
rect 11990 9610 12050 9620
rect 11990 9570 12000 9610
rect 12000 9570 12040 9610
rect 12040 9570 12050 9610
rect 11990 9560 12050 9570
rect 11990 9480 12050 9540
rect 11990 9400 12050 9460
rect 12350 9610 12410 9620
rect 12350 9570 12360 9610
rect 12360 9570 12400 9610
rect 12400 9570 12410 9610
rect 12350 9560 12410 9570
rect 12350 9480 12410 9540
rect 12350 9400 12410 9460
rect 12710 9610 12770 9620
rect 12710 9570 12720 9610
rect 12720 9570 12760 9610
rect 12760 9570 12770 9610
rect 12710 9560 12770 9570
rect 12710 9480 12770 9540
rect 12710 9400 12770 9460
rect 13070 9610 13130 9620
rect 13070 9570 13080 9610
rect 13080 9570 13120 9610
rect 13120 9570 13130 9610
rect 13070 9560 13130 9570
rect 13070 9480 13130 9540
rect 13070 9400 13130 9460
rect 13430 9610 13490 9620
rect 13430 9570 13440 9610
rect 13440 9570 13480 9610
rect 13480 9570 13490 9610
rect 13430 9560 13490 9570
rect 13430 9480 13490 9540
rect 13430 9400 13490 9460
rect 13790 9610 13850 9620
rect 13790 9570 13800 9610
rect 13800 9570 13840 9610
rect 13840 9570 13850 9610
rect 13790 9560 13850 9570
rect 13790 9480 13850 9540
rect 13790 9400 13850 9460
rect 14150 9610 14210 9620
rect 14150 9570 14160 9610
rect 14160 9570 14200 9610
rect 14200 9570 14210 9610
rect 14150 9560 14210 9570
rect 14150 9480 14210 9540
rect 14150 9400 14210 9460
rect 14510 9610 14570 9620
rect 14510 9570 14520 9610
rect 14520 9570 14560 9610
rect 14560 9570 14570 9610
rect 14510 9560 14570 9570
rect 14510 9480 14570 9540
rect 14510 9400 14570 9460
rect 14870 9610 14930 9620
rect 14870 9570 14880 9610
rect 14880 9570 14920 9610
rect 14920 9570 14930 9610
rect 14870 9560 14930 9570
rect 14870 9480 14930 9540
rect 14870 9400 14930 9460
rect 15500 9560 15560 9620
rect 15500 9480 15560 9540
rect 15500 9400 15560 9460
rect 15940 9560 16000 9620
rect 15940 9480 16000 9540
rect 15940 9400 16000 9460
rect 11808 9342 11860 9350
rect 11808 9308 11818 9342
rect 11818 9308 11852 9342
rect 11852 9308 11860 9342
rect 11808 9298 11860 9308
rect 11918 9342 11970 9350
rect 11918 9308 11928 9342
rect 11928 9308 11962 9342
rect 11962 9308 11970 9342
rect 11918 9298 11970 9308
rect 12028 9342 12080 9350
rect 12028 9308 12038 9342
rect 12038 9308 12072 9342
rect 12072 9308 12080 9342
rect 12028 9298 12080 9308
rect 12138 9342 12190 9350
rect 12138 9308 12148 9342
rect 12148 9308 12182 9342
rect 12182 9308 12190 9342
rect 12138 9298 12190 9308
rect 12248 9342 12300 9350
rect 12248 9308 12258 9342
rect 12258 9308 12292 9342
rect 12292 9308 12300 9342
rect 12248 9298 12300 9308
rect 12358 9342 12410 9350
rect 12358 9308 12368 9342
rect 12368 9308 12402 9342
rect 12402 9308 12410 9342
rect 12358 9298 12410 9308
rect 12468 9342 12520 9350
rect 12468 9308 12478 9342
rect 12478 9308 12512 9342
rect 12512 9308 12520 9342
rect 12468 9298 12520 9308
rect 12578 9342 12630 9350
rect 12578 9308 12588 9342
rect 12588 9308 12622 9342
rect 12622 9308 12630 9342
rect 12578 9298 12630 9308
rect 12688 9342 12740 9350
rect 12688 9308 12698 9342
rect 12698 9308 12732 9342
rect 12732 9308 12740 9342
rect 12688 9298 12740 9308
rect 12798 9342 12850 9350
rect 12798 9308 12808 9342
rect 12808 9308 12842 9342
rect 12842 9308 12850 9342
rect 12798 9298 12850 9308
rect 13708 9342 13760 9350
rect 13708 9308 13718 9342
rect 13718 9308 13752 9342
rect 13752 9308 13760 9342
rect 13708 9298 13760 9308
rect 13818 9342 13870 9350
rect 13818 9308 13828 9342
rect 13828 9308 13862 9342
rect 13862 9308 13870 9342
rect 13818 9298 13870 9308
rect 13928 9342 13980 9350
rect 13928 9308 13938 9342
rect 13938 9308 13972 9342
rect 13972 9308 13980 9342
rect 13928 9298 13980 9308
rect 14038 9342 14090 9350
rect 14038 9308 14048 9342
rect 14048 9308 14082 9342
rect 14082 9308 14090 9342
rect 14038 9298 14090 9308
rect 14148 9342 14200 9350
rect 14148 9308 14158 9342
rect 14158 9308 14192 9342
rect 14192 9308 14200 9342
rect 14148 9298 14200 9308
rect 14258 9342 14310 9350
rect 14258 9308 14268 9342
rect 14268 9308 14302 9342
rect 14302 9308 14310 9342
rect 14258 9298 14310 9308
rect 14368 9342 14420 9350
rect 14368 9308 14378 9342
rect 14378 9308 14412 9342
rect 14412 9308 14420 9342
rect 14368 9298 14420 9308
rect 14478 9342 14530 9350
rect 14478 9308 14488 9342
rect 14488 9308 14522 9342
rect 14522 9308 14530 9342
rect 14478 9298 14530 9308
rect 14588 9342 14640 9350
rect 14588 9308 14598 9342
rect 14598 9308 14632 9342
rect 14632 9308 14640 9342
rect 14588 9298 14640 9308
rect 14698 9342 14750 9350
rect 14698 9308 14708 9342
rect 14708 9308 14742 9342
rect 14742 9308 14750 9342
rect 14698 9298 14750 9308
rect 11640 9010 11700 9020
rect 11640 8970 11650 9010
rect 11650 8970 11690 9010
rect 11690 8970 11700 9010
rect 11640 8960 11700 8970
rect 11860 8960 11920 9020
rect 12080 8960 12140 9020
rect 12300 8960 12360 9020
rect 12520 8960 12580 9020
rect 12740 8960 12800 9020
rect 12960 9010 13020 9020
rect 12960 8970 12970 9010
rect 12970 8970 13010 9010
rect 13010 8970 13020 9010
rect 12960 8960 13020 8970
rect 13540 9010 13600 9020
rect 13540 8970 13550 9010
rect 13550 8970 13590 9010
rect 13590 8970 13600 9010
rect 13540 8960 13600 8970
rect 9690 8850 9750 8910
rect 11750 8850 11810 8910
rect 11970 8850 12030 8910
rect 12190 8850 12250 8910
rect 12410 8850 12470 8910
rect 12630 8850 12690 8910
rect 13760 8960 13820 9020
rect 13980 8960 14040 9020
rect 14200 8960 14260 9020
rect 14420 8960 14480 9020
rect 14640 8960 14700 9020
rect 14860 9010 14920 9020
rect 14860 8970 14870 9010
rect 14870 8970 14910 9010
rect 14910 8970 14920 9010
rect 14860 8960 14920 8970
rect 12850 8850 12910 8910
rect 13650 8840 13710 8900
rect 13650 8760 13710 8820
rect 13650 8680 13710 8740
rect 13870 8840 13930 8900
rect 13870 8760 13930 8820
rect 13870 8680 13930 8740
rect 14090 8840 14150 8900
rect 14090 8760 14150 8820
rect 14090 8680 14150 8740
rect 14310 8840 14370 8900
rect 14310 8760 14370 8820
rect 14310 8680 14370 8740
rect 14530 8840 14590 8900
rect 14530 8760 14590 8820
rect 14530 8680 14590 8740
rect 14750 8840 14810 8900
rect 14750 8760 14810 8820
rect 14750 8680 14810 8740
<< metal2 >>
rect 9170 19190 18270 19200
rect 9170 19130 9180 19190
rect 9240 19130 18200 19190
rect 18260 19130 18270 19190
rect 9170 19120 18270 19130
rect 8790 19080 17650 19090
rect 8790 19020 8800 19080
rect 8860 19020 9580 19080
rect 9640 19020 10690 19080
rect 10750 19020 13250 19080
rect 13310 19020 15680 19080
rect 15740 19020 16790 19080
rect 16850 19020 17580 19080
rect 17640 19020 17650 19080
rect 8790 19000 17650 19020
rect 8790 18940 8800 19000
rect 8860 18940 9580 19000
rect 9640 18940 10690 19000
rect 10750 18940 13250 19000
rect 13310 18940 15680 19000
rect 15740 18940 16790 19000
rect 16850 18940 17580 19000
rect 17640 18940 17650 19000
rect 8790 18920 17650 18940
rect 8790 18860 8800 18920
rect 8860 18860 9580 18920
rect 9640 18860 10690 18920
rect 10750 18860 13250 18920
rect 13310 18860 15680 18920
rect 15740 18860 16790 18920
rect 16850 18860 17580 18920
rect 17640 18860 17650 18920
rect 8790 18850 17650 18860
rect 18190 18850 18270 18860
rect 18190 18790 18200 18850
rect 18260 18790 18270 18850
rect 18190 18780 18270 18790
rect 8770 18450 9250 18460
rect 8770 18420 9180 18450
rect 8770 18050 8790 18420
rect 8870 18390 9180 18420
rect 9240 18390 9250 18450
rect 8870 18370 9250 18390
rect 8870 18310 9180 18370
rect 9240 18310 9250 18370
rect 8870 18280 9250 18310
rect 8870 18220 9180 18280
rect 9240 18220 9250 18280
rect 8870 18190 9250 18220
rect 8870 18130 9180 18190
rect 9240 18130 9250 18190
rect 8870 18110 9250 18130
rect 8870 18050 9180 18110
rect 9240 18050 9250 18110
rect 8770 18030 9250 18050
rect 17550 18450 18030 18460
rect 17550 18420 17960 18450
rect 17550 18050 17570 18420
rect 17650 18390 17960 18420
rect 18020 18390 18030 18450
rect 17650 18370 18030 18390
rect 17650 18310 17960 18370
rect 18020 18310 18030 18370
rect 17650 18280 18030 18310
rect 17650 18220 17960 18280
rect 18020 18220 18030 18280
rect 17650 18190 18030 18220
rect 17650 18130 17960 18190
rect 18020 18130 18030 18190
rect 17650 18110 18030 18130
rect 17650 18050 17960 18110
rect 18020 18050 18030 18110
rect 18640 18150 18740 18170
rect 18640 18090 18660 18150
rect 18720 18090 18740 18150
rect 18640 18070 18740 18090
rect 17550 18030 18030 18050
rect 18120 17450 18200 17460
rect 18120 17390 18130 17450
rect 18190 17390 18200 17450
rect 18120 17380 18200 17390
rect 11140 16810 11650 16820
rect 11140 16750 11150 16810
rect 11210 16750 11580 16810
rect 11640 16750 11650 16810
rect 11140 16740 11650 16750
rect 13240 16810 15420 16820
rect 13240 16750 13250 16810
rect 13310 16750 15350 16810
rect 15410 16750 15420 16810
rect 13240 16740 15420 16750
rect 17560 16760 18880 16770
rect 17560 16680 17570 16760
rect 17650 16750 18880 16760
rect 17650 16690 18800 16750
rect 18860 16690 18880 16750
rect 17650 16680 18880 16690
rect 17560 16670 18880 16680
rect 17950 16050 19070 16060
rect 17950 15990 17960 16050
rect 18020 15990 19000 16050
rect 19060 15990 19070 16050
rect 17950 15980 19070 15990
rect 16350 15350 18880 15370
rect 16350 15290 16360 15350
rect 16420 15290 16440 15350
rect 16500 15290 16520 15350
rect 16580 15290 18800 15350
rect 18860 15290 18880 15350
rect 16350 15270 18880 15290
rect 15340 14800 16320 14810
rect 15340 14740 15350 14800
rect 15410 14740 16010 14800
rect 16070 14740 16250 14800
rect 16310 14740 16320 14800
rect 15340 14730 16320 14740
rect 10350 14720 15020 14730
rect 10350 14660 10360 14720
rect 10420 14660 14590 14720
rect 14650 14660 14680 14720
rect 14740 14660 14770 14720
rect 14830 14660 14860 14720
rect 14920 14660 14950 14720
rect 15010 14660 15020 14720
rect 10350 14650 15020 14660
rect 11140 14410 11980 14420
rect 11140 14350 11150 14410
rect 11210 14402 11980 14410
rect 11210 14350 11560 14402
rect 11960 14350 11980 14402
rect 11140 14340 11980 14350
rect 14580 14410 16230 14420
rect 14580 14402 16160 14410
rect 14580 14350 14600 14402
rect 15000 14350 16160 14402
rect 16220 14350 16230 14410
rect 14580 14340 16230 14350
rect 9680 14090 16860 14100
rect 9680 14030 9690 14090
rect 9750 14030 16790 14090
rect 16850 14030 16860 14090
rect 9680 14020 16860 14030
rect 10620 13980 18730 13990
rect 10620 13920 10630 13980
rect 10690 13920 11040 13980
rect 11100 13920 18660 13980
rect 18720 13920 18730 13980
rect 10620 13910 18730 13920
rect 15470 13850 15550 13860
rect 9460 13810 11160 13820
rect 9460 13750 9470 13810
rect 9530 13750 11090 13810
rect 11150 13750 11160 13810
rect 9460 13740 11160 13750
rect 15470 13790 15480 13850
rect 15540 13790 15550 13850
rect 15470 13770 15550 13790
rect 15470 13710 15480 13770
rect 15540 13710 15550 13770
rect 15470 13700 15550 13710
rect 11160 13640 11240 13650
rect 11160 13580 11170 13640
rect 11230 13630 11240 13640
rect 11320 13640 11400 13650
rect 11320 13630 11330 13640
rect 11230 13590 11330 13630
rect 11230 13580 11240 13590
rect 11160 13570 11240 13580
rect 11320 13580 11330 13590
rect 11390 13630 11400 13640
rect 11480 13640 11560 13650
rect 11480 13630 11490 13640
rect 11390 13590 11490 13630
rect 11390 13580 11400 13590
rect 11320 13570 11400 13580
rect 11480 13580 11490 13590
rect 11550 13630 11560 13640
rect 11640 13640 11720 13650
rect 11640 13630 11650 13640
rect 11550 13590 11650 13630
rect 11550 13580 11560 13590
rect 11480 13570 11560 13580
rect 11640 13580 11650 13590
rect 11710 13630 11720 13640
rect 11800 13640 11880 13650
rect 11800 13630 11810 13640
rect 11710 13590 11810 13630
rect 11710 13580 11720 13590
rect 11640 13570 11720 13580
rect 11800 13580 11810 13590
rect 11870 13630 11880 13640
rect 11960 13640 12040 13650
rect 11960 13630 11970 13640
rect 11870 13590 11970 13630
rect 11870 13580 11880 13590
rect 11800 13570 11880 13580
rect 11960 13580 11970 13590
rect 12030 13630 12040 13640
rect 12120 13640 12200 13650
rect 12120 13630 12130 13640
rect 12030 13590 12130 13630
rect 12030 13580 12040 13590
rect 11960 13570 12040 13580
rect 12120 13580 12130 13590
rect 12190 13630 12200 13640
rect 12280 13640 12360 13650
rect 12280 13630 12290 13640
rect 12190 13590 12290 13630
rect 12190 13580 12200 13590
rect 12120 13570 12200 13580
rect 12280 13580 12290 13590
rect 12350 13630 12360 13640
rect 12440 13640 12520 13650
rect 12440 13630 12450 13640
rect 12350 13590 12450 13630
rect 12350 13580 12360 13590
rect 12280 13570 12360 13580
rect 12440 13580 12450 13590
rect 12510 13630 12520 13640
rect 12600 13640 12680 13650
rect 12600 13630 12610 13640
rect 12510 13590 12610 13630
rect 12510 13580 12520 13590
rect 12440 13570 12520 13580
rect 12600 13580 12610 13590
rect 12670 13630 12680 13640
rect 12760 13640 12840 13650
rect 12760 13630 12770 13640
rect 12670 13590 12770 13630
rect 12670 13580 12680 13590
rect 12600 13570 12680 13580
rect 12760 13580 12770 13590
rect 12830 13630 12840 13640
rect 12920 13640 13000 13650
rect 12920 13630 12930 13640
rect 12830 13590 12930 13630
rect 12830 13580 12840 13590
rect 12760 13570 12840 13580
rect 12920 13580 12930 13590
rect 12990 13630 13000 13640
rect 13080 13640 13160 13650
rect 13080 13630 13090 13640
rect 12990 13590 13090 13630
rect 12990 13580 13000 13590
rect 12920 13570 13000 13580
rect 13080 13580 13090 13590
rect 13150 13580 13160 13640
rect 13080 13570 13160 13580
rect 13240 13640 13320 13650
rect 13240 13580 13250 13640
rect 13310 13630 13320 13640
rect 13400 13640 13480 13650
rect 13400 13630 13410 13640
rect 13310 13590 13410 13630
rect 13310 13580 13320 13590
rect 13240 13570 13320 13580
rect 13400 13580 13410 13590
rect 13470 13630 13480 13640
rect 13560 13640 13640 13650
rect 13560 13630 13570 13640
rect 13470 13590 13570 13630
rect 13470 13580 13480 13590
rect 13400 13570 13480 13580
rect 13560 13580 13570 13590
rect 13630 13630 13640 13640
rect 13720 13640 13800 13650
rect 13720 13630 13730 13640
rect 13630 13590 13730 13630
rect 13630 13580 13640 13590
rect 13560 13570 13640 13580
rect 13720 13580 13730 13590
rect 13790 13630 13800 13640
rect 13880 13640 13960 13650
rect 13880 13630 13890 13640
rect 13790 13590 13890 13630
rect 13790 13580 13800 13590
rect 13720 13570 13800 13580
rect 13880 13580 13890 13590
rect 13950 13630 13960 13640
rect 14040 13640 14120 13650
rect 14040 13630 14050 13640
rect 13950 13590 14050 13630
rect 13950 13580 13960 13590
rect 13880 13570 13960 13580
rect 14040 13580 14050 13590
rect 14110 13630 14120 13640
rect 14200 13640 14280 13650
rect 14200 13630 14210 13640
rect 14110 13590 14210 13630
rect 14110 13580 14120 13590
rect 14040 13570 14120 13580
rect 14200 13580 14210 13590
rect 14270 13630 14280 13640
rect 14360 13640 14440 13650
rect 14360 13630 14370 13640
rect 14270 13590 14370 13630
rect 14270 13580 14280 13590
rect 14200 13570 14280 13580
rect 14360 13580 14370 13590
rect 14430 13630 14440 13640
rect 14520 13640 14600 13650
rect 14520 13630 14530 13640
rect 14430 13590 14530 13630
rect 14430 13580 14440 13590
rect 14360 13570 14440 13580
rect 14520 13580 14530 13590
rect 14590 13630 14600 13640
rect 14680 13640 14760 13650
rect 14680 13630 14690 13640
rect 14590 13590 14690 13630
rect 14590 13580 14600 13590
rect 14520 13570 14600 13580
rect 14680 13580 14690 13590
rect 14750 13630 14760 13640
rect 14840 13640 14920 13650
rect 14840 13630 14850 13640
rect 14750 13590 14850 13630
rect 14750 13580 14760 13590
rect 14680 13570 14760 13580
rect 14840 13580 14850 13590
rect 14910 13630 14920 13640
rect 15000 13640 15080 13650
rect 15000 13630 15010 13640
rect 14910 13590 15010 13630
rect 14910 13580 14920 13590
rect 14840 13570 14920 13580
rect 15000 13580 15010 13590
rect 15070 13630 15080 13640
rect 15160 13640 15240 13650
rect 15160 13630 15170 13640
rect 15070 13590 15170 13630
rect 15070 13580 15080 13590
rect 15000 13570 15080 13580
rect 15160 13580 15170 13590
rect 15230 13580 15240 13640
rect 15160 13570 15240 13580
rect 11900 13530 14660 13540
rect 11900 13470 11910 13530
rect 11970 13470 13170 13530
rect 13230 13470 13250 13530
rect 13310 13470 13330 13530
rect 13390 13470 14590 13530
rect 14650 13470 14660 13530
rect 11900 13450 14660 13470
rect 11900 13390 11910 13450
rect 11970 13390 13170 13450
rect 13230 13390 13250 13450
rect 13310 13390 13330 13450
rect 13390 13390 14590 13450
rect 14650 13390 14660 13450
rect 11900 13370 14660 13390
rect 11900 13310 11910 13370
rect 11970 13310 13170 13370
rect 13230 13310 13250 13370
rect 13310 13310 13330 13370
rect 13390 13310 14590 13370
rect 14650 13310 14660 13370
rect 11900 13300 14660 13310
rect 10920 12730 15640 12740
rect 10920 12670 10930 12730
rect 10990 12670 11170 12730
rect 11230 12670 11410 12730
rect 11470 12670 11650 12730
rect 11710 12670 12290 12730
rect 12350 12670 12530 12730
rect 12590 12670 12770 12730
rect 12830 12670 13730 12730
rect 13790 12670 13970 12730
rect 14030 12670 14210 12730
rect 14270 12670 14850 12730
rect 14910 12670 15090 12730
rect 15150 12670 15330 12730
rect 15390 12670 15570 12730
rect 15630 12670 15640 12730
rect 10920 12650 15640 12670
rect 10920 12590 10930 12650
rect 10990 12590 11170 12650
rect 11230 12590 11410 12650
rect 11470 12590 11650 12650
rect 11710 12590 12290 12650
rect 12350 12590 12530 12650
rect 12590 12590 12770 12650
rect 12830 12590 13730 12650
rect 13790 12590 13970 12650
rect 14030 12590 14210 12650
rect 14270 12590 14850 12650
rect 14910 12590 15090 12650
rect 15150 12590 15330 12650
rect 15390 12590 15570 12650
rect 15630 12590 15640 12650
rect 10920 12570 15640 12590
rect 10920 12510 10930 12570
rect 10990 12510 11170 12570
rect 11230 12510 11410 12570
rect 11470 12510 11650 12570
rect 11710 12510 12290 12570
rect 12350 12510 12530 12570
rect 12590 12510 12770 12570
rect 12830 12510 13730 12570
rect 13790 12510 13970 12570
rect 14030 12510 14210 12570
rect 14270 12510 14850 12570
rect 14910 12510 15090 12570
rect 15150 12510 15330 12570
rect 15390 12510 15570 12570
rect 15630 12510 15640 12570
rect 10920 12500 15640 12510
rect 10740 12460 12530 12470
rect 10740 12400 10750 12460
rect 10810 12400 11500 12460
rect 11560 12400 11720 12460
rect 11780 12400 11980 12460
rect 12040 12400 12200 12460
rect 12260 12400 12460 12460
rect 12520 12400 12530 12460
rect 10740 12390 12530 12400
rect 14030 12460 15820 12470
rect 14030 12400 14040 12460
rect 14100 12400 14300 12460
rect 14360 12400 14520 12460
rect 14580 12400 14780 12460
rect 14840 12400 15000 12460
rect 15060 12400 15750 12460
rect 15810 12400 15820 12460
rect 14030 12390 15820 12400
rect 9680 12350 12449 12360
rect 9680 12290 9690 12350
rect 9750 12298 11433 12350
rect 11485 12298 11793 12350
rect 11845 12298 11913 12350
rect 11965 12298 12273 12350
rect 12325 12298 12393 12350
rect 12445 12298 12449 12350
rect 14111 12350 16230 12360
rect 9750 12290 12449 12298
rect 12800 12330 13760 12340
rect 9680 12280 9760 12290
rect 12800 12270 12810 12330
rect 12870 12270 13170 12330
rect 13230 12270 13250 12330
rect 13310 12270 13330 12330
rect 13390 12270 13690 12330
rect 13750 12270 13760 12330
rect 14111 12298 14115 12350
rect 14167 12298 14235 12350
rect 14287 12298 14595 12350
rect 14647 12298 14715 12350
rect 14767 12298 15075 12350
rect 15127 12298 16160 12350
rect 14111 12290 16160 12298
rect 16220 12290 16230 12350
rect 16150 12280 16230 12290
rect 12800 12250 13760 12270
rect 12800 12190 12810 12250
rect 12870 12190 13170 12250
rect 13230 12190 13250 12250
rect 13310 12190 13330 12250
rect 13390 12190 13690 12250
rect 13750 12190 13760 12250
rect 12800 12170 13760 12190
rect 9570 12122 12550 12130
rect 9570 12120 11536 12122
rect 9570 12060 9580 12120
rect 9640 12070 11536 12120
rect 11588 12070 11694 12122
rect 11746 12070 12018 12122
rect 12070 12070 12172 12122
rect 12224 12070 12496 12122
rect 12548 12070 12550 12122
rect 12800 12110 12810 12170
rect 12870 12110 13170 12170
rect 13230 12110 13250 12170
rect 13310 12110 13330 12170
rect 13390 12110 13690 12170
rect 13750 12110 13760 12170
rect 12800 12100 13760 12110
rect 14010 12122 16320 12130
rect 9640 12060 12550 12070
rect 14010 12070 14012 12122
rect 14064 12070 14336 12122
rect 14388 12070 14490 12122
rect 14542 12070 14814 12122
rect 14866 12070 14972 12122
rect 15024 12120 16320 12122
rect 15024 12070 16250 12120
rect 14010 12060 16250 12070
rect 16310 12060 16320 12120
rect 9570 12050 9650 12060
rect 16240 12050 16320 12060
rect 11600 12020 12640 12030
rect 11600 11960 11610 12020
rect 11670 11960 12090 12020
rect 12150 11960 12570 12020
rect 12630 11960 12640 12020
rect 11600 11950 12640 11960
rect 13920 12020 14960 12030
rect 13920 11960 13930 12020
rect 13990 11960 14410 12020
rect 14470 11960 14890 12020
rect 14950 11960 14960 12020
rect 13920 11950 14960 11960
rect 11360 11910 12400 11920
rect 11360 11850 11370 11910
rect 11430 11850 11850 11910
rect 11910 11850 12330 11910
rect 12390 11850 12400 11910
rect 11360 11840 12400 11850
rect 14160 11910 15200 11920
rect 14160 11850 14170 11910
rect 14230 11850 14650 11910
rect 14710 11850 15130 11910
rect 15190 11850 15200 11910
rect 14160 11840 15200 11850
rect 13740 11800 16590 11810
rect 13740 11740 13750 11800
rect 13810 11740 13930 11800
rect 13990 11740 14170 11800
rect 14230 11740 14410 11800
rect 14470 11740 14650 11800
rect 14710 11740 15130 11800
rect 15190 11740 15370 11800
rect 15430 11740 15790 11800
rect 15850 11740 16360 11800
rect 16420 11740 16440 11800
rect 16500 11740 16520 11800
rect 16580 11740 16590 11800
rect 13740 11720 16590 11740
rect 13740 11660 13750 11720
rect 13810 11660 13930 11720
rect 13990 11660 14170 11720
rect 14230 11660 14410 11720
rect 14470 11660 14650 11720
rect 14710 11660 15130 11720
rect 15190 11660 15370 11720
rect 15430 11660 15790 11720
rect 15850 11660 16360 11720
rect 16420 11660 16440 11720
rect 16500 11660 16520 11720
rect 16580 11660 16590 11720
rect 10620 11640 12820 11650
rect 10620 11580 10630 11640
rect 10690 11580 10710 11640
rect 10770 11580 11130 11640
rect 11190 11580 11370 11640
rect 11430 11580 11850 11640
rect 11910 11580 12090 11640
rect 12150 11580 12570 11640
rect 12630 11580 12750 11640
rect 12810 11580 12820 11640
rect 10620 11570 12820 11580
rect 13740 11640 16590 11660
rect 13740 11580 13750 11640
rect 13810 11580 13930 11640
rect 13990 11580 14170 11640
rect 14230 11580 14410 11640
rect 14470 11580 14650 11640
rect 14710 11580 15130 11640
rect 15190 11580 15370 11640
rect 15430 11580 15790 11640
rect 15850 11580 16360 11640
rect 16420 11580 16440 11640
rect 16500 11580 16520 11640
rect 16580 11580 16590 11640
rect 13740 11570 16590 11580
rect 10880 11520 10960 11530
rect 10880 11460 10890 11520
rect 10950 11510 10960 11520
rect 11600 11520 11680 11530
rect 11600 11510 11610 11520
rect 10950 11470 11610 11510
rect 10950 11460 10960 11470
rect 10880 11450 10960 11460
rect 11600 11460 11610 11470
rect 11670 11510 11680 11520
rect 12320 11520 12400 11530
rect 12320 11510 12330 11520
rect 11670 11470 12330 11510
rect 11670 11460 11680 11470
rect 11600 11450 11680 11460
rect 12320 11460 12330 11470
rect 12390 11460 12400 11520
rect 12320 11450 12400 11460
rect 14160 11520 14240 11530
rect 14160 11460 14170 11520
rect 14230 11510 14240 11520
rect 14880 11520 14960 11530
rect 14880 11510 14890 11520
rect 14230 11470 14890 11510
rect 14230 11460 14240 11470
rect 14160 11450 14240 11460
rect 14880 11460 14890 11470
rect 14950 11510 14960 11520
rect 15600 11520 15680 11530
rect 15600 11510 15610 11520
rect 14950 11470 15610 11510
rect 14950 11460 14960 11470
rect 14880 11450 14960 11460
rect 15600 11460 15610 11470
rect 15670 11460 15680 11520
rect 15600 11450 15680 11460
rect 11370 11190 11430 11220
rect 15130 11190 15190 11230
rect 8790 11180 13140 11190
rect 8790 11120 8800 11180
rect 8860 11120 10650 11180
rect 10710 11120 11370 11180
rect 11430 11120 12090 11180
rect 12150 11120 12810 11180
rect 12870 11120 13070 11180
rect 13130 11120 13140 11180
rect 8790 11110 13140 11120
rect 13420 11180 17650 11190
rect 13420 11120 13430 11180
rect 13490 11120 13690 11180
rect 13750 11120 14410 11180
rect 14470 11120 15130 11180
rect 15190 11120 15850 11180
rect 15910 11120 17580 11180
rect 17640 11120 17650 11180
rect 13420 11110 17650 11120
rect 10520 11070 16040 11080
rect 10520 11010 10530 11070
rect 10590 11010 10770 11070
rect 10830 11010 11010 11070
rect 11070 11010 11250 11070
rect 11310 11010 11490 11070
rect 11550 11010 11730 11070
rect 11790 11010 11970 11070
rect 12030 11010 12210 11070
rect 12270 11010 12450 11070
rect 12510 11010 12690 11070
rect 12750 11010 12930 11070
rect 12990 11010 13570 11070
rect 13630 11010 13810 11070
rect 13870 11010 14050 11070
rect 14110 11010 14290 11070
rect 14350 11010 14530 11070
rect 14590 11010 14770 11070
rect 14830 11010 15010 11070
rect 15070 11010 15250 11070
rect 15310 11010 15490 11070
rect 15550 11010 15730 11070
rect 15790 11010 15970 11070
rect 16030 11010 16040 11070
rect 10520 10990 16040 11010
rect 10520 10930 10530 10990
rect 10590 10930 10770 10990
rect 10830 10930 11010 10990
rect 11070 10930 11250 10990
rect 11310 10930 11490 10990
rect 11550 10930 11730 10990
rect 11790 10930 11970 10990
rect 12030 10930 12210 10990
rect 12270 10930 12450 10990
rect 12510 10930 12690 10990
rect 12750 10930 12930 10990
rect 12990 10930 13570 10990
rect 13630 10930 13810 10990
rect 13870 10930 14050 10990
rect 14110 10930 14290 10990
rect 14350 10930 14530 10990
rect 14590 10930 14770 10990
rect 14830 10930 15010 10990
rect 15070 10930 15250 10990
rect 15310 10930 15490 10990
rect 15550 10930 15730 10990
rect 15790 10930 15970 10990
rect 16030 10930 16040 10990
rect 10520 10910 16040 10930
rect 10520 10850 10530 10910
rect 10590 10850 10770 10910
rect 10830 10850 11010 10910
rect 11070 10850 11250 10910
rect 11310 10850 11490 10910
rect 11550 10850 11730 10910
rect 11790 10850 11970 10910
rect 12030 10850 12210 10910
rect 12270 10850 12450 10910
rect 12510 10850 12690 10910
rect 12750 10850 12930 10910
rect 12990 10850 13570 10910
rect 13630 10850 13810 10910
rect 13870 10850 14050 10910
rect 14110 10850 14290 10910
rect 14350 10850 14530 10910
rect 14590 10850 14770 10910
rect 14830 10850 15010 10910
rect 15070 10850 15250 10910
rect 15310 10850 15490 10910
rect 15550 10850 15730 10910
rect 15790 10850 15970 10910
rect 16030 10850 16040 10910
rect 10520 10840 16040 10850
rect 9570 10800 14760 10810
rect 9570 10740 9580 10800
rect 9640 10740 11810 10800
rect 11870 10740 13250 10800
rect 13310 10740 14690 10800
rect 14750 10740 14760 10800
rect 9570 10730 14760 10740
rect 9460 10690 15790 10700
rect 9460 10630 9470 10690
rect 9530 10630 12170 10690
rect 12230 10630 14330 10690
rect 14390 10630 15720 10690
rect 15780 10630 15790 10690
rect 9460 10620 15790 10630
rect 12520 10580 16320 10590
rect 12520 10520 12530 10580
rect 12590 10520 13970 10580
rect 14030 10520 15250 10580
rect 15310 10520 16250 10580
rect 16310 10520 16320 10580
rect 12520 10510 16320 10520
rect 12880 10470 16230 10480
rect 12880 10410 12890 10470
rect 12950 10410 13610 10470
rect 13670 10410 16160 10470
rect 16220 10410 16230 10470
rect 12880 10400 16230 10410
rect 11900 10360 14660 10370
rect 11960 10300 12080 10360
rect 12140 10300 12260 10360
rect 12320 10300 12440 10360
rect 12500 10300 12620 10360
rect 12680 10300 12800 10360
rect 12860 10300 12980 10360
rect 13040 10300 13160 10360
rect 13220 10300 13340 10360
rect 13400 10300 13430 10360
rect 13490 10300 13520 10360
rect 13580 10300 13700 10360
rect 13760 10300 13880 10360
rect 13940 10300 14060 10360
rect 14120 10300 14240 10360
rect 14300 10300 14420 10360
rect 14480 10300 14600 10360
rect 11900 10290 14660 10300
rect 15590 10160 15910 10170
rect 15590 10100 15600 10160
rect 15660 10100 15840 10160
rect 15900 10100 15910 10160
rect 15590 10090 15910 10100
rect 15240 9820 15320 9830
rect 15240 9760 15250 9820
rect 15310 9810 15320 9820
rect 15710 9820 15790 9830
rect 15710 9810 15720 9820
rect 15310 9770 15720 9810
rect 15310 9760 15320 9770
rect 15240 9750 15320 9760
rect 15710 9760 15720 9770
rect 15780 9760 15790 9820
rect 15710 9750 15790 9760
rect 11620 9620 16010 9630
rect 11620 9560 11630 9620
rect 11690 9560 11990 9620
rect 12050 9560 12350 9620
rect 12410 9560 12710 9620
rect 12770 9560 13070 9620
rect 13130 9560 13430 9620
rect 13490 9560 13790 9620
rect 13850 9560 14150 9620
rect 14210 9560 14510 9620
rect 14570 9560 14870 9620
rect 14930 9560 15500 9620
rect 15560 9560 15940 9620
rect 16000 9560 16010 9620
rect 11620 9540 16010 9560
rect 11620 9480 11630 9540
rect 11690 9480 11990 9540
rect 12050 9480 12350 9540
rect 12410 9480 12710 9540
rect 12770 9480 13070 9540
rect 13130 9480 13430 9540
rect 13490 9480 13790 9540
rect 13850 9480 14150 9540
rect 14210 9480 14510 9540
rect 14570 9480 14870 9540
rect 14930 9480 15500 9540
rect 15560 9480 15940 9540
rect 16000 9480 16010 9540
rect 11620 9460 16010 9480
rect 11620 9400 11630 9460
rect 11690 9400 11990 9460
rect 12050 9400 12350 9460
rect 12410 9400 12710 9460
rect 12770 9400 13070 9460
rect 13130 9400 13430 9460
rect 13490 9400 13790 9460
rect 13850 9400 14150 9460
rect 14210 9400 14510 9460
rect 14570 9400 14870 9460
rect 14930 9400 15500 9460
rect 15560 9400 15940 9460
rect 16000 9400 16010 9460
rect 11620 9390 16010 9400
rect 8790 9300 8800 9360
rect 8860 9350 14754 9360
rect 8860 9300 11808 9350
rect 8790 9298 11808 9300
rect 11860 9298 11918 9350
rect 11970 9298 12028 9350
rect 12080 9298 12138 9350
rect 12190 9298 12248 9350
rect 12300 9298 12358 9350
rect 12410 9298 12468 9350
rect 12520 9298 12578 9350
rect 12630 9298 12688 9350
rect 12740 9298 12798 9350
rect 12850 9298 13708 9350
rect 13760 9298 13818 9350
rect 13870 9298 13928 9350
rect 13980 9298 14038 9350
rect 14090 9298 14148 9350
rect 14200 9298 14258 9350
rect 14310 9298 14368 9350
rect 14420 9298 14478 9350
rect 14530 9298 14588 9350
rect 14640 9298 14698 9350
rect 14750 9298 14754 9350
rect 8790 9290 14754 9298
rect 11630 9020 14930 9030
rect 11630 8960 11640 9020
rect 11700 8960 11860 9020
rect 11920 8960 12080 9020
rect 12140 8960 12300 9020
rect 12360 8960 12520 9020
rect 12580 8960 12740 9020
rect 12800 8960 12960 9020
rect 13020 8960 13540 9020
rect 13600 8960 13760 9020
rect 13820 8960 13980 9020
rect 14040 8960 14200 9020
rect 14260 8960 14420 9020
rect 14480 8960 14640 9020
rect 14700 8960 14860 9020
rect 14920 8960 14930 9020
rect 11630 8950 14930 8960
rect 9680 8910 12920 8920
rect 9680 8850 9690 8910
rect 9750 8850 11750 8910
rect 11810 8850 11970 8910
rect 12030 8850 12190 8910
rect 12250 8850 12410 8910
rect 12470 8850 12630 8910
rect 12690 8850 12850 8910
rect 12910 8850 12920 8910
rect 9680 8840 12920 8850
rect 13640 8900 14820 8910
rect 13640 8840 13650 8900
rect 13710 8840 13870 8900
rect 13930 8840 14090 8900
rect 14150 8840 14310 8900
rect 14370 8840 14530 8900
rect 14590 8840 14750 8900
rect 14810 8840 14820 8900
rect 13640 8820 14820 8840
rect 13640 8760 13650 8820
rect 13710 8760 13870 8820
rect 13930 8760 14090 8820
rect 14150 8760 14310 8820
rect 14370 8760 14530 8820
rect 14590 8760 14750 8820
rect 14810 8760 14820 8820
rect 13640 8740 14820 8760
rect 13640 8680 13650 8740
rect 13710 8680 13870 8740
rect 13930 8680 14090 8740
rect 14150 8680 14310 8740
rect 14370 8680 14530 8740
rect 14590 8680 14750 8740
rect 14810 8680 14820 8740
rect 13640 8670 14820 8680
<< via2 >>
rect 18200 18790 18260 18850
rect 18660 18090 18720 18150
rect 18130 17390 18190 17450
rect 18800 16690 18860 16750
rect 19000 15990 19060 16050
rect 18800 15290 18860 15350
<< metal3 >>
rect 19120 18870 19580 19040
rect 19820 18870 20280 19040
rect 20520 18870 20980 19040
rect 21220 18870 21680 19040
rect 21920 18870 22380 19040
rect 22620 18870 23080 19040
rect 23320 18870 23780 19040
rect 24020 18870 24480 19040
rect 24720 18870 25180 19040
rect 25420 18870 25880 19040
rect 19120 18860 25880 18870
rect 18190 18850 25880 18860
rect 18190 18790 18200 18850
rect 18260 18790 25880 18850
rect 18190 18780 25880 18790
rect 19120 18770 25880 18780
rect 19120 18580 19580 18770
rect 19820 18580 20280 18770
rect 20520 18580 20980 18770
rect 21220 18580 21680 18770
rect 21920 18580 22380 18770
rect 22620 18580 23080 18770
rect 23320 18580 23780 18770
rect 24020 18580 24480 18770
rect 24720 18580 25180 18770
rect 25420 18580 25880 18770
rect 25600 18340 25700 18580
rect 19120 18170 19580 18340
rect 19820 18170 20280 18340
rect 20520 18170 20980 18340
rect 21220 18170 21680 18340
rect 21920 18170 22380 18340
rect 22620 18170 23080 18340
rect 23320 18170 23780 18340
rect 24020 18170 24480 18340
rect 24720 18170 25180 18340
rect 25420 18170 25880 18340
rect 18640 18160 18740 18170
rect 18640 18080 18650 18160
rect 18730 18080 18740 18160
rect 18640 18070 18740 18080
rect 19120 18070 25880 18170
rect 19120 17880 19580 18070
rect 19820 17880 20280 18070
rect 20520 17880 20980 18070
rect 21220 17880 21680 18070
rect 21920 17880 22380 18070
rect 22620 17880 23080 18070
rect 23320 17880 23780 18070
rect 24020 17880 24480 18070
rect 24720 17880 25180 18070
rect 25420 17880 25880 18070
rect 19120 17470 19580 17640
rect 19820 17470 20280 17640
rect 20520 17470 20980 17640
rect 21220 17470 21680 17640
rect 21920 17470 22380 17640
rect 22620 17470 23080 17640
rect 23320 17470 23780 17640
rect 24020 17470 24480 17640
rect 24720 17470 25180 17640
rect 25420 17470 25880 17640
rect 19120 17460 25880 17470
rect 18120 17450 25880 17460
rect 18120 17390 18130 17450
rect 18190 17390 25880 17450
rect 18120 17380 25880 17390
rect 19120 17370 25880 17380
rect 19120 17180 19580 17370
rect 19820 17180 20280 17370
rect 20520 17180 20980 17370
rect 21220 17180 21680 17370
rect 21920 17180 22380 17370
rect 22620 17180 23080 17370
rect 23320 17180 23780 17370
rect 24020 17180 24480 17370
rect 24720 17180 25180 17370
rect 25420 17180 25880 17370
rect 25600 16940 25700 17180
rect 19120 16770 19580 16940
rect 19820 16770 20280 16940
rect 20520 16770 20980 16940
rect 21220 16770 21680 16940
rect 21920 16770 22380 16940
rect 22620 16770 23080 16940
rect 23320 16770 23780 16940
rect 24020 16770 24480 16940
rect 24720 16770 25180 16940
rect 25420 16770 25880 16940
rect 18780 16760 18880 16770
rect 18780 16680 18790 16760
rect 18870 16680 18880 16760
rect 18780 16670 18880 16680
rect 19120 16670 25880 16770
rect 19120 16480 19580 16670
rect 19820 16480 20280 16670
rect 20520 16480 20980 16670
rect 21220 16480 21680 16670
rect 21920 16480 22380 16670
rect 22620 16480 23080 16670
rect 23320 16480 23780 16670
rect 24020 16480 24480 16670
rect 24720 16480 25180 16670
rect 25420 16480 25880 16670
rect 19120 16070 19580 16240
rect 19820 16070 20280 16240
rect 20520 16070 20980 16240
rect 21220 16070 21680 16240
rect 21920 16070 22380 16240
rect 22620 16070 23080 16240
rect 23320 16070 23780 16240
rect 24020 16070 24480 16240
rect 24720 16070 25180 16240
rect 25420 16070 25880 16240
rect 19120 16060 25880 16070
rect 18990 16050 25880 16060
rect 18990 15990 19000 16050
rect 19060 15990 25880 16050
rect 18990 15980 25880 15990
rect 19120 15970 25880 15980
rect 19120 15780 19580 15970
rect 19820 15780 20280 15970
rect 20520 15780 20980 15970
rect 21220 15780 21680 15970
rect 21920 15780 22380 15970
rect 22620 15780 23080 15970
rect 23320 15780 23780 15970
rect 24020 15780 24480 15970
rect 24720 15780 25180 15970
rect 25420 15780 25880 15970
rect 25600 15540 25700 15780
rect 19120 15370 19580 15540
rect 19820 15370 20280 15540
rect 20520 15370 20980 15540
rect 21220 15370 21680 15540
rect 21920 15370 22380 15540
rect 22620 15370 23080 15540
rect 23320 15370 23780 15540
rect 24020 15370 24480 15540
rect 24720 15370 25180 15540
rect 25420 15370 25880 15540
rect 18780 15360 18880 15370
rect 18780 15280 18790 15360
rect 18870 15280 18880 15360
rect 18780 15270 18880 15280
rect 19120 15270 25880 15370
rect 19120 15080 19580 15270
rect 19820 15080 20280 15270
rect 20520 15080 20980 15270
rect 21220 15080 21680 15270
rect 21920 15080 22380 15270
rect 22620 15080 23080 15270
rect 23320 15080 23780 15270
rect 24020 15080 24480 15270
rect 24720 15080 25180 15270
rect 25420 15080 25880 15270
<< via3 >>
rect 18650 18150 18730 18160
rect 18650 18090 18660 18150
rect 18660 18090 18720 18150
rect 18720 18090 18730 18150
rect 18650 18080 18730 18090
rect 18790 16750 18870 16760
rect 18790 16690 18800 16750
rect 18800 16690 18860 16750
rect 18860 16690 18870 16750
rect 18790 16680 18870 16690
rect 18790 15350 18870 15360
rect 18790 15290 18800 15350
rect 18800 15290 18860 15350
rect 18860 15290 18870 15350
rect 18790 15280 18870 15290
<< mimcap >>
rect 19150 18860 19550 19010
rect 19150 18780 19320 18860
rect 19400 18780 19550 18860
rect 19150 18610 19550 18780
rect 19850 18860 20250 19010
rect 19850 18780 20010 18860
rect 20090 18780 20250 18860
rect 19850 18610 20250 18780
rect 20550 18860 20950 19010
rect 20550 18780 20710 18860
rect 20790 18780 20950 18860
rect 20550 18610 20950 18780
rect 21250 18860 21650 19010
rect 21250 18780 21410 18860
rect 21490 18780 21650 18860
rect 21250 18610 21650 18780
rect 21950 18860 22350 19010
rect 21950 18780 22110 18860
rect 22190 18780 22350 18860
rect 21950 18610 22350 18780
rect 22650 18860 23050 19010
rect 22650 18780 22810 18860
rect 22890 18780 23050 18860
rect 22650 18610 23050 18780
rect 23350 18860 23750 19010
rect 23350 18780 23510 18860
rect 23590 18780 23750 18860
rect 23350 18610 23750 18780
rect 24050 18860 24450 19010
rect 24050 18780 24210 18860
rect 24290 18780 24450 18860
rect 24050 18610 24450 18780
rect 24750 18860 25150 19010
rect 24750 18780 24910 18860
rect 24990 18780 25150 18860
rect 24750 18610 25150 18780
rect 25450 18860 25850 19010
rect 25450 18780 25610 18860
rect 25690 18780 25850 18860
rect 25450 18610 25850 18780
rect 19150 18160 19550 18310
rect 19150 18080 19320 18160
rect 19400 18080 19550 18160
rect 19150 17910 19550 18080
rect 19850 18160 20250 18310
rect 19850 18080 20010 18160
rect 20090 18080 20250 18160
rect 19850 17910 20250 18080
rect 20550 18160 20950 18310
rect 20550 18080 20710 18160
rect 20790 18080 20950 18160
rect 20550 17910 20950 18080
rect 21250 18160 21650 18310
rect 21250 18080 21410 18160
rect 21490 18080 21650 18160
rect 21250 17910 21650 18080
rect 21950 18160 22350 18310
rect 21950 18080 22110 18160
rect 22190 18080 22350 18160
rect 21950 17910 22350 18080
rect 22650 18160 23050 18310
rect 22650 18080 22810 18160
rect 22890 18080 23050 18160
rect 22650 17910 23050 18080
rect 23350 18160 23750 18310
rect 23350 18080 23510 18160
rect 23590 18080 23750 18160
rect 23350 17910 23750 18080
rect 24050 18160 24450 18310
rect 24050 18080 24210 18160
rect 24290 18080 24450 18160
rect 24050 17910 24450 18080
rect 24750 18160 25150 18310
rect 24750 18080 24910 18160
rect 24990 18080 25150 18160
rect 24750 17910 25150 18080
rect 25450 18160 25850 18310
rect 25450 18080 25610 18160
rect 25690 18080 25850 18160
rect 25450 17910 25850 18080
rect 19150 17460 19550 17610
rect 19150 17380 19320 17460
rect 19400 17380 19550 17460
rect 19150 17210 19550 17380
rect 19850 17460 20250 17610
rect 19850 17380 20010 17460
rect 20090 17380 20250 17460
rect 19850 17210 20250 17380
rect 20550 17460 20950 17610
rect 20550 17380 20710 17460
rect 20790 17380 20950 17460
rect 20550 17210 20950 17380
rect 21250 17460 21650 17610
rect 21250 17380 21410 17460
rect 21490 17380 21650 17460
rect 21250 17210 21650 17380
rect 21950 17460 22350 17610
rect 21950 17380 22110 17460
rect 22190 17380 22350 17460
rect 21950 17210 22350 17380
rect 22650 17460 23050 17610
rect 22650 17380 22810 17460
rect 22890 17380 23050 17460
rect 22650 17210 23050 17380
rect 23350 17460 23750 17610
rect 23350 17380 23510 17460
rect 23590 17380 23750 17460
rect 23350 17210 23750 17380
rect 24050 17460 24450 17610
rect 24050 17380 24210 17460
rect 24290 17380 24450 17460
rect 24050 17210 24450 17380
rect 24750 17460 25150 17610
rect 24750 17380 24910 17460
rect 24990 17380 25150 17460
rect 24750 17210 25150 17380
rect 25450 17460 25850 17610
rect 25450 17380 25610 17460
rect 25690 17380 25850 17460
rect 25450 17210 25850 17380
rect 19150 16760 19550 16910
rect 19150 16680 19320 16760
rect 19400 16680 19550 16760
rect 19150 16510 19550 16680
rect 19850 16760 20250 16910
rect 19850 16680 20010 16760
rect 20090 16680 20250 16760
rect 19850 16510 20250 16680
rect 20550 16760 20950 16910
rect 20550 16680 20710 16760
rect 20790 16680 20950 16760
rect 20550 16510 20950 16680
rect 21250 16760 21650 16910
rect 21250 16680 21410 16760
rect 21490 16680 21650 16760
rect 21250 16510 21650 16680
rect 21950 16760 22350 16910
rect 21950 16680 22110 16760
rect 22190 16680 22350 16760
rect 21950 16510 22350 16680
rect 22650 16760 23050 16910
rect 22650 16680 22810 16760
rect 22890 16680 23050 16760
rect 22650 16510 23050 16680
rect 23350 16760 23750 16910
rect 23350 16680 23510 16760
rect 23590 16680 23750 16760
rect 23350 16510 23750 16680
rect 24050 16760 24450 16910
rect 24050 16680 24210 16760
rect 24290 16680 24450 16760
rect 24050 16510 24450 16680
rect 24750 16760 25150 16910
rect 24750 16680 24910 16760
rect 24990 16680 25150 16760
rect 24750 16510 25150 16680
rect 25450 16760 25850 16910
rect 25450 16680 25610 16760
rect 25690 16680 25850 16760
rect 25450 16510 25850 16680
rect 19150 16060 19550 16210
rect 19150 15980 19320 16060
rect 19400 15980 19550 16060
rect 19150 15810 19550 15980
rect 19850 16060 20250 16210
rect 19850 15980 20010 16060
rect 20090 15980 20250 16060
rect 19850 15810 20250 15980
rect 20550 16060 20950 16210
rect 20550 15980 20710 16060
rect 20790 15980 20950 16060
rect 20550 15810 20950 15980
rect 21250 16060 21650 16210
rect 21250 15980 21410 16060
rect 21490 15980 21650 16060
rect 21250 15810 21650 15980
rect 21950 16060 22350 16210
rect 21950 15980 22110 16060
rect 22190 15980 22350 16060
rect 21950 15810 22350 15980
rect 22650 16060 23050 16210
rect 22650 15980 22810 16060
rect 22890 15980 23050 16060
rect 22650 15810 23050 15980
rect 23350 16060 23750 16210
rect 23350 15980 23510 16060
rect 23590 15980 23750 16060
rect 23350 15810 23750 15980
rect 24050 16060 24450 16210
rect 24050 15980 24210 16060
rect 24290 15980 24450 16060
rect 24050 15810 24450 15980
rect 24750 16060 25150 16210
rect 24750 15980 24910 16060
rect 24990 15980 25150 16060
rect 24750 15810 25150 15980
rect 25450 16060 25850 16210
rect 25450 15980 25610 16060
rect 25690 15980 25850 16060
rect 25450 15810 25850 15980
rect 19150 15360 19550 15510
rect 19150 15280 19320 15360
rect 19400 15280 19550 15360
rect 19150 15110 19550 15280
rect 19850 15360 20250 15510
rect 19850 15280 20010 15360
rect 20090 15280 20250 15360
rect 19850 15110 20250 15280
rect 20550 15360 20950 15510
rect 20550 15280 20710 15360
rect 20790 15280 20950 15360
rect 20550 15110 20950 15280
rect 21250 15360 21650 15510
rect 21250 15280 21410 15360
rect 21490 15280 21650 15360
rect 21250 15110 21650 15280
rect 21950 15360 22350 15510
rect 21950 15280 22110 15360
rect 22190 15280 22350 15360
rect 21950 15110 22350 15280
rect 22650 15360 23050 15510
rect 22650 15280 22810 15360
rect 22890 15280 23050 15360
rect 22650 15110 23050 15280
rect 23350 15360 23750 15510
rect 23350 15280 23510 15360
rect 23590 15280 23750 15360
rect 23350 15110 23750 15280
rect 24050 15360 24450 15510
rect 24050 15280 24210 15360
rect 24290 15280 24450 15360
rect 24050 15110 24450 15280
rect 24750 15360 25150 15510
rect 24750 15280 24910 15360
rect 24990 15280 25150 15360
rect 24750 15110 25150 15280
rect 25450 15360 25850 15510
rect 25450 15280 25610 15360
rect 25690 15280 25850 15360
rect 25450 15110 25850 15280
<< mimcapcontact >>
rect 19320 18780 19400 18860
rect 20010 18780 20090 18860
rect 20710 18780 20790 18860
rect 21410 18780 21490 18860
rect 22110 18780 22190 18860
rect 22810 18780 22890 18860
rect 23510 18780 23590 18860
rect 24210 18780 24290 18860
rect 24910 18780 24990 18860
rect 25610 18780 25690 18860
rect 19320 18080 19400 18160
rect 20010 18080 20090 18160
rect 20710 18080 20790 18160
rect 21410 18080 21490 18160
rect 22110 18080 22190 18160
rect 22810 18080 22890 18160
rect 23510 18080 23590 18160
rect 24210 18080 24290 18160
rect 24910 18080 24990 18160
rect 25610 18080 25690 18160
rect 19320 17380 19400 17460
rect 20010 17380 20090 17460
rect 20710 17380 20790 17460
rect 21410 17380 21490 17460
rect 22110 17380 22190 17460
rect 22810 17380 22890 17460
rect 23510 17380 23590 17460
rect 24210 17380 24290 17460
rect 24910 17380 24990 17460
rect 25610 17380 25690 17460
rect 19320 16680 19400 16760
rect 20010 16680 20090 16760
rect 20710 16680 20790 16760
rect 21410 16680 21490 16760
rect 22110 16680 22190 16760
rect 22810 16680 22890 16760
rect 23510 16680 23590 16760
rect 24210 16680 24290 16760
rect 24910 16680 24990 16760
rect 25610 16680 25690 16760
rect 19320 15980 19400 16060
rect 20010 15980 20090 16060
rect 20710 15980 20790 16060
rect 21410 15980 21490 16060
rect 22110 15980 22190 16060
rect 22810 15980 22890 16060
rect 23510 15980 23590 16060
rect 24210 15980 24290 16060
rect 24910 15980 24990 16060
rect 25610 15980 25690 16060
rect 19320 15280 19400 15360
rect 20010 15280 20090 15360
rect 20710 15280 20790 15360
rect 21410 15280 21490 15360
rect 22110 15280 22190 15360
rect 22810 15280 22890 15360
rect 23510 15280 23590 15360
rect 24210 15280 24290 15360
rect 24910 15280 24990 15360
rect 25610 15280 25690 15360
<< metal4 >>
rect 19310 18860 25700 18870
rect 19310 18780 19320 18860
rect 19400 18780 20010 18860
rect 20090 18780 20710 18860
rect 20790 18780 21410 18860
rect 21490 18780 22110 18860
rect 22190 18780 22810 18860
rect 22890 18780 23510 18860
rect 23590 18780 24210 18860
rect 24290 18780 24910 18860
rect 24990 18780 25610 18860
rect 25690 18780 25700 18860
rect 19310 18770 25700 18780
rect 25600 18170 25700 18770
rect 18640 18160 25700 18170
rect 18640 18080 18650 18160
rect 18730 18080 19320 18160
rect 19400 18080 20010 18160
rect 20090 18080 20710 18160
rect 20790 18080 21410 18160
rect 21490 18080 22110 18160
rect 22190 18080 22810 18160
rect 22890 18080 23510 18160
rect 23590 18080 24210 18160
rect 24290 18080 24910 18160
rect 24990 18080 25610 18160
rect 25690 18080 25700 18160
rect 18640 18070 25700 18080
rect 19310 17460 25700 17470
rect 19310 17380 19320 17460
rect 19400 17380 20010 17460
rect 20090 17380 20710 17460
rect 20790 17380 21410 17460
rect 21490 17380 22110 17460
rect 22190 17380 22810 17460
rect 22890 17380 23510 17460
rect 23590 17380 24210 17460
rect 24290 17380 24910 17460
rect 24990 17380 25610 17460
rect 25690 17380 25700 17460
rect 19310 17370 25700 17380
rect 25600 16770 25700 17370
rect 18780 16760 25700 16770
rect 18780 16680 18790 16760
rect 18870 16680 19320 16760
rect 19400 16680 20010 16760
rect 20090 16680 20710 16760
rect 20790 16680 21410 16760
rect 21490 16680 22110 16760
rect 22190 16680 22810 16760
rect 22890 16680 23510 16760
rect 23590 16680 24210 16760
rect 24290 16680 24910 16760
rect 24990 16680 25610 16760
rect 25690 16680 25700 16760
rect 18780 16670 25700 16680
rect 19310 16060 25700 16070
rect 19310 15980 19320 16060
rect 19400 15980 20010 16060
rect 20090 15980 20710 16060
rect 20790 15980 21410 16060
rect 21490 15980 22110 16060
rect 22190 15980 22810 16060
rect 22890 15980 23510 16060
rect 23590 15980 24210 16060
rect 24290 15980 24910 16060
rect 24990 15980 25610 16060
rect 25690 15980 25700 16060
rect 19310 15970 25700 15980
rect 25600 15370 25700 15970
rect 18780 15360 25700 15370
rect 18780 15280 18790 15360
rect 18870 15280 19320 15360
rect 19400 15280 20010 15360
rect 20090 15280 20710 15360
rect 20790 15280 21410 15360
rect 21490 15280 22110 15360
rect 22190 15280 22810 15360
rect 22890 15280 23510 15360
rect 23590 15280 24210 15360
rect 24290 15280 24910 15360
rect 24990 15280 25610 15360
rect 25690 15280 25700 15360
rect 18780 15270 25700 15280
<< labels >>
flabel metal2 13290 9290 13290 9290 5 FreeSans 1600 0 0 -800 PFET_GATE
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
