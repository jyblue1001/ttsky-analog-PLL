magic
tech sky130A
magscale 1 2
timestamp 1757393363
<< nwell >>
rect 54817 19209 57503 19733
<< nsubdiff >>
rect 54853 19663 54949 19697
rect 57371 19663 57467 19697
rect 54853 19601 54887 19663
rect 57433 19601 57467 19663
rect 54853 19279 54887 19341
rect 57433 19279 57467 19341
rect 54853 19245 54949 19279
rect 57371 19245 57467 19279
<< nsubdiffcont >>
rect 54949 19663 57371 19697
rect 54853 19341 54887 19601
rect 57433 19341 57467 19601
rect 54949 19245 57371 19279
<< xpolycontact >>
rect 54992 19436 55424 19506
rect 56896 19436 57328 19506
<< xpolyres >>
rect 55424 19436 56896 19506
<< locali >>
rect 56120 19697 56200 19700
rect 54853 19663 54949 19697
rect 57371 19663 57467 19697
rect 54853 19601 54887 19663
rect 56120 19640 56140 19663
rect 56180 19640 56200 19663
rect 56120 19620 56200 19640
rect 57433 19601 57467 19663
rect 54853 19279 54887 19341
rect 57433 19279 57467 19341
rect 54853 19245 54949 19279
rect 57371 19245 57467 19279
<< viali >>
rect 56140 19663 56180 19680
rect 56140 19640 56180 19663
rect 55010 19452 55407 19490
rect 56913 19452 57310 19490
<< metal1 >>
rect 56120 19690 56200 19700
rect 56120 19630 56130 19690
rect 56190 19630 56200 19690
rect 56120 19620 56200 19630
rect 54990 19500 55420 19510
rect 54990 19440 55000 19500
rect 55410 19440 55420 19500
rect 54990 19430 55420 19440
rect 56900 19500 57330 19510
rect 56900 19440 56910 19500
rect 57320 19440 57330 19500
rect 56900 19430 57330 19440
rect 65990 19500 66090 19520
rect 65990 19440 66010 19500
rect 66070 19440 66090 19500
rect 65990 19420 66090 19440
<< via1 >>
rect 56130 19680 56190 19690
rect 56130 19640 56140 19680
rect 56140 19640 56180 19680
rect 56180 19640 56190 19680
rect 56130 19630 56190 19640
rect 55000 19490 55410 19500
rect 55000 19452 55010 19490
rect 55010 19452 55407 19490
rect 55407 19452 55410 19490
rect 55000 19440 55410 19452
rect 56910 19490 57320 19500
rect 56910 19452 56913 19490
rect 56913 19452 57310 19490
rect 57310 19452 57320 19490
rect 56910 19440 57320 19452
rect 66010 19440 66070 19500
<< metal2 >>
rect 47720 19790 63410 19810
rect 47720 19720 62820 19790
rect 62890 19720 63320 19790
rect 63390 19720 63410 19790
rect 47720 19700 63410 19720
rect 56120 19690 56200 19700
rect 56120 19630 56130 19690
rect 56190 19630 56200 19690
rect 56120 19620 56200 19630
rect 48920 19510 49020 19520
rect 65990 19510 66090 19520
rect 48920 19500 55420 19510
rect 48920 19440 48940 19500
rect 49000 19440 55000 19500
rect 55410 19440 55420 19500
rect 48920 19430 55420 19440
rect 56900 19500 66090 19510
rect 56900 19440 56910 19500
rect 57320 19440 66010 19500
rect 66070 19440 66090 19500
rect 56900 19430 66090 19440
rect 48920 19420 49020 19430
rect 65990 19420 66090 19430
<< via2 >>
rect 62820 19720 62890 19790
rect 63320 19720 63390 19790
rect 48940 19440 49000 19500
rect 66010 19440 66070 19500
<< metal3 >>
rect 48920 20050 62940 32110
rect 63270 20050 66090 32110
rect 48920 19500 49020 20050
rect 62800 19790 62910 19810
rect 62800 19720 62820 19790
rect 62890 19720 62910 19790
rect 62800 19700 62910 19720
rect 63300 19790 63410 19810
rect 63300 19720 63320 19790
rect 63390 19720 63410 19790
rect 63300 19700 63410 19720
rect 48920 19440 48940 19500
rect 49000 19440 49020 19500
rect 48920 19420 49020 19440
rect 65990 19500 66090 20050
rect 65990 19440 66010 19500
rect 66070 19440 66090 19500
rect 65990 19420 66090 19440
<< via3 >>
rect 62820 19720 62890 19790
rect 63320 19720 63390 19790
<< mimcap >>
rect 48950 20170 62910 32080
rect 48950 20100 62820 20170
rect 62890 20100 62910 20170
rect 48950 20080 62910 20100
rect 63300 20170 66060 32080
rect 63300 20100 63320 20170
rect 63390 20100 66060 20170
rect 63300 20080 66060 20100
<< mimcapcontact >>
rect 62820 20100 62890 20170
rect 63320 20100 63390 20170
<< metal4 >>
rect 62800 20170 62910 20180
rect 62800 20100 62820 20170
rect 62890 20100 62910 20170
rect 62800 19790 62910 20100
rect 62800 19720 62820 19790
rect 62890 19720 62910 19790
rect 62800 19700 62910 19720
rect 63300 20170 63410 20180
rect 63300 20100 63320 20170
rect 63390 20100 63410 20170
rect 63300 19790 63410 20100
rect 63300 19720 63320 19790
rect 63390 19720 63410 19790
rect 63300 19700 63410 19720
<< end >>
