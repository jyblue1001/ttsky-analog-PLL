magic
tech sky130A
timestamp 1757393487
<< nwell >>
rect 21565 3235 24055 3855
rect 24695 3250 26305 3540
<< nmos >>
rect 21665 3945 21680 4045
rect 21720 3945 21735 4045
rect 21925 3945 21940 4045
rect 21980 3945 21995 4045
rect 22115 3945 22130 4045
rect 22170 3945 22185 4045
rect 22375 3945 22390 4045
rect 22430 3945 22445 4045
rect 22630 3945 22645 4045
rect 22795 3945 22810 4045
rect 22960 3945 22975 4045
rect 23240 3945 23255 4045
rect 23435 3945 23450 4045
rect 23630 3945 23645 4045
rect 23775 3945 23790 4045
rect 23970 3945 23985 4045
rect 24715 3820 24775 4020
rect 24825 3820 24885 4020
rect 24935 3820 24995 4020
rect 25045 3820 25105 4020
rect 25255 3820 25315 4020
rect 25365 3820 25425 4020
rect 25475 3820 25535 4020
rect 25585 3820 25645 4020
rect 25795 3820 25855 4020
rect 25905 3820 25965 4020
rect 26015 3820 26075 4020
rect 26125 3820 26185 4020
rect 21665 3045 21680 3145
rect 21720 3045 21735 3145
rect 21925 3045 21940 3145
rect 21980 3045 21995 3145
rect 22115 3045 22130 3145
rect 22170 3045 22185 3145
rect 22375 3045 22390 3145
rect 22430 3045 22445 3145
rect 22635 3045 22650 3145
rect 22690 3045 22705 3145
rect 22855 3045 22870 3145
rect 23020 3045 23035 3145
rect 23240 3045 23255 3145
rect 23435 3045 23450 3145
rect 23630 3045 23645 3145
rect 23775 3045 23790 3145
<< pmos >>
rect 21665 3635 21680 3835
rect 21720 3635 21735 3835
rect 21925 3635 21940 3835
rect 21980 3635 21995 3835
rect 22115 3635 22130 3835
rect 22170 3635 22185 3835
rect 22375 3635 22390 3835
rect 22430 3635 22445 3835
rect 22630 3635 22645 3835
rect 22795 3635 22810 3835
rect 22960 3635 22975 3835
rect 23240 3635 23255 3835
rect 23435 3635 23450 3835
rect 23630 3635 23645 3835
rect 23775 3635 23790 3835
rect 21665 3255 21680 3455
rect 21720 3255 21735 3455
rect 21925 3255 21940 3455
rect 21980 3255 21995 3455
rect 22115 3255 22130 3455
rect 22170 3255 22185 3455
rect 22375 3255 22390 3455
rect 22430 3255 22445 3455
rect 22635 3255 22650 3455
rect 22690 3255 22705 3455
rect 22855 3255 22870 3455
rect 23020 3255 23035 3455
rect 23240 3255 23255 3455
rect 23435 3255 23450 3455
rect 23630 3255 23645 3455
rect 23775 3255 23790 3455
rect 23970 3255 23985 3455
rect 24815 3270 24875 3470
rect 24925 3270 24985 3470
rect 25035 3270 25095 3470
rect 25145 3270 25205 3470
rect 25255 3270 25315 3470
rect 25365 3270 25425 3470
rect 25575 3270 25635 3470
rect 25685 3270 25745 3470
rect 25795 3270 25855 3470
rect 25905 3270 25965 3470
rect 26015 3270 26075 3470
rect 26125 3270 26185 3470
<< ndiff >>
rect 21625 4030 21665 4045
rect 21625 4010 21635 4030
rect 21655 4010 21665 4030
rect 21625 3980 21665 4010
rect 21625 3960 21635 3980
rect 21655 3960 21665 3980
rect 21625 3945 21665 3960
rect 21680 4030 21720 4045
rect 21680 4010 21690 4030
rect 21710 4010 21720 4030
rect 21680 3980 21720 4010
rect 21680 3960 21690 3980
rect 21710 3960 21720 3980
rect 21680 3945 21720 3960
rect 21735 4030 21775 4045
rect 21735 4010 21745 4030
rect 21765 4010 21775 4030
rect 21735 3980 21775 4010
rect 21735 3960 21745 3980
rect 21765 3960 21775 3980
rect 21735 3945 21775 3960
rect 21885 4030 21925 4045
rect 21885 4010 21895 4030
rect 21915 4010 21925 4030
rect 21885 3980 21925 4010
rect 21885 3960 21895 3980
rect 21915 3960 21925 3980
rect 21885 3945 21925 3960
rect 21940 4030 21980 4045
rect 21940 4010 21950 4030
rect 21970 4010 21980 4030
rect 21940 3980 21980 4010
rect 21940 3960 21950 3980
rect 21970 3960 21980 3980
rect 21940 3945 21980 3960
rect 21995 4030 22035 4045
rect 22075 4030 22115 4045
rect 21995 4010 22005 4030
rect 22025 4010 22035 4030
rect 22075 4010 22085 4030
rect 22105 4010 22115 4030
rect 21995 3980 22035 4010
rect 22075 3980 22115 4010
rect 21995 3960 22005 3980
rect 22025 3960 22035 3980
rect 22075 3960 22085 3980
rect 22105 3960 22115 3980
rect 21995 3945 22035 3960
rect 22075 3945 22115 3960
rect 22130 4030 22170 4045
rect 22130 4010 22140 4030
rect 22160 4010 22170 4030
rect 22130 3980 22170 4010
rect 22130 3960 22140 3980
rect 22160 3960 22170 3980
rect 22130 3945 22170 3960
rect 22185 4030 22225 4045
rect 22185 4010 22195 4030
rect 22215 4010 22225 4030
rect 22185 3980 22225 4010
rect 22185 3960 22195 3980
rect 22215 3960 22225 3980
rect 22185 3945 22225 3960
rect 22335 4030 22375 4045
rect 22335 4010 22345 4030
rect 22365 4010 22375 4030
rect 22335 3980 22375 4010
rect 22335 3960 22345 3980
rect 22365 3960 22375 3980
rect 22335 3945 22375 3960
rect 22390 4030 22430 4045
rect 22390 4010 22400 4030
rect 22420 4010 22430 4030
rect 22390 3980 22430 4010
rect 22390 3960 22400 3980
rect 22420 3960 22430 3980
rect 22390 3945 22430 3960
rect 22445 4030 22485 4045
rect 22445 4010 22455 4030
rect 22475 4010 22485 4030
rect 22445 3980 22485 4010
rect 22445 3960 22455 3980
rect 22475 3960 22485 3980
rect 22445 3945 22485 3960
rect 22590 4030 22630 4045
rect 22590 4010 22600 4030
rect 22620 4010 22630 4030
rect 22590 3980 22630 4010
rect 22590 3960 22600 3980
rect 22620 3960 22630 3980
rect 22590 3945 22630 3960
rect 22645 4030 22685 4045
rect 22645 4010 22655 4030
rect 22675 4010 22685 4030
rect 22645 3980 22685 4010
rect 22645 3960 22655 3980
rect 22675 3960 22685 3980
rect 22645 3945 22685 3960
rect 22755 4030 22795 4045
rect 22755 4010 22765 4030
rect 22785 4010 22795 4030
rect 22755 3980 22795 4010
rect 22755 3960 22765 3980
rect 22785 3960 22795 3980
rect 22755 3945 22795 3960
rect 22810 4030 22850 4045
rect 22810 4010 22820 4030
rect 22840 4010 22850 4030
rect 22810 3980 22850 4010
rect 22810 3960 22820 3980
rect 22840 3960 22850 3980
rect 22810 3945 22850 3960
rect 22920 4030 22960 4045
rect 22920 4010 22930 4030
rect 22950 4010 22960 4030
rect 22920 3980 22960 4010
rect 22920 3960 22930 3980
rect 22950 3960 22960 3980
rect 22920 3945 22960 3960
rect 22975 4030 23015 4045
rect 22975 4010 22985 4030
rect 23005 4010 23015 4030
rect 22975 3980 23015 4010
rect 22975 3960 22985 3980
rect 23005 3960 23015 3980
rect 22975 3945 23015 3960
rect 23190 4030 23240 4045
rect 23190 4010 23205 4030
rect 23225 4010 23240 4030
rect 23190 3980 23240 4010
rect 23190 3960 23205 3980
rect 23225 3960 23240 3980
rect 23190 3945 23240 3960
rect 23255 4030 23305 4045
rect 23255 4010 23270 4030
rect 23290 4010 23305 4030
rect 23255 3980 23305 4010
rect 23255 3960 23270 3980
rect 23290 3960 23305 3980
rect 23255 3945 23305 3960
rect 23385 4030 23435 4045
rect 23385 4010 23400 4030
rect 23420 4010 23435 4030
rect 23385 3980 23435 4010
rect 23385 3960 23400 3980
rect 23420 3960 23435 3980
rect 23385 3945 23435 3960
rect 23450 4030 23500 4045
rect 23450 4010 23465 4030
rect 23485 4010 23500 4030
rect 23450 3980 23500 4010
rect 23450 3960 23465 3980
rect 23485 3960 23500 3980
rect 23450 3945 23500 3960
rect 23580 4030 23630 4045
rect 23580 4010 23595 4030
rect 23615 4010 23630 4030
rect 23580 3980 23630 4010
rect 23580 3960 23595 3980
rect 23615 3960 23630 3980
rect 23580 3945 23630 3960
rect 23645 4030 23695 4045
rect 23645 4010 23660 4030
rect 23680 4010 23695 4030
rect 23645 3980 23695 4010
rect 23645 3960 23660 3980
rect 23680 3960 23695 3980
rect 23645 3945 23695 3960
rect 23725 4030 23775 4045
rect 23725 4010 23740 4030
rect 23760 4010 23775 4030
rect 23725 3980 23775 4010
rect 23725 3960 23740 3980
rect 23760 3960 23775 3980
rect 23725 3945 23775 3960
rect 23790 4030 23840 4045
rect 23790 4010 23805 4030
rect 23825 4010 23840 4030
rect 23790 3980 23840 4010
rect 23790 3960 23805 3980
rect 23825 3960 23840 3980
rect 23790 3945 23840 3960
rect 23920 4030 23970 4045
rect 23920 4010 23935 4030
rect 23955 4010 23970 4030
rect 23920 3980 23970 4010
rect 23920 3960 23935 3980
rect 23955 3960 23970 3980
rect 23920 3945 23970 3960
rect 23985 4030 24035 4045
rect 23985 4010 24000 4030
rect 24020 4010 24035 4030
rect 23985 3980 24035 4010
rect 23985 3960 24000 3980
rect 24020 3960 24035 3980
rect 23985 3945 24035 3960
rect 24665 4005 24715 4020
rect 24665 3985 24680 4005
rect 24700 3985 24715 4005
rect 24665 3955 24715 3985
rect 24665 3935 24680 3955
rect 24700 3935 24715 3955
rect 24665 3905 24715 3935
rect 24665 3885 24680 3905
rect 24700 3885 24715 3905
rect 24665 3855 24715 3885
rect 24665 3835 24680 3855
rect 24700 3835 24715 3855
rect 24665 3820 24715 3835
rect 24775 4005 24825 4020
rect 24775 3985 24790 4005
rect 24810 3985 24825 4005
rect 24775 3955 24825 3985
rect 24775 3935 24790 3955
rect 24810 3935 24825 3955
rect 24775 3905 24825 3935
rect 24775 3885 24790 3905
rect 24810 3885 24825 3905
rect 24775 3855 24825 3885
rect 24775 3835 24790 3855
rect 24810 3835 24825 3855
rect 24775 3820 24825 3835
rect 24885 4005 24935 4020
rect 24885 3985 24900 4005
rect 24920 3985 24935 4005
rect 24885 3955 24935 3985
rect 24885 3935 24900 3955
rect 24920 3935 24935 3955
rect 24885 3905 24935 3935
rect 24885 3885 24900 3905
rect 24920 3885 24935 3905
rect 24885 3855 24935 3885
rect 24885 3835 24900 3855
rect 24920 3835 24935 3855
rect 24885 3820 24935 3835
rect 24995 4005 25045 4020
rect 24995 3985 25010 4005
rect 25030 3985 25045 4005
rect 24995 3955 25045 3985
rect 24995 3935 25010 3955
rect 25030 3935 25045 3955
rect 24995 3905 25045 3935
rect 24995 3885 25010 3905
rect 25030 3885 25045 3905
rect 24995 3855 25045 3885
rect 24995 3835 25010 3855
rect 25030 3835 25045 3855
rect 24995 3820 25045 3835
rect 25105 4005 25155 4020
rect 25205 4005 25255 4020
rect 25105 3985 25120 4005
rect 25140 3985 25155 4005
rect 25205 3985 25220 4005
rect 25240 3985 25255 4005
rect 25105 3955 25155 3985
rect 25205 3955 25255 3985
rect 25105 3935 25120 3955
rect 25140 3935 25155 3955
rect 25205 3935 25220 3955
rect 25240 3935 25255 3955
rect 25105 3905 25155 3935
rect 25205 3905 25255 3935
rect 25105 3885 25120 3905
rect 25140 3885 25155 3905
rect 25205 3885 25220 3905
rect 25240 3885 25255 3905
rect 25105 3855 25155 3885
rect 25205 3855 25255 3885
rect 25105 3835 25120 3855
rect 25140 3835 25155 3855
rect 25205 3835 25220 3855
rect 25240 3835 25255 3855
rect 25105 3820 25155 3835
rect 25205 3820 25255 3835
rect 25315 4005 25365 4020
rect 25315 3985 25330 4005
rect 25350 3985 25365 4005
rect 25315 3955 25365 3985
rect 25315 3935 25330 3955
rect 25350 3935 25365 3955
rect 25315 3905 25365 3935
rect 25315 3885 25330 3905
rect 25350 3885 25365 3905
rect 25315 3855 25365 3885
rect 25315 3835 25330 3855
rect 25350 3835 25365 3855
rect 25315 3820 25365 3835
rect 25425 4005 25475 4020
rect 25425 3985 25440 4005
rect 25460 3985 25475 4005
rect 25425 3955 25475 3985
rect 25425 3935 25440 3955
rect 25460 3935 25475 3955
rect 25425 3905 25475 3935
rect 25425 3885 25440 3905
rect 25460 3885 25475 3905
rect 25425 3855 25475 3885
rect 25425 3835 25440 3855
rect 25460 3835 25475 3855
rect 25425 3820 25475 3835
rect 25535 4005 25585 4020
rect 25535 3985 25550 4005
rect 25570 3985 25585 4005
rect 25535 3955 25585 3985
rect 25535 3935 25550 3955
rect 25570 3935 25585 3955
rect 25535 3905 25585 3935
rect 25535 3885 25550 3905
rect 25570 3885 25585 3905
rect 25535 3855 25585 3885
rect 25535 3835 25550 3855
rect 25570 3835 25585 3855
rect 25535 3820 25585 3835
rect 25645 4005 25695 4020
rect 25745 4005 25795 4020
rect 25645 3985 25660 4005
rect 25680 3985 25695 4005
rect 25745 3985 25760 4005
rect 25780 3985 25795 4005
rect 25645 3955 25695 3985
rect 25745 3955 25795 3985
rect 25645 3935 25660 3955
rect 25680 3935 25695 3955
rect 25745 3935 25760 3955
rect 25780 3935 25795 3955
rect 25645 3905 25695 3935
rect 25745 3905 25795 3935
rect 25645 3885 25660 3905
rect 25680 3885 25695 3905
rect 25745 3885 25760 3905
rect 25780 3885 25795 3905
rect 25645 3855 25695 3885
rect 25745 3855 25795 3885
rect 25645 3835 25660 3855
rect 25680 3835 25695 3855
rect 25745 3835 25760 3855
rect 25780 3835 25795 3855
rect 25645 3820 25695 3835
rect 25745 3820 25795 3835
rect 25855 4005 25905 4020
rect 25855 3985 25870 4005
rect 25890 3985 25905 4005
rect 25855 3955 25905 3985
rect 25855 3935 25870 3955
rect 25890 3935 25905 3955
rect 25855 3905 25905 3935
rect 25855 3885 25870 3905
rect 25890 3885 25905 3905
rect 25855 3855 25905 3885
rect 25855 3835 25870 3855
rect 25890 3835 25905 3855
rect 25855 3820 25905 3835
rect 25965 4005 26015 4020
rect 25965 3985 25980 4005
rect 26000 3985 26015 4005
rect 25965 3955 26015 3985
rect 25965 3935 25980 3955
rect 26000 3935 26015 3955
rect 25965 3905 26015 3935
rect 25965 3885 25980 3905
rect 26000 3885 26015 3905
rect 25965 3855 26015 3885
rect 25965 3835 25980 3855
rect 26000 3835 26015 3855
rect 25965 3820 26015 3835
rect 26075 4005 26125 4020
rect 26075 3985 26090 4005
rect 26110 3985 26125 4005
rect 26075 3955 26125 3985
rect 26075 3935 26090 3955
rect 26110 3935 26125 3955
rect 26075 3905 26125 3935
rect 26075 3885 26090 3905
rect 26110 3885 26125 3905
rect 26075 3855 26125 3885
rect 26075 3835 26090 3855
rect 26110 3835 26125 3855
rect 26075 3820 26125 3835
rect 26185 4005 26235 4020
rect 26185 3985 26200 4005
rect 26220 3985 26235 4005
rect 26185 3955 26235 3985
rect 26185 3935 26200 3955
rect 26220 3935 26235 3955
rect 26185 3905 26235 3935
rect 26185 3885 26200 3905
rect 26220 3885 26235 3905
rect 26185 3855 26235 3885
rect 26185 3835 26200 3855
rect 26220 3835 26235 3855
rect 26185 3820 26235 3835
rect 21625 3130 21665 3145
rect 21625 3110 21635 3130
rect 21655 3110 21665 3130
rect 21625 3080 21665 3110
rect 21625 3060 21635 3080
rect 21655 3060 21665 3080
rect 21625 3045 21665 3060
rect 21680 3130 21720 3145
rect 21680 3110 21690 3130
rect 21710 3110 21720 3130
rect 21680 3080 21720 3110
rect 21680 3060 21690 3080
rect 21710 3060 21720 3080
rect 21680 3045 21720 3060
rect 21735 3130 21775 3145
rect 21735 3110 21745 3130
rect 21765 3110 21775 3130
rect 21735 3080 21775 3110
rect 21735 3060 21745 3080
rect 21765 3060 21775 3080
rect 21735 3045 21775 3060
rect 21885 3130 21925 3145
rect 21885 3110 21895 3130
rect 21915 3110 21925 3130
rect 21885 3080 21925 3110
rect 21885 3060 21895 3080
rect 21915 3060 21925 3080
rect 21885 3045 21925 3060
rect 21940 3130 21980 3145
rect 21940 3110 21950 3130
rect 21970 3110 21980 3130
rect 21940 3080 21980 3110
rect 21940 3060 21950 3080
rect 21970 3060 21980 3080
rect 21940 3045 21980 3060
rect 21995 3130 22035 3145
rect 22075 3130 22115 3145
rect 21995 3110 22005 3130
rect 22025 3110 22035 3130
rect 22075 3110 22085 3130
rect 22105 3110 22115 3130
rect 21995 3080 22035 3110
rect 22075 3080 22115 3110
rect 21995 3060 22005 3080
rect 22025 3060 22035 3080
rect 22075 3060 22085 3080
rect 22105 3060 22115 3080
rect 21995 3045 22035 3060
rect 22075 3045 22115 3060
rect 22130 3130 22170 3145
rect 22130 3110 22140 3130
rect 22160 3110 22170 3130
rect 22130 3080 22170 3110
rect 22130 3060 22140 3080
rect 22160 3060 22170 3080
rect 22130 3045 22170 3060
rect 22185 3130 22225 3145
rect 22185 3110 22195 3130
rect 22215 3110 22225 3130
rect 22185 3080 22225 3110
rect 22185 3060 22195 3080
rect 22215 3060 22225 3080
rect 22185 3045 22225 3060
rect 22335 3130 22375 3145
rect 22335 3110 22345 3130
rect 22365 3110 22375 3130
rect 22335 3080 22375 3110
rect 22335 3060 22345 3080
rect 22365 3060 22375 3080
rect 22335 3045 22375 3060
rect 22390 3130 22430 3145
rect 22390 3110 22400 3130
rect 22420 3110 22430 3130
rect 22390 3080 22430 3110
rect 22390 3060 22400 3080
rect 22420 3060 22430 3080
rect 22390 3045 22430 3060
rect 22445 3130 22485 3145
rect 22445 3110 22455 3130
rect 22475 3110 22485 3130
rect 22445 3080 22485 3110
rect 22445 3060 22455 3080
rect 22475 3060 22485 3080
rect 22445 3045 22485 3060
rect 22595 3130 22635 3145
rect 22595 3110 22605 3130
rect 22625 3110 22635 3130
rect 22595 3080 22635 3110
rect 22595 3060 22605 3080
rect 22625 3060 22635 3080
rect 22595 3045 22635 3060
rect 22650 3130 22690 3145
rect 22650 3110 22660 3130
rect 22680 3110 22690 3130
rect 22650 3080 22690 3110
rect 22650 3060 22660 3080
rect 22680 3060 22690 3080
rect 22650 3045 22690 3060
rect 22705 3130 22745 3145
rect 22705 3110 22715 3130
rect 22735 3110 22745 3130
rect 22705 3080 22745 3110
rect 22705 3060 22715 3080
rect 22735 3060 22745 3080
rect 22705 3045 22745 3060
rect 22815 3130 22855 3145
rect 22815 3110 22825 3130
rect 22845 3110 22855 3130
rect 22815 3080 22855 3110
rect 22815 3060 22825 3080
rect 22845 3060 22855 3080
rect 22815 3045 22855 3060
rect 22870 3130 22910 3145
rect 22870 3110 22880 3130
rect 22900 3110 22910 3130
rect 22870 3080 22910 3110
rect 22870 3060 22880 3080
rect 22900 3060 22910 3080
rect 22870 3045 22910 3060
rect 22980 3130 23020 3145
rect 22980 3110 22990 3130
rect 23010 3110 23020 3130
rect 22980 3080 23020 3110
rect 22980 3060 22990 3080
rect 23010 3060 23020 3080
rect 22980 3045 23020 3060
rect 23035 3130 23075 3145
rect 23035 3110 23045 3130
rect 23065 3110 23075 3130
rect 23035 3080 23075 3110
rect 23035 3060 23045 3080
rect 23065 3060 23075 3080
rect 23035 3045 23075 3060
rect 23190 3130 23240 3145
rect 23190 3110 23205 3130
rect 23225 3110 23240 3130
rect 23190 3080 23240 3110
rect 23190 3060 23205 3080
rect 23225 3060 23240 3080
rect 23190 3045 23240 3060
rect 23255 3130 23305 3145
rect 23255 3110 23270 3130
rect 23290 3110 23305 3130
rect 23255 3080 23305 3110
rect 23255 3060 23270 3080
rect 23290 3060 23305 3080
rect 23255 3045 23305 3060
rect 23385 3130 23435 3145
rect 23385 3110 23400 3130
rect 23420 3110 23435 3130
rect 23385 3080 23435 3110
rect 23385 3060 23400 3080
rect 23420 3060 23435 3080
rect 23385 3045 23435 3060
rect 23450 3130 23500 3145
rect 23450 3110 23465 3130
rect 23485 3110 23500 3130
rect 23450 3080 23500 3110
rect 23450 3060 23465 3080
rect 23485 3060 23500 3080
rect 23450 3045 23500 3060
rect 23580 3130 23630 3145
rect 23580 3110 23595 3130
rect 23615 3110 23630 3130
rect 23580 3080 23630 3110
rect 23580 3060 23595 3080
rect 23615 3060 23630 3080
rect 23580 3045 23630 3060
rect 23645 3130 23695 3145
rect 23645 3110 23660 3130
rect 23680 3110 23695 3130
rect 23645 3080 23695 3110
rect 23645 3060 23660 3080
rect 23680 3060 23695 3080
rect 23645 3045 23695 3060
rect 23725 3130 23775 3145
rect 23725 3110 23740 3130
rect 23760 3110 23775 3130
rect 23725 3080 23775 3110
rect 23725 3060 23740 3080
rect 23760 3060 23775 3080
rect 23725 3045 23775 3060
rect 23790 3130 23840 3145
rect 23790 3110 23805 3130
rect 23825 3110 23840 3130
rect 23790 3080 23840 3110
rect 23790 3060 23805 3080
rect 23825 3060 23840 3080
rect 23790 3045 23840 3060
<< pdiff >>
rect 21625 3820 21665 3835
rect 21625 3800 21635 3820
rect 21655 3800 21665 3820
rect 21625 3770 21665 3800
rect 21625 3750 21635 3770
rect 21655 3750 21665 3770
rect 21625 3720 21665 3750
rect 21625 3700 21635 3720
rect 21655 3700 21665 3720
rect 21625 3670 21665 3700
rect 21625 3650 21635 3670
rect 21655 3650 21665 3670
rect 21625 3635 21665 3650
rect 21680 3820 21720 3835
rect 21680 3800 21690 3820
rect 21710 3800 21720 3820
rect 21680 3770 21720 3800
rect 21680 3750 21690 3770
rect 21710 3750 21720 3770
rect 21680 3720 21720 3750
rect 21680 3700 21690 3720
rect 21710 3700 21720 3720
rect 21680 3670 21720 3700
rect 21680 3650 21690 3670
rect 21710 3650 21720 3670
rect 21680 3635 21720 3650
rect 21735 3820 21775 3835
rect 21735 3800 21745 3820
rect 21765 3800 21775 3820
rect 21735 3770 21775 3800
rect 21735 3750 21745 3770
rect 21765 3750 21775 3770
rect 21735 3720 21775 3750
rect 21735 3700 21745 3720
rect 21765 3700 21775 3720
rect 21735 3670 21775 3700
rect 21735 3650 21745 3670
rect 21765 3650 21775 3670
rect 21735 3635 21775 3650
rect 21885 3820 21925 3835
rect 21885 3800 21895 3820
rect 21915 3800 21925 3820
rect 21885 3770 21925 3800
rect 21885 3750 21895 3770
rect 21915 3750 21925 3770
rect 21885 3720 21925 3750
rect 21885 3700 21895 3720
rect 21915 3700 21925 3720
rect 21885 3670 21925 3700
rect 21885 3650 21895 3670
rect 21915 3650 21925 3670
rect 21885 3635 21925 3650
rect 21940 3820 21980 3835
rect 21940 3800 21950 3820
rect 21970 3800 21980 3820
rect 21940 3770 21980 3800
rect 21940 3750 21950 3770
rect 21970 3750 21980 3770
rect 21940 3720 21980 3750
rect 21940 3700 21950 3720
rect 21970 3700 21980 3720
rect 21940 3670 21980 3700
rect 21940 3650 21950 3670
rect 21970 3650 21980 3670
rect 21940 3635 21980 3650
rect 21995 3820 22035 3835
rect 22075 3820 22115 3835
rect 21995 3800 22005 3820
rect 22025 3800 22035 3820
rect 22075 3800 22085 3820
rect 22105 3800 22115 3820
rect 21995 3770 22035 3800
rect 22075 3770 22115 3800
rect 21995 3750 22005 3770
rect 22025 3750 22035 3770
rect 22075 3750 22085 3770
rect 22105 3750 22115 3770
rect 21995 3720 22035 3750
rect 22075 3720 22115 3750
rect 21995 3700 22005 3720
rect 22025 3700 22035 3720
rect 22075 3700 22085 3720
rect 22105 3700 22115 3720
rect 21995 3670 22035 3700
rect 22075 3670 22115 3700
rect 21995 3650 22005 3670
rect 22025 3650 22035 3670
rect 22075 3650 22085 3670
rect 22105 3650 22115 3670
rect 21995 3635 22035 3650
rect 22075 3635 22115 3650
rect 22130 3820 22170 3835
rect 22130 3800 22140 3820
rect 22160 3800 22170 3820
rect 22130 3770 22170 3800
rect 22130 3750 22140 3770
rect 22160 3750 22170 3770
rect 22130 3720 22170 3750
rect 22130 3700 22140 3720
rect 22160 3700 22170 3720
rect 22130 3670 22170 3700
rect 22130 3650 22140 3670
rect 22160 3650 22170 3670
rect 22130 3635 22170 3650
rect 22185 3820 22225 3835
rect 22185 3800 22195 3820
rect 22215 3800 22225 3820
rect 22185 3770 22225 3800
rect 22185 3750 22195 3770
rect 22215 3750 22225 3770
rect 22185 3720 22225 3750
rect 22185 3700 22195 3720
rect 22215 3700 22225 3720
rect 22185 3670 22225 3700
rect 22185 3650 22195 3670
rect 22215 3650 22225 3670
rect 22185 3635 22225 3650
rect 22335 3820 22375 3835
rect 22335 3800 22345 3820
rect 22365 3800 22375 3820
rect 22335 3770 22375 3800
rect 22335 3750 22345 3770
rect 22365 3750 22375 3770
rect 22335 3720 22375 3750
rect 22335 3700 22345 3720
rect 22365 3700 22375 3720
rect 22335 3670 22375 3700
rect 22335 3650 22345 3670
rect 22365 3650 22375 3670
rect 22335 3635 22375 3650
rect 22390 3820 22430 3835
rect 22390 3800 22400 3820
rect 22420 3800 22430 3820
rect 22390 3770 22430 3800
rect 22390 3750 22400 3770
rect 22420 3750 22430 3770
rect 22390 3720 22430 3750
rect 22390 3700 22400 3720
rect 22420 3700 22430 3720
rect 22390 3670 22430 3700
rect 22390 3650 22400 3670
rect 22420 3650 22430 3670
rect 22390 3635 22430 3650
rect 22445 3820 22485 3835
rect 22445 3800 22455 3820
rect 22475 3800 22485 3820
rect 22445 3770 22485 3800
rect 22445 3750 22455 3770
rect 22475 3750 22485 3770
rect 22445 3720 22485 3750
rect 22445 3700 22455 3720
rect 22475 3700 22485 3720
rect 22445 3670 22485 3700
rect 22445 3650 22455 3670
rect 22475 3650 22485 3670
rect 22445 3635 22485 3650
rect 22590 3820 22630 3835
rect 22590 3800 22600 3820
rect 22620 3800 22630 3820
rect 22590 3770 22630 3800
rect 22590 3750 22600 3770
rect 22620 3750 22630 3770
rect 22590 3720 22630 3750
rect 22590 3700 22600 3720
rect 22620 3700 22630 3720
rect 22590 3670 22630 3700
rect 22590 3650 22600 3670
rect 22620 3650 22630 3670
rect 22590 3635 22630 3650
rect 22645 3820 22685 3835
rect 22645 3800 22655 3820
rect 22675 3800 22685 3820
rect 22645 3770 22685 3800
rect 22645 3750 22655 3770
rect 22675 3750 22685 3770
rect 22645 3720 22685 3750
rect 22645 3700 22655 3720
rect 22675 3700 22685 3720
rect 22645 3670 22685 3700
rect 22645 3650 22655 3670
rect 22675 3650 22685 3670
rect 22645 3635 22685 3650
rect 22755 3820 22795 3835
rect 22755 3800 22765 3820
rect 22785 3800 22795 3820
rect 22755 3770 22795 3800
rect 22755 3750 22765 3770
rect 22785 3750 22795 3770
rect 22755 3720 22795 3750
rect 22755 3700 22765 3720
rect 22785 3700 22795 3720
rect 22755 3670 22795 3700
rect 22755 3650 22765 3670
rect 22785 3650 22795 3670
rect 22755 3635 22795 3650
rect 22810 3820 22850 3835
rect 22810 3800 22820 3820
rect 22840 3800 22850 3820
rect 22810 3770 22850 3800
rect 22810 3750 22820 3770
rect 22840 3750 22850 3770
rect 22810 3720 22850 3750
rect 22810 3700 22820 3720
rect 22840 3700 22850 3720
rect 22810 3670 22850 3700
rect 22810 3650 22820 3670
rect 22840 3650 22850 3670
rect 22810 3635 22850 3650
rect 22920 3820 22960 3835
rect 22920 3800 22930 3820
rect 22950 3800 22960 3820
rect 22920 3770 22960 3800
rect 22920 3750 22930 3770
rect 22950 3750 22960 3770
rect 22920 3720 22960 3750
rect 22920 3700 22930 3720
rect 22950 3700 22960 3720
rect 22920 3670 22960 3700
rect 22920 3650 22930 3670
rect 22950 3650 22960 3670
rect 22920 3635 22960 3650
rect 22975 3820 23015 3835
rect 22975 3800 22985 3820
rect 23005 3800 23015 3820
rect 22975 3770 23015 3800
rect 22975 3750 22985 3770
rect 23005 3750 23015 3770
rect 22975 3720 23015 3750
rect 22975 3700 22985 3720
rect 23005 3700 23015 3720
rect 22975 3670 23015 3700
rect 22975 3650 22985 3670
rect 23005 3650 23015 3670
rect 22975 3635 23015 3650
rect 23190 3820 23240 3835
rect 23190 3800 23205 3820
rect 23225 3800 23240 3820
rect 23190 3770 23240 3800
rect 23190 3750 23205 3770
rect 23225 3750 23240 3770
rect 23190 3720 23240 3750
rect 23190 3700 23205 3720
rect 23225 3700 23240 3720
rect 23190 3670 23240 3700
rect 23190 3650 23205 3670
rect 23225 3650 23240 3670
rect 23190 3635 23240 3650
rect 23255 3820 23305 3835
rect 23255 3800 23270 3820
rect 23290 3800 23305 3820
rect 23255 3770 23305 3800
rect 23255 3750 23270 3770
rect 23290 3750 23305 3770
rect 23255 3720 23305 3750
rect 23255 3700 23270 3720
rect 23290 3700 23305 3720
rect 23255 3670 23305 3700
rect 23255 3650 23270 3670
rect 23290 3650 23305 3670
rect 23255 3635 23305 3650
rect 23385 3820 23435 3835
rect 23385 3800 23400 3820
rect 23420 3800 23435 3820
rect 23385 3770 23435 3800
rect 23385 3750 23400 3770
rect 23420 3750 23435 3770
rect 23385 3720 23435 3750
rect 23385 3700 23400 3720
rect 23420 3700 23435 3720
rect 23385 3670 23435 3700
rect 23385 3650 23400 3670
rect 23420 3650 23435 3670
rect 23385 3635 23435 3650
rect 23450 3820 23500 3835
rect 23450 3800 23465 3820
rect 23485 3800 23500 3820
rect 23450 3770 23500 3800
rect 23450 3750 23465 3770
rect 23485 3750 23500 3770
rect 23450 3720 23500 3750
rect 23450 3700 23465 3720
rect 23485 3700 23500 3720
rect 23450 3670 23500 3700
rect 23450 3650 23465 3670
rect 23485 3650 23500 3670
rect 23450 3635 23500 3650
rect 23580 3820 23630 3835
rect 23580 3800 23595 3820
rect 23615 3800 23630 3820
rect 23580 3770 23630 3800
rect 23580 3750 23595 3770
rect 23615 3750 23630 3770
rect 23580 3720 23630 3750
rect 23580 3700 23595 3720
rect 23615 3700 23630 3720
rect 23580 3670 23630 3700
rect 23580 3650 23595 3670
rect 23615 3650 23630 3670
rect 23580 3635 23630 3650
rect 23645 3820 23695 3835
rect 23645 3800 23660 3820
rect 23680 3800 23695 3820
rect 23645 3770 23695 3800
rect 23645 3750 23660 3770
rect 23680 3750 23695 3770
rect 23645 3720 23695 3750
rect 23645 3700 23660 3720
rect 23680 3700 23695 3720
rect 23645 3670 23695 3700
rect 23645 3650 23660 3670
rect 23680 3650 23695 3670
rect 23645 3635 23695 3650
rect 23725 3820 23775 3835
rect 23725 3800 23740 3820
rect 23760 3800 23775 3820
rect 23725 3770 23775 3800
rect 23725 3750 23740 3770
rect 23760 3750 23775 3770
rect 23725 3720 23775 3750
rect 23725 3700 23740 3720
rect 23760 3700 23775 3720
rect 23725 3670 23775 3700
rect 23725 3650 23740 3670
rect 23760 3650 23775 3670
rect 23725 3635 23775 3650
rect 23790 3820 23840 3835
rect 23790 3800 23805 3820
rect 23825 3800 23840 3820
rect 23790 3770 23840 3800
rect 23790 3750 23805 3770
rect 23825 3750 23840 3770
rect 23790 3720 23840 3750
rect 23790 3700 23805 3720
rect 23825 3700 23840 3720
rect 23790 3670 23840 3700
rect 23790 3650 23805 3670
rect 23825 3650 23840 3670
rect 23790 3635 23840 3650
rect 24765 3455 24815 3470
rect 21625 3440 21665 3455
rect 21625 3420 21635 3440
rect 21655 3420 21665 3440
rect 21625 3390 21665 3420
rect 21625 3370 21635 3390
rect 21655 3370 21665 3390
rect 21625 3340 21665 3370
rect 21625 3320 21635 3340
rect 21655 3320 21665 3340
rect 21625 3290 21665 3320
rect 21625 3270 21635 3290
rect 21655 3270 21665 3290
rect 21625 3255 21665 3270
rect 21680 3440 21720 3455
rect 21680 3420 21690 3440
rect 21710 3420 21720 3440
rect 21680 3390 21720 3420
rect 21680 3370 21690 3390
rect 21710 3370 21720 3390
rect 21680 3340 21720 3370
rect 21680 3320 21690 3340
rect 21710 3320 21720 3340
rect 21680 3290 21720 3320
rect 21680 3270 21690 3290
rect 21710 3270 21720 3290
rect 21680 3255 21720 3270
rect 21735 3440 21775 3455
rect 21735 3420 21745 3440
rect 21765 3420 21775 3440
rect 21735 3390 21775 3420
rect 21735 3370 21745 3390
rect 21765 3370 21775 3390
rect 21735 3340 21775 3370
rect 21735 3320 21745 3340
rect 21765 3320 21775 3340
rect 21735 3290 21775 3320
rect 21735 3270 21745 3290
rect 21765 3270 21775 3290
rect 21735 3255 21775 3270
rect 21885 3440 21925 3455
rect 21885 3420 21895 3440
rect 21915 3420 21925 3440
rect 21885 3390 21925 3420
rect 21885 3370 21895 3390
rect 21915 3370 21925 3390
rect 21885 3340 21925 3370
rect 21885 3320 21895 3340
rect 21915 3320 21925 3340
rect 21885 3290 21925 3320
rect 21885 3270 21895 3290
rect 21915 3270 21925 3290
rect 21885 3255 21925 3270
rect 21940 3440 21980 3455
rect 21940 3420 21950 3440
rect 21970 3420 21980 3440
rect 21940 3390 21980 3420
rect 21940 3370 21950 3390
rect 21970 3370 21980 3390
rect 21940 3340 21980 3370
rect 21940 3320 21950 3340
rect 21970 3320 21980 3340
rect 21940 3290 21980 3320
rect 21940 3270 21950 3290
rect 21970 3270 21980 3290
rect 21940 3255 21980 3270
rect 21995 3440 22035 3455
rect 22075 3440 22115 3455
rect 21995 3420 22005 3440
rect 22025 3420 22035 3440
rect 22075 3420 22085 3440
rect 22105 3420 22115 3440
rect 21995 3390 22035 3420
rect 22075 3390 22115 3420
rect 21995 3370 22005 3390
rect 22025 3370 22035 3390
rect 22075 3370 22085 3390
rect 22105 3370 22115 3390
rect 21995 3340 22035 3370
rect 22075 3340 22115 3370
rect 21995 3320 22005 3340
rect 22025 3320 22035 3340
rect 22075 3320 22085 3340
rect 22105 3320 22115 3340
rect 21995 3290 22035 3320
rect 22075 3290 22115 3320
rect 21995 3270 22005 3290
rect 22025 3270 22035 3290
rect 22075 3270 22085 3290
rect 22105 3270 22115 3290
rect 21995 3255 22035 3270
rect 22075 3255 22115 3270
rect 22130 3440 22170 3455
rect 22130 3420 22140 3440
rect 22160 3420 22170 3440
rect 22130 3390 22170 3420
rect 22130 3370 22140 3390
rect 22160 3370 22170 3390
rect 22130 3340 22170 3370
rect 22130 3320 22140 3340
rect 22160 3320 22170 3340
rect 22130 3290 22170 3320
rect 22130 3270 22140 3290
rect 22160 3270 22170 3290
rect 22130 3255 22170 3270
rect 22185 3440 22225 3455
rect 22185 3420 22195 3440
rect 22215 3420 22225 3440
rect 22185 3390 22225 3420
rect 22185 3370 22195 3390
rect 22215 3370 22225 3390
rect 22185 3340 22225 3370
rect 22185 3320 22195 3340
rect 22215 3320 22225 3340
rect 22185 3290 22225 3320
rect 22185 3270 22195 3290
rect 22215 3270 22225 3290
rect 22185 3255 22225 3270
rect 22335 3440 22375 3455
rect 22335 3420 22345 3440
rect 22365 3420 22375 3440
rect 22335 3390 22375 3420
rect 22335 3370 22345 3390
rect 22365 3370 22375 3390
rect 22335 3340 22375 3370
rect 22335 3320 22345 3340
rect 22365 3320 22375 3340
rect 22335 3290 22375 3320
rect 22335 3270 22345 3290
rect 22365 3270 22375 3290
rect 22335 3255 22375 3270
rect 22390 3440 22430 3455
rect 22390 3420 22400 3440
rect 22420 3420 22430 3440
rect 22390 3390 22430 3420
rect 22390 3370 22400 3390
rect 22420 3370 22430 3390
rect 22390 3340 22430 3370
rect 22390 3320 22400 3340
rect 22420 3320 22430 3340
rect 22390 3290 22430 3320
rect 22390 3270 22400 3290
rect 22420 3270 22430 3290
rect 22390 3255 22430 3270
rect 22445 3440 22485 3455
rect 22445 3420 22455 3440
rect 22475 3420 22485 3440
rect 22445 3390 22485 3420
rect 22445 3370 22455 3390
rect 22475 3370 22485 3390
rect 22445 3340 22485 3370
rect 22445 3320 22455 3340
rect 22475 3320 22485 3340
rect 22445 3290 22485 3320
rect 22445 3270 22455 3290
rect 22475 3270 22485 3290
rect 22445 3255 22485 3270
rect 22595 3440 22635 3455
rect 22595 3420 22605 3440
rect 22625 3420 22635 3440
rect 22595 3390 22635 3420
rect 22595 3370 22605 3390
rect 22625 3370 22635 3390
rect 22595 3340 22635 3370
rect 22595 3320 22605 3340
rect 22625 3320 22635 3340
rect 22595 3290 22635 3320
rect 22595 3270 22605 3290
rect 22625 3270 22635 3290
rect 22595 3255 22635 3270
rect 22650 3440 22690 3455
rect 22650 3420 22660 3440
rect 22680 3420 22690 3440
rect 22650 3390 22690 3420
rect 22650 3370 22660 3390
rect 22680 3370 22690 3390
rect 22650 3340 22690 3370
rect 22650 3320 22660 3340
rect 22680 3320 22690 3340
rect 22650 3290 22690 3320
rect 22650 3270 22660 3290
rect 22680 3270 22690 3290
rect 22650 3255 22690 3270
rect 22705 3440 22745 3455
rect 22705 3420 22715 3440
rect 22735 3420 22745 3440
rect 22705 3390 22745 3420
rect 22705 3370 22715 3390
rect 22735 3370 22745 3390
rect 22705 3340 22745 3370
rect 22705 3320 22715 3340
rect 22735 3320 22745 3340
rect 22705 3290 22745 3320
rect 22705 3270 22715 3290
rect 22735 3270 22745 3290
rect 22705 3255 22745 3270
rect 22815 3440 22855 3455
rect 22815 3420 22825 3440
rect 22845 3420 22855 3440
rect 22815 3390 22855 3420
rect 22815 3370 22825 3390
rect 22845 3370 22855 3390
rect 22815 3340 22855 3370
rect 22815 3320 22825 3340
rect 22845 3320 22855 3340
rect 22815 3290 22855 3320
rect 22815 3270 22825 3290
rect 22845 3270 22855 3290
rect 22815 3255 22855 3270
rect 22870 3440 22910 3455
rect 22870 3420 22880 3440
rect 22900 3420 22910 3440
rect 22870 3390 22910 3420
rect 22870 3370 22880 3390
rect 22900 3370 22910 3390
rect 22870 3340 22910 3370
rect 22870 3320 22880 3340
rect 22900 3320 22910 3340
rect 22870 3290 22910 3320
rect 22870 3270 22880 3290
rect 22900 3270 22910 3290
rect 22870 3255 22910 3270
rect 22980 3440 23020 3455
rect 22980 3420 22990 3440
rect 23010 3420 23020 3440
rect 22980 3390 23020 3420
rect 22980 3370 22990 3390
rect 23010 3370 23020 3390
rect 22980 3340 23020 3370
rect 22980 3320 22990 3340
rect 23010 3320 23020 3340
rect 22980 3290 23020 3320
rect 22980 3270 22990 3290
rect 23010 3270 23020 3290
rect 22980 3255 23020 3270
rect 23035 3440 23075 3455
rect 23035 3420 23045 3440
rect 23065 3420 23075 3440
rect 23035 3390 23075 3420
rect 23035 3370 23045 3390
rect 23065 3370 23075 3390
rect 23035 3340 23075 3370
rect 23035 3320 23045 3340
rect 23065 3320 23075 3340
rect 23035 3290 23075 3320
rect 23035 3270 23045 3290
rect 23065 3270 23075 3290
rect 23035 3255 23075 3270
rect 23190 3440 23240 3455
rect 23190 3420 23205 3440
rect 23225 3420 23240 3440
rect 23190 3390 23240 3420
rect 23190 3370 23205 3390
rect 23225 3370 23240 3390
rect 23190 3340 23240 3370
rect 23190 3320 23205 3340
rect 23225 3320 23240 3340
rect 23190 3290 23240 3320
rect 23190 3270 23205 3290
rect 23225 3270 23240 3290
rect 23190 3255 23240 3270
rect 23255 3440 23305 3455
rect 23255 3420 23270 3440
rect 23290 3420 23305 3440
rect 23255 3390 23305 3420
rect 23255 3370 23270 3390
rect 23290 3370 23305 3390
rect 23255 3340 23305 3370
rect 23255 3320 23270 3340
rect 23290 3320 23305 3340
rect 23255 3290 23305 3320
rect 23255 3270 23270 3290
rect 23290 3270 23305 3290
rect 23255 3255 23305 3270
rect 23385 3440 23435 3455
rect 23385 3420 23400 3440
rect 23420 3420 23435 3440
rect 23385 3390 23435 3420
rect 23385 3370 23400 3390
rect 23420 3370 23435 3390
rect 23385 3340 23435 3370
rect 23385 3320 23400 3340
rect 23420 3320 23435 3340
rect 23385 3290 23435 3320
rect 23385 3270 23400 3290
rect 23420 3270 23435 3290
rect 23385 3255 23435 3270
rect 23450 3440 23500 3455
rect 23450 3420 23465 3440
rect 23485 3420 23500 3440
rect 23450 3390 23500 3420
rect 23450 3370 23465 3390
rect 23485 3370 23500 3390
rect 23450 3340 23500 3370
rect 23450 3320 23465 3340
rect 23485 3320 23500 3340
rect 23450 3290 23500 3320
rect 23450 3270 23465 3290
rect 23485 3270 23500 3290
rect 23450 3255 23500 3270
rect 23580 3440 23630 3455
rect 23580 3420 23595 3440
rect 23615 3420 23630 3440
rect 23580 3390 23630 3420
rect 23580 3370 23595 3390
rect 23615 3370 23630 3390
rect 23580 3340 23630 3370
rect 23580 3320 23595 3340
rect 23615 3320 23630 3340
rect 23580 3290 23630 3320
rect 23580 3270 23595 3290
rect 23615 3270 23630 3290
rect 23580 3255 23630 3270
rect 23645 3440 23695 3455
rect 23645 3420 23660 3440
rect 23680 3420 23695 3440
rect 23645 3390 23695 3420
rect 23645 3370 23660 3390
rect 23680 3370 23695 3390
rect 23645 3340 23695 3370
rect 23645 3320 23660 3340
rect 23680 3320 23695 3340
rect 23645 3290 23695 3320
rect 23645 3270 23660 3290
rect 23680 3270 23695 3290
rect 23645 3255 23695 3270
rect 23725 3440 23775 3455
rect 23725 3420 23740 3440
rect 23760 3420 23775 3440
rect 23725 3390 23775 3420
rect 23725 3370 23740 3390
rect 23760 3370 23775 3390
rect 23725 3340 23775 3370
rect 23725 3320 23740 3340
rect 23760 3320 23775 3340
rect 23725 3290 23775 3320
rect 23725 3270 23740 3290
rect 23760 3270 23775 3290
rect 23725 3255 23775 3270
rect 23790 3440 23840 3455
rect 23790 3420 23805 3440
rect 23825 3420 23840 3440
rect 23790 3390 23840 3420
rect 23790 3370 23805 3390
rect 23825 3370 23840 3390
rect 23790 3340 23840 3370
rect 23790 3320 23805 3340
rect 23825 3320 23840 3340
rect 23790 3290 23840 3320
rect 23790 3270 23805 3290
rect 23825 3270 23840 3290
rect 23790 3255 23840 3270
rect 23920 3440 23970 3455
rect 23920 3420 23935 3440
rect 23955 3420 23970 3440
rect 23920 3390 23970 3420
rect 23920 3370 23935 3390
rect 23955 3370 23970 3390
rect 23920 3340 23970 3370
rect 23920 3320 23935 3340
rect 23955 3320 23970 3340
rect 23920 3290 23970 3320
rect 23920 3270 23935 3290
rect 23955 3270 23970 3290
rect 23920 3255 23970 3270
rect 23985 3440 24035 3455
rect 23985 3420 24000 3440
rect 24020 3420 24035 3440
rect 23985 3390 24035 3420
rect 23985 3370 24000 3390
rect 24020 3370 24035 3390
rect 23985 3340 24035 3370
rect 23985 3320 24000 3340
rect 24020 3320 24035 3340
rect 23985 3290 24035 3320
rect 23985 3270 24000 3290
rect 24020 3270 24035 3290
rect 24765 3435 24780 3455
rect 24800 3435 24815 3455
rect 24765 3405 24815 3435
rect 24765 3385 24780 3405
rect 24800 3385 24815 3405
rect 24765 3355 24815 3385
rect 24765 3335 24780 3355
rect 24800 3335 24815 3355
rect 24765 3305 24815 3335
rect 24765 3285 24780 3305
rect 24800 3285 24815 3305
rect 24765 3270 24815 3285
rect 24875 3455 24925 3470
rect 24875 3435 24890 3455
rect 24910 3435 24925 3455
rect 24875 3405 24925 3435
rect 24875 3385 24890 3405
rect 24910 3385 24925 3405
rect 24875 3355 24925 3385
rect 24875 3335 24890 3355
rect 24910 3335 24925 3355
rect 24875 3305 24925 3335
rect 24875 3285 24890 3305
rect 24910 3285 24925 3305
rect 24875 3270 24925 3285
rect 24985 3455 25035 3470
rect 24985 3435 25000 3455
rect 25020 3435 25035 3455
rect 24985 3405 25035 3435
rect 24985 3385 25000 3405
rect 25020 3385 25035 3405
rect 24985 3355 25035 3385
rect 24985 3335 25000 3355
rect 25020 3335 25035 3355
rect 24985 3305 25035 3335
rect 24985 3285 25000 3305
rect 25020 3285 25035 3305
rect 24985 3270 25035 3285
rect 25095 3455 25145 3470
rect 25095 3435 25110 3455
rect 25130 3435 25145 3455
rect 25095 3405 25145 3435
rect 25095 3385 25110 3405
rect 25130 3385 25145 3405
rect 25095 3355 25145 3385
rect 25095 3335 25110 3355
rect 25130 3335 25145 3355
rect 25095 3305 25145 3335
rect 25095 3285 25110 3305
rect 25130 3285 25145 3305
rect 25095 3270 25145 3285
rect 25205 3455 25255 3470
rect 25205 3435 25220 3455
rect 25240 3435 25255 3455
rect 25205 3405 25255 3435
rect 25205 3385 25220 3405
rect 25240 3385 25255 3405
rect 25205 3355 25255 3385
rect 25205 3335 25220 3355
rect 25240 3335 25255 3355
rect 25205 3305 25255 3335
rect 25205 3285 25220 3305
rect 25240 3285 25255 3305
rect 25205 3270 25255 3285
rect 25315 3455 25365 3470
rect 25315 3435 25330 3455
rect 25350 3435 25365 3455
rect 25315 3405 25365 3435
rect 25315 3385 25330 3405
rect 25350 3385 25365 3405
rect 25315 3355 25365 3385
rect 25315 3335 25330 3355
rect 25350 3335 25365 3355
rect 25315 3305 25365 3335
rect 25315 3285 25330 3305
rect 25350 3285 25365 3305
rect 25315 3270 25365 3285
rect 25425 3455 25475 3470
rect 25525 3455 25575 3470
rect 25425 3435 25440 3455
rect 25460 3435 25475 3455
rect 25525 3435 25540 3455
rect 25560 3435 25575 3455
rect 25425 3405 25475 3435
rect 25525 3405 25575 3435
rect 25425 3385 25440 3405
rect 25460 3385 25475 3405
rect 25525 3385 25540 3405
rect 25560 3385 25575 3405
rect 25425 3355 25475 3385
rect 25525 3355 25575 3385
rect 25425 3335 25440 3355
rect 25460 3335 25475 3355
rect 25525 3335 25540 3355
rect 25560 3335 25575 3355
rect 25425 3305 25475 3335
rect 25525 3305 25575 3335
rect 25425 3285 25440 3305
rect 25460 3285 25475 3305
rect 25525 3285 25540 3305
rect 25560 3285 25575 3305
rect 25425 3270 25475 3285
rect 25525 3270 25575 3285
rect 25635 3455 25685 3470
rect 25635 3435 25650 3455
rect 25670 3435 25685 3455
rect 25635 3405 25685 3435
rect 25635 3385 25650 3405
rect 25670 3385 25685 3405
rect 25635 3355 25685 3385
rect 25635 3335 25650 3355
rect 25670 3335 25685 3355
rect 25635 3305 25685 3335
rect 25635 3285 25650 3305
rect 25670 3285 25685 3305
rect 25635 3270 25685 3285
rect 25745 3455 25795 3470
rect 25745 3435 25760 3455
rect 25780 3435 25795 3455
rect 25745 3405 25795 3435
rect 25745 3385 25760 3405
rect 25780 3385 25795 3405
rect 25745 3355 25795 3385
rect 25745 3335 25760 3355
rect 25780 3335 25795 3355
rect 25745 3305 25795 3335
rect 25745 3285 25760 3305
rect 25780 3285 25795 3305
rect 25745 3270 25795 3285
rect 25855 3455 25905 3470
rect 25855 3435 25870 3455
rect 25890 3435 25905 3455
rect 25855 3405 25905 3435
rect 25855 3385 25870 3405
rect 25890 3385 25905 3405
rect 25855 3355 25905 3385
rect 25855 3335 25870 3355
rect 25890 3335 25905 3355
rect 25855 3305 25905 3335
rect 25855 3285 25870 3305
rect 25890 3285 25905 3305
rect 25855 3270 25905 3285
rect 25965 3455 26015 3470
rect 25965 3435 25980 3455
rect 26000 3435 26015 3455
rect 25965 3405 26015 3435
rect 25965 3385 25980 3405
rect 26000 3385 26015 3405
rect 25965 3355 26015 3385
rect 25965 3335 25980 3355
rect 26000 3335 26015 3355
rect 25965 3305 26015 3335
rect 25965 3285 25980 3305
rect 26000 3285 26015 3305
rect 25965 3270 26015 3285
rect 26075 3455 26125 3470
rect 26075 3435 26090 3455
rect 26110 3435 26125 3455
rect 26075 3405 26125 3435
rect 26075 3385 26090 3405
rect 26110 3385 26125 3405
rect 26075 3355 26125 3385
rect 26075 3335 26090 3355
rect 26110 3335 26125 3355
rect 26075 3305 26125 3335
rect 26075 3285 26090 3305
rect 26110 3285 26125 3305
rect 26075 3270 26125 3285
rect 26185 3455 26235 3470
rect 26185 3435 26200 3455
rect 26220 3435 26235 3455
rect 26185 3405 26235 3435
rect 26185 3385 26200 3405
rect 26220 3385 26235 3405
rect 26185 3355 26235 3385
rect 26185 3335 26200 3355
rect 26220 3335 26235 3355
rect 26185 3305 26235 3335
rect 26185 3285 26200 3305
rect 26220 3285 26235 3305
rect 26185 3270 26235 3285
rect 23985 3255 24035 3270
<< ndiffc >>
rect 21635 4010 21655 4030
rect 21635 3960 21655 3980
rect 21690 4010 21710 4030
rect 21690 3960 21710 3980
rect 21745 4010 21765 4030
rect 21745 3960 21765 3980
rect 21895 4010 21915 4030
rect 21895 3960 21915 3980
rect 21950 4010 21970 4030
rect 21950 3960 21970 3980
rect 22005 4010 22025 4030
rect 22085 4010 22105 4030
rect 22005 3960 22025 3980
rect 22085 3960 22105 3980
rect 22140 4010 22160 4030
rect 22140 3960 22160 3980
rect 22195 4010 22215 4030
rect 22195 3960 22215 3980
rect 22345 4010 22365 4030
rect 22345 3960 22365 3980
rect 22400 4010 22420 4030
rect 22400 3960 22420 3980
rect 22455 4010 22475 4030
rect 22455 3960 22475 3980
rect 22600 4010 22620 4030
rect 22600 3960 22620 3980
rect 22655 4010 22675 4030
rect 22655 3960 22675 3980
rect 22765 4010 22785 4030
rect 22765 3960 22785 3980
rect 22820 4010 22840 4030
rect 22820 3960 22840 3980
rect 22930 4010 22950 4030
rect 22930 3960 22950 3980
rect 22985 4010 23005 4030
rect 22985 3960 23005 3980
rect 23205 4010 23225 4030
rect 23205 3960 23225 3980
rect 23270 4010 23290 4030
rect 23270 3960 23290 3980
rect 23400 4010 23420 4030
rect 23400 3960 23420 3980
rect 23465 4010 23485 4030
rect 23465 3960 23485 3980
rect 23595 4010 23615 4030
rect 23595 3960 23615 3980
rect 23660 4010 23680 4030
rect 23660 3960 23680 3980
rect 23740 4010 23760 4030
rect 23740 3960 23760 3980
rect 23805 4010 23825 4030
rect 23805 3960 23825 3980
rect 23935 4010 23955 4030
rect 23935 3960 23955 3980
rect 24000 4010 24020 4030
rect 24000 3960 24020 3980
rect 24680 3985 24700 4005
rect 24680 3935 24700 3955
rect 24680 3885 24700 3905
rect 24680 3835 24700 3855
rect 24790 3985 24810 4005
rect 24790 3935 24810 3955
rect 24790 3885 24810 3905
rect 24790 3835 24810 3855
rect 24900 3985 24920 4005
rect 24900 3935 24920 3955
rect 24900 3885 24920 3905
rect 24900 3835 24920 3855
rect 25010 3985 25030 4005
rect 25010 3935 25030 3955
rect 25010 3885 25030 3905
rect 25010 3835 25030 3855
rect 25120 3985 25140 4005
rect 25220 3985 25240 4005
rect 25120 3935 25140 3955
rect 25220 3935 25240 3955
rect 25120 3885 25140 3905
rect 25220 3885 25240 3905
rect 25120 3835 25140 3855
rect 25220 3835 25240 3855
rect 25330 3985 25350 4005
rect 25330 3935 25350 3955
rect 25330 3885 25350 3905
rect 25330 3835 25350 3855
rect 25440 3985 25460 4005
rect 25440 3935 25460 3955
rect 25440 3885 25460 3905
rect 25440 3835 25460 3855
rect 25550 3985 25570 4005
rect 25550 3935 25570 3955
rect 25550 3885 25570 3905
rect 25550 3835 25570 3855
rect 25660 3985 25680 4005
rect 25760 3985 25780 4005
rect 25660 3935 25680 3955
rect 25760 3935 25780 3955
rect 25660 3885 25680 3905
rect 25760 3885 25780 3905
rect 25660 3835 25680 3855
rect 25760 3835 25780 3855
rect 25870 3985 25890 4005
rect 25870 3935 25890 3955
rect 25870 3885 25890 3905
rect 25870 3835 25890 3855
rect 25980 3985 26000 4005
rect 25980 3935 26000 3955
rect 25980 3885 26000 3905
rect 25980 3835 26000 3855
rect 26090 3985 26110 4005
rect 26090 3935 26110 3955
rect 26090 3885 26110 3905
rect 26090 3835 26110 3855
rect 26200 3985 26220 4005
rect 26200 3935 26220 3955
rect 26200 3885 26220 3905
rect 26200 3835 26220 3855
rect 21635 3110 21655 3130
rect 21635 3060 21655 3080
rect 21690 3110 21710 3130
rect 21690 3060 21710 3080
rect 21745 3110 21765 3130
rect 21745 3060 21765 3080
rect 21895 3110 21915 3130
rect 21895 3060 21915 3080
rect 21950 3110 21970 3130
rect 21950 3060 21970 3080
rect 22005 3110 22025 3130
rect 22085 3110 22105 3130
rect 22005 3060 22025 3080
rect 22085 3060 22105 3080
rect 22140 3110 22160 3130
rect 22140 3060 22160 3080
rect 22195 3110 22215 3130
rect 22195 3060 22215 3080
rect 22345 3110 22365 3130
rect 22345 3060 22365 3080
rect 22400 3110 22420 3130
rect 22400 3060 22420 3080
rect 22455 3110 22475 3130
rect 22455 3060 22475 3080
rect 22605 3110 22625 3130
rect 22605 3060 22625 3080
rect 22660 3110 22680 3130
rect 22660 3060 22680 3080
rect 22715 3110 22735 3130
rect 22715 3060 22735 3080
rect 22825 3110 22845 3130
rect 22825 3060 22845 3080
rect 22880 3110 22900 3130
rect 22880 3060 22900 3080
rect 22990 3110 23010 3130
rect 22990 3060 23010 3080
rect 23045 3110 23065 3130
rect 23045 3060 23065 3080
rect 23205 3110 23225 3130
rect 23205 3060 23225 3080
rect 23270 3110 23290 3130
rect 23270 3060 23290 3080
rect 23400 3110 23420 3130
rect 23400 3060 23420 3080
rect 23465 3110 23485 3130
rect 23465 3060 23485 3080
rect 23595 3110 23615 3130
rect 23595 3060 23615 3080
rect 23660 3110 23680 3130
rect 23660 3060 23680 3080
rect 23740 3110 23760 3130
rect 23740 3060 23760 3080
rect 23805 3110 23825 3130
rect 23805 3060 23825 3080
<< pdiffc >>
rect 21635 3800 21655 3820
rect 21635 3750 21655 3770
rect 21635 3700 21655 3720
rect 21635 3650 21655 3670
rect 21690 3800 21710 3820
rect 21690 3750 21710 3770
rect 21690 3700 21710 3720
rect 21690 3650 21710 3670
rect 21745 3800 21765 3820
rect 21745 3750 21765 3770
rect 21745 3700 21765 3720
rect 21745 3650 21765 3670
rect 21895 3800 21915 3820
rect 21895 3750 21915 3770
rect 21895 3700 21915 3720
rect 21895 3650 21915 3670
rect 21950 3800 21970 3820
rect 21950 3750 21970 3770
rect 21950 3700 21970 3720
rect 21950 3650 21970 3670
rect 22005 3800 22025 3820
rect 22085 3800 22105 3820
rect 22005 3750 22025 3770
rect 22085 3750 22105 3770
rect 22005 3700 22025 3720
rect 22085 3700 22105 3720
rect 22005 3650 22025 3670
rect 22085 3650 22105 3670
rect 22140 3800 22160 3820
rect 22140 3750 22160 3770
rect 22140 3700 22160 3720
rect 22140 3650 22160 3670
rect 22195 3800 22215 3820
rect 22195 3750 22215 3770
rect 22195 3700 22215 3720
rect 22195 3650 22215 3670
rect 22345 3800 22365 3820
rect 22345 3750 22365 3770
rect 22345 3700 22365 3720
rect 22345 3650 22365 3670
rect 22400 3800 22420 3820
rect 22400 3750 22420 3770
rect 22400 3700 22420 3720
rect 22400 3650 22420 3670
rect 22455 3800 22475 3820
rect 22455 3750 22475 3770
rect 22455 3700 22475 3720
rect 22455 3650 22475 3670
rect 22600 3800 22620 3820
rect 22600 3750 22620 3770
rect 22600 3700 22620 3720
rect 22600 3650 22620 3670
rect 22655 3800 22675 3820
rect 22655 3750 22675 3770
rect 22655 3700 22675 3720
rect 22655 3650 22675 3670
rect 22765 3800 22785 3820
rect 22765 3750 22785 3770
rect 22765 3700 22785 3720
rect 22765 3650 22785 3670
rect 22820 3800 22840 3820
rect 22820 3750 22840 3770
rect 22820 3700 22840 3720
rect 22820 3650 22840 3670
rect 22930 3800 22950 3820
rect 22930 3750 22950 3770
rect 22930 3700 22950 3720
rect 22930 3650 22950 3670
rect 22985 3800 23005 3820
rect 22985 3750 23005 3770
rect 22985 3700 23005 3720
rect 22985 3650 23005 3670
rect 23205 3800 23225 3820
rect 23205 3750 23225 3770
rect 23205 3700 23225 3720
rect 23205 3650 23225 3670
rect 23270 3800 23290 3820
rect 23270 3750 23290 3770
rect 23270 3700 23290 3720
rect 23270 3650 23290 3670
rect 23400 3800 23420 3820
rect 23400 3750 23420 3770
rect 23400 3700 23420 3720
rect 23400 3650 23420 3670
rect 23465 3800 23485 3820
rect 23465 3750 23485 3770
rect 23465 3700 23485 3720
rect 23465 3650 23485 3670
rect 23595 3800 23615 3820
rect 23595 3750 23615 3770
rect 23595 3700 23615 3720
rect 23595 3650 23615 3670
rect 23660 3800 23680 3820
rect 23660 3750 23680 3770
rect 23660 3700 23680 3720
rect 23660 3650 23680 3670
rect 23740 3800 23760 3820
rect 23740 3750 23760 3770
rect 23740 3700 23760 3720
rect 23740 3650 23760 3670
rect 23805 3800 23825 3820
rect 23805 3750 23825 3770
rect 23805 3700 23825 3720
rect 23805 3650 23825 3670
rect 21635 3420 21655 3440
rect 21635 3370 21655 3390
rect 21635 3320 21655 3340
rect 21635 3270 21655 3290
rect 21690 3420 21710 3440
rect 21690 3370 21710 3390
rect 21690 3320 21710 3340
rect 21690 3270 21710 3290
rect 21745 3420 21765 3440
rect 21745 3370 21765 3390
rect 21745 3320 21765 3340
rect 21745 3270 21765 3290
rect 21895 3420 21915 3440
rect 21895 3370 21915 3390
rect 21895 3320 21915 3340
rect 21895 3270 21915 3290
rect 21950 3420 21970 3440
rect 21950 3370 21970 3390
rect 21950 3320 21970 3340
rect 21950 3270 21970 3290
rect 22005 3420 22025 3440
rect 22085 3420 22105 3440
rect 22005 3370 22025 3390
rect 22085 3370 22105 3390
rect 22005 3320 22025 3340
rect 22085 3320 22105 3340
rect 22005 3270 22025 3290
rect 22085 3270 22105 3290
rect 22140 3420 22160 3440
rect 22140 3370 22160 3390
rect 22140 3320 22160 3340
rect 22140 3270 22160 3290
rect 22195 3420 22215 3440
rect 22195 3370 22215 3390
rect 22195 3320 22215 3340
rect 22195 3270 22215 3290
rect 22345 3420 22365 3440
rect 22345 3370 22365 3390
rect 22345 3320 22365 3340
rect 22345 3270 22365 3290
rect 22400 3420 22420 3440
rect 22400 3370 22420 3390
rect 22400 3320 22420 3340
rect 22400 3270 22420 3290
rect 22455 3420 22475 3440
rect 22455 3370 22475 3390
rect 22455 3320 22475 3340
rect 22455 3270 22475 3290
rect 22605 3420 22625 3440
rect 22605 3370 22625 3390
rect 22605 3320 22625 3340
rect 22605 3270 22625 3290
rect 22660 3420 22680 3440
rect 22660 3370 22680 3390
rect 22660 3320 22680 3340
rect 22660 3270 22680 3290
rect 22715 3420 22735 3440
rect 22715 3370 22735 3390
rect 22715 3320 22735 3340
rect 22715 3270 22735 3290
rect 22825 3420 22845 3440
rect 22825 3370 22845 3390
rect 22825 3320 22845 3340
rect 22825 3270 22845 3290
rect 22880 3420 22900 3440
rect 22880 3370 22900 3390
rect 22880 3320 22900 3340
rect 22880 3270 22900 3290
rect 22990 3420 23010 3440
rect 22990 3370 23010 3390
rect 22990 3320 23010 3340
rect 22990 3270 23010 3290
rect 23045 3420 23065 3440
rect 23045 3370 23065 3390
rect 23045 3320 23065 3340
rect 23045 3270 23065 3290
rect 23205 3420 23225 3440
rect 23205 3370 23225 3390
rect 23205 3320 23225 3340
rect 23205 3270 23225 3290
rect 23270 3420 23290 3440
rect 23270 3370 23290 3390
rect 23270 3320 23290 3340
rect 23270 3270 23290 3290
rect 23400 3420 23420 3440
rect 23400 3370 23420 3390
rect 23400 3320 23420 3340
rect 23400 3270 23420 3290
rect 23465 3420 23485 3440
rect 23465 3370 23485 3390
rect 23465 3320 23485 3340
rect 23465 3270 23485 3290
rect 23595 3420 23615 3440
rect 23595 3370 23615 3390
rect 23595 3320 23615 3340
rect 23595 3270 23615 3290
rect 23660 3420 23680 3440
rect 23660 3370 23680 3390
rect 23660 3320 23680 3340
rect 23660 3270 23680 3290
rect 23740 3420 23760 3440
rect 23740 3370 23760 3390
rect 23740 3320 23760 3340
rect 23740 3270 23760 3290
rect 23805 3420 23825 3440
rect 23805 3370 23825 3390
rect 23805 3320 23825 3340
rect 23805 3270 23825 3290
rect 23935 3420 23955 3440
rect 23935 3370 23955 3390
rect 23935 3320 23955 3340
rect 23935 3270 23955 3290
rect 24000 3420 24020 3440
rect 24000 3370 24020 3390
rect 24000 3320 24020 3340
rect 24000 3270 24020 3290
rect 24780 3435 24800 3455
rect 24780 3385 24800 3405
rect 24780 3335 24800 3355
rect 24780 3285 24800 3305
rect 24890 3435 24910 3455
rect 24890 3385 24910 3405
rect 24890 3335 24910 3355
rect 24890 3285 24910 3305
rect 25000 3435 25020 3455
rect 25000 3385 25020 3405
rect 25000 3335 25020 3355
rect 25000 3285 25020 3305
rect 25110 3435 25130 3455
rect 25110 3385 25130 3405
rect 25110 3335 25130 3355
rect 25110 3285 25130 3305
rect 25220 3435 25240 3455
rect 25220 3385 25240 3405
rect 25220 3335 25240 3355
rect 25220 3285 25240 3305
rect 25330 3435 25350 3455
rect 25330 3385 25350 3405
rect 25330 3335 25350 3355
rect 25330 3285 25350 3305
rect 25440 3435 25460 3455
rect 25540 3435 25560 3455
rect 25440 3385 25460 3405
rect 25540 3385 25560 3405
rect 25440 3335 25460 3355
rect 25540 3335 25560 3355
rect 25440 3285 25460 3305
rect 25540 3285 25560 3305
rect 25650 3435 25670 3455
rect 25650 3385 25670 3405
rect 25650 3335 25670 3355
rect 25650 3285 25670 3305
rect 25760 3435 25780 3455
rect 25760 3385 25780 3405
rect 25760 3335 25780 3355
rect 25760 3285 25780 3305
rect 25870 3435 25890 3455
rect 25870 3385 25890 3405
rect 25870 3335 25890 3355
rect 25870 3285 25890 3305
rect 25980 3435 26000 3455
rect 25980 3385 26000 3405
rect 25980 3335 26000 3355
rect 25980 3285 26000 3305
rect 26090 3435 26110 3455
rect 26090 3385 26110 3405
rect 26090 3335 26110 3355
rect 26090 3285 26110 3305
rect 26200 3435 26220 3455
rect 26200 3385 26220 3405
rect 26200 3335 26220 3355
rect 26200 3285 26220 3305
<< psubdiff >>
rect 21585 4030 21625 4045
rect 21585 4010 21595 4030
rect 21615 4010 21625 4030
rect 21585 3980 21625 4010
rect 21585 3960 21595 3980
rect 21615 3960 21625 3980
rect 21585 3945 21625 3960
rect 22035 4030 22075 4045
rect 22035 4010 22045 4030
rect 22065 4010 22075 4030
rect 22035 3980 22075 4010
rect 22035 3960 22045 3980
rect 22065 3960 22075 3980
rect 22035 3945 22075 3960
rect 22485 4030 22525 4045
rect 22485 4010 22495 4030
rect 22515 4010 22525 4030
rect 22485 3980 22525 4010
rect 22485 3960 22495 3980
rect 22515 3960 22525 3980
rect 22485 3945 22525 3960
rect 22685 4030 22725 4045
rect 22685 4010 22695 4030
rect 22715 4010 22725 4030
rect 22685 3980 22725 4010
rect 22685 3960 22695 3980
rect 22715 3960 22725 3980
rect 22685 3945 22725 3960
rect 22850 4030 22890 4045
rect 22850 4010 22860 4030
rect 22880 4010 22890 4030
rect 22850 3980 22890 4010
rect 22850 3960 22860 3980
rect 22880 3960 22890 3980
rect 22850 3945 22890 3960
rect 23015 4030 23055 4045
rect 23015 4010 23025 4030
rect 23045 4010 23055 4030
rect 23015 3980 23055 4010
rect 23015 3960 23025 3980
rect 23045 3960 23055 3980
rect 23015 3945 23055 3960
rect 23140 4030 23190 4045
rect 23140 4010 23155 4030
rect 23175 4010 23190 4030
rect 23140 3980 23190 4010
rect 23140 3960 23155 3980
rect 23175 3960 23190 3980
rect 23140 3945 23190 3960
rect 23530 4030 23580 4045
rect 23530 4010 23545 4030
rect 23565 4010 23580 4030
rect 23530 3980 23580 4010
rect 23530 3960 23545 3980
rect 23565 3960 23580 3980
rect 23530 3945 23580 3960
rect 23870 4030 23920 4045
rect 23870 4010 23885 4030
rect 23905 4010 23920 4030
rect 23870 3980 23920 4010
rect 23870 3960 23885 3980
rect 23905 3960 23920 3980
rect 23870 3945 23920 3960
rect 24615 4005 24665 4020
rect 24615 3985 24630 4005
rect 24650 3985 24665 4005
rect 24615 3955 24665 3985
rect 24615 3935 24630 3955
rect 24650 3935 24665 3955
rect 24615 3905 24665 3935
rect 24615 3885 24630 3905
rect 24650 3885 24665 3905
rect 24615 3855 24665 3885
rect 24615 3835 24630 3855
rect 24650 3835 24665 3855
rect 24615 3820 24665 3835
rect 25155 4005 25205 4020
rect 25155 3985 25170 4005
rect 25190 3985 25205 4005
rect 25155 3955 25205 3985
rect 25155 3935 25170 3955
rect 25190 3935 25205 3955
rect 25155 3905 25205 3935
rect 25155 3885 25170 3905
rect 25190 3885 25205 3905
rect 25155 3855 25205 3885
rect 25155 3835 25170 3855
rect 25190 3835 25205 3855
rect 25155 3820 25205 3835
rect 25695 4005 25745 4020
rect 25695 3985 25710 4005
rect 25730 3985 25745 4005
rect 25695 3955 25745 3985
rect 25695 3935 25710 3955
rect 25730 3935 25745 3955
rect 25695 3905 25745 3935
rect 25695 3885 25710 3905
rect 25730 3885 25745 3905
rect 25695 3855 25745 3885
rect 25695 3835 25710 3855
rect 25730 3835 25745 3855
rect 25695 3820 25745 3835
rect 26235 4005 26285 4020
rect 26235 3985 26250 4005
rect 26270 3985 26285 4005
rect 26235 3955 26285 3985
rect 26235 3935 26250 3955
rect 26270 3935 26285 3955
rect 26235 3905 26285 3935
rect 26235 3885 26250 3905
rect 26270 3885 26285 3905
rect 26235 3855 26285 3885
rect 26235 3835 26250 3855
rect 26270 3835 26285 3855
rect 26235 3820 26285 3835
rect 21585 3130 21625 3145
rect 21585 3110 21595 3130
rect 21615 3110 21625 3130
rect 21585 3080 21625 3110
rect 21585 3060 21595 3080
rect 21615 3060 21625 3080
rect 21585 3045 21625 3060
rect 22035 3130 22075 3145
rect 22035 3110 22045 3130
rect 22065 3110 22075 3130
rect 22035 3080 22075 3110
rect 22035 3060 22045 3080
rect 22065 3060 22075 3080
rect 22035 3045 22075 3060
rect 22485 3130 22525 3145
rect 22485 3110 22495 3130
rect 22515 3110 22525 3130
rect 22485 3080 22525 3110
rect 22485 3060 22495 3080
rect 22515 3060 22525 3080
rect 22485 3045 22525 3060
rect 22555 3130 22595 3145
rect 22555 3110 22565 3130
rect 22585 3110 22595 3130
rect 22555 3080 22595 3110
rect 22555 3060 22565 3080
rect 22585 3060 22595 3080
rect 22555 3045 22595 3060
rect 22775 3130 22815 3145
rect 22775 3110 22785 3130
rect 22805 3110 22815 3130
rect 22775 3080 22815 3110
rect 22775 3060 22785 3080
rect 22805 3060 22815 3080
rect 22775 3045 22815 3060
rect 22940 3130 22980 3145
rect 22940 3110 22950 3130
rect 22970 3110 22980 3130
rect 22940 3080 22980 3110
rect 22940 3060 22950 3080
rect 22970 3060 22980 3080
rect 22940 3045 22980 3060
rect 23150 3130 23190 3145
rect 23150 3110 23160 3130
rect 23180 3110 23190 3130
rect 23150 3080 23190 3110
rect 23150 3060 23160 3080
rect 23180 3060 23190 3080
rect 23150 3045 23190 3060
rect 23345 3130 23385 3145
rect 23345 3110 23355 3130
rect 23375 3110 23385 3130
rect 23345 3080 23385 3110
rect 23345 3060 23355 3080
rect 23375 3060 23385 3080
rect 23345 3045 23385 3060
rect 23540 3130 23580 3145
rect 23540 3110 23550 3130
rect 23570 3110 23580 3130
rect 23540 3080 23580 3110
rect 23540 3060 23550 3080
rect 23570 3060 23580 3080
rect 23540 3045 23580 3060
<< nsubdiff >>
rect 21585 3820 21625 3835
rect 21585 3800 21595 3820
rect 21615 3800 21625 3820
rect 21585 3770 21625 3800
rect 21585 3750 21595 3770
rect 21615 3750 21625 3770
rect 21585 3720 21625 3750
rect 21585 3700 21595 3720
rect 21615 3700 21625 3720
rect 21585 3670 21625 3700
rect 21585 3650 21595 3670
rect 21615 3650 21625 3670
rect 21585 3635 21625 3650
rect 22035 3820 22075 3835
rect 22035 3800 22045 3820
rect 22065 3800 22075 3820
rect 22035 3770 22075 3800
rect 22035 3750 22045 3770
rect 22065 3750 22075 3770
rect 22035 3720 22075 3750
rect 22035 3700 22045 3720
rect 22065 3700 22075 3720
rect 22035 3670 22075 3700
rect 22035 3650 22045 3670
rect 22065 3650 22075 3670
rect 22035 3635 22075 3650
rect 22485 3820 22525 3835
rect 22485 3800 22495 3820
rect 22515 3800 22525 3820
rect 22485 3770 22525 3800
rect 22485 3750 22495 3770
rect 22515 3750 22525 3770
rect 22485 3720 22525 3750
rect 22485 3700 22495 3720
rect 22515 3700 22525 3720
rect 22485 3670 22525 3700
rect 22485 3650 22495 3670
rect 22515 3650 22525 3670
rect 22485 3635 22525 3650
rect 22685 3820 22725 3835
rect 22685 3800 22695 3820
rect 22715 3800 22725 3820
rect 22685 3770 22725 3800
rect 22685 3750 22695 3770
rect 22715 3750 22725 3770
rect 22685 3720 22725 3750
rect 22685 3700 22695 3720
rect 22715 3700 22725 3720
rect 22685 3670 22725 3700
rect 22685 3650 22695 3670
rect 22715 3650 22725 3670
rect 22685 3635 22725 3650
rect 22850 3820 22890 3835
rect 22850 3800 22860 3820
rect 22880 3800 22890 3820
rect 22850 3770 22890 3800
rect 22850 3750 22860 3770
rect 22880 3750 22890 3770
rect 22850 3720 22890 3750
rect 22850 3700 22860 3720
rect 22880 3700 22890 3720
rect 22850 3670 22890 3700
rect 22850 3650 22860 3670
rect 22880 3650 22890 3670
rect 22850 3635 22890 3650
rect 23015 3820 23055 3835
rect 23015 3800 23025 3820
rect 23045 3800 23055 3820
rect 23015 3770 23055 3800
rect 23015 3750 23025 3770
rect 23045 3750 23055 3770
rect 23015 3720 23055 3750
rect 23015 3700 23025 3720
rect 23045 3700 23055 3720
rect 23015 3670 23055 3700
rect 23015 3650 23025 3670
rect 23045 3650 23055 3670
rect 23015 3635 23055 3650
rect 23140 3820 23190 3835
rect 23140 3800 23155 3820
rect 23175 3800 23190 3820
rect 23140 3770 23190 3800
rect 23140 3750 23155 3770
rect 23175 3750 23190 3770
rect 23140 3720 23190 3750
rect 23140 3700 23155 3720
rect 23175 3700 23190 3720
rect 23140 3670 23190 3700
rect 23140 3650 23155 3670
rect 23175 3650 23190 3670
rect 23140 3635 23190 3650
rect 23530 3820 23580 3835
rect 23530 3800 23545 3820
rect 23565 3800 23580 3820
rect 23530 3770 23580 3800
rect 23530 3750 23545 3770
rect 23565 3750 23580 3770
rect 23530 3720 23580 3750
rect 23530 3700 23545 3720
rect 23565 3700 23580 3720
rect 23530 3670 23580 3700
rect 23530 3650 23545 3670
rect 23565 3650 23580 3670
rect 23530 3635 23580 3650
rect 24715 3455 24765 3470
rect 21585 3440 21625 3455
rect 21585 3420 21595 3440
rect 21615 3420 21625 3440
rect 21585 3390 21625 3420
rect 21585 3370 21595 3390
rect 21615 3370 21625 3390
rect 21585 3340 21625 3370
rect 21585 3320 21595 3340
rect 21615 3320 21625 3340
rect 21585 3290 21625 3320
rect 21585 3270 21595 3290
rect 21615 3270 21625 3290
rect 21585 3255 21625 3270
rect 22035 3440 22075 3455
rect 22035 3420 22045 3440
rect 22065 3420 22075 3440
rect 22035 3390 22075 3420
rect 22035 3370 22045 3390
rect 22065 3370 22075 3390
rect 22035 3340 22075 3370
rect 22035 3320 22045 3340
rect 22065 3320 22075 3340
rect 22035 3290 22075 3320
rect 22035 3270 22045 3290
rect 22065 3270 22075 3290
rect 22035 3255 22075 3270
rect 22485 3440 22525 3455
rect 22485 3420 22495 3440
rect 22515 3420 22525 3440
rect 22485 3390 22525 3420
rect 22485 3370 22495 3390
rect 22515 3370 22525 3390
rect 22485 3340 22525 3370
rect 22485 3320 22495 3340
rect 22515 3320 22525 3340
rect 22485 3290 22525 3320
rect 22485 3270 22495 3290
rect 22515 3270 22525 3290
rect 22485 3255 22525 3270
rect 22555 3440 22595 3455
rect 22555 3420 22565 3440
rect 22585 3420 22595 3440
rect 22555 3390 22595 3420
rect 22555 3370 22565 3390
rect 22585 3370 22595 3390
rect 22555 3340 22595 3370
rect 22555 3320 22565 3340
rect 22585 3320 22595 3340
rect 22555 3290 22595 3320
rect 22555 3270 22565 3290
rect 22585 3270 22595 3290
rect 22555 3255 22595 3270
rect 22775 3440 22815 3455
rect 22775 3420 22785 3440
rect 22805 3420 22815 3440
rect 22775 3390 22815 3420
rect 22775 3370 22785 3390
rect 22805 3370 22815 3390
rect 22775 3340 22815 3370
rect 22775 3320 22785 3340
rect 22805 3320 22815 3340
rect 22775 3290 22815 3320
rect 22775 3270 22785 3290
rect 22805 3270 22815 3290
rect 22775 3255 22815 3270
rect 22940 3440 22980 3455
rect 22940 3420 22950 3440
rect 22970 3420 22980 3440
rect 22940 3390 22980 3420
rect 22940 3370 22950 3390
rect 22970 3370 22980 3390
rect 22940 3340 22980 3370
rect 22940 3320 22950 3340
rect 22970 3320 22980 3340
rect 22940 3290 22980 3320
rect 22940 3270 22950 3290
rect 22970 3270 22980 3290
rect 22940 3255 22980 3270
rect 23140 3440 23190 3455
rect 23140 3420 23155 3440
rect 23175 3420 23190 3440
rect 23140 3390 23190 3420
rect 23140 3370 23155 3390
rect 23175 3370 23190 3390
rect 23140 3340 23190 3370
rect 23140 3320 23155 3340
rect 23175 3320 23190 3340
rect 23140 3290 23190 3320
rect 23140 3270 23155 3290
rect 23175 3270 23190 3290
rect 23140 3255 23190 3270
rect 23335 3440 23385 3455
rect 23335 3420 23350 3440
rect 23370 3420 23385 3440
rect 23335 3390 23385 3420
rect 23335 3370 23350 3390
rect 23370 3370 23385 3390
rect 23335 3340 23385 3370
rect 23335 3320 23350 3340
rect 23370 3320 23385 3340
rect 23335 3290 23385 3320
rect 23335 3270 23350 3290
rect 23370 3270 23385 3290
rect 23335 3255 23385 3270
rect 23530 3440 23580 3455
rect 23530 3420 23545 3440
rect 23565 3420 23580 3440
rect 23530 3390 23580 3420
rect 23530 3370 23545 3390
rect 23565 3370 23580 3390
rect 23530 3340 23580 3370
rect 23530 3320 23545 3340
rect 23565 3320 23580 3340
rect 23530 3290 23580 3320
rect 23530 3270 23545 3290
rect 23565 3270 23580 3290
rect 23530 3255 23580 3270
rect 23870 3440 23920 3455
rect 23870 3420 23885 3440
rect 23905 3420 23920 3440
rect 23870 3390 23920 3420
rect 23870 3370 23885 3390
rect 23905 3370 23920 3390
rect 23870 3340 23920 3370
rect 23870 3320 23885 3340
rect 23905 3320 23920 3340
rect 23870 3290 23920 3320
rect 23870 3270 23885 3290
rect 23905 3270 23920 3290
rect 23870 3255 23920 3270
rect 24715 3435 24730 3455
rect 24750 3435 24765 3455
rect 24715 3405 24765 3435
rect 24715 3385 24730 3405
rect 24750 3385 24765 3405
rect 24715 3355 24765 3385
rect 24715 3335 24730 3355
rect 24750 3335 24765 3355
rect 24715 3305 24765 3335
rect 24715 3285 24730 3305
rect 24750 3285 24765 3305
rect 24715 3270 24765 3285
rect 25475 3455 25525 3470
rect 25475 3435 25490 3455
rect 25510 3435 25525 3455
rect 25475 3405 25525 3435
rect 25475 3385 25490 3405
rect 25510 3385 25525 3405
rect 25475 3355 25525 3385
rect 25475 3335 25490 3355
rect 25510 3335 25525 3355
rect 25475 3305 25525 3335
rect 25475 3285 25490 3305
rect 25510 3285 25525 3305
rect 25475 3270 25525 3285
rect 26235 3455 26285 3470
rect 26235 3435 26250 3455
rect 26270 3435 26285 3455
rect 26235 3405 26285 3435
rect 26235 3385 26250 3405
rect 26270 3385 26285 3405
rect 26235 3355 26285 3385
rect 26235 3335 26250 3355
rect 26270 3335 26285 3355
rect 26235 3305 26285 3335
rect 26235 3285 26250 3305
rect 26270 3285 26285 3305
rect 26235 3270 26285 3285
<< psubdiffcont >>
rect 21595 4010 21615 4030
rect 21595 3960 21615 3980
rect 22045 4010 22065 4030
rect 22045 3960 22065 3980
rect 22495 4010 22515 4030
rect 22495 3960 22515 3980
rect 22695 4010 22715 4030
rect 22695 3960 22715 3980
rect 22860 4010 22880 4030
rect 22860 3960 22880 3980
rect 23025 4010 23045 4030
rect 23025 3960 23045 3980
rect 23155 4010 23175 4030
rect 23155 3960 23175 3980
rect 23545 4010 23565 4030
rect 23545 3960 23565 3980
rect 23885 4010 23905 4030
rect 23885 3960 23905 3980
rect 24630 3985 24650 4005
rect 24630 3935 24650 3955
rect 24630 3885 24650 3905
rect 24630 3835 24650 3855
rect 25170 3985 25190 4005
rect 25170 3935 25190 3955
rect 25170 3885 25190 3905
rect 25170 3835 25190 3855
rect 25710 3985 25730 4005
rect 25710 3935 25730 3955
rect 25710 3885 25730 3905
rect 25710 3835 25730 3855
rect 26250 3985 26270 4005
rect 26250 3935 26270 3955
rect 26250 3885 26270 3905
rect 26250 3835 26270 3855
rect 21595 3110 21615 3130
rect 21595 3060 21615 3080
rect 22045 3110 22065 3130
rect 22045 3060 22065 3080
rect 22495 3110 22515 3130
rect 22495 3060 22515 3080
rect 22565 3110 22585 3130
rect 22565 3060 22585 3080
rect 22785 3110 22805 3130
rect 22785 3060 22805 3080
rect 22950 3110 22970 3130
rect 22950 3060 22970 3080
rect 23160 3110 23180 3130
rect 23160 3060 23180 3080
rect 23355 3110 23375 3130
rect 23355 3060 23375 3080
rect 23550 3110 23570 3130
rect 23550 3060 23570 3080
<< nsubdiffcont >>
rect 21595 3800 21615 3820
rect 21595 3750 21615 3770
rect 21595 3700 21615 3720
rect 21595 3650 21615 3670
rect 22045 3800 22065 3820
rect 22045 3750 22065 3770
rect 22045 3700 22065 3720
rect 22045 3650 22065 3670
rect 22495 3800 22515 3820
rect 22495 3750 22515 3770
rect 22495 3700 22515 3720
rect 22495 3650 22515 3670
rect 22695 3800 22715 3820
rect 22695 3750 22715 3770
rect 22695 3700 22715 3720
rect 22695 3650 22715 3670
rect 22860 3800 22880 3820
rect 22860 3750 22880 3770
rect 22860 3700 22880 3720
rect 22860 3650 22880 3670
rect 23025 3800 23045 3820
rect 23025 3750 23045 3770
rect 23025 3700 23045 3720
rect 23025 3650 23045 3670
rect 23155 3800 23175 3820
rect 23155 3750 23175 3770
rect 23155 3700 23175 3720
rect 23155 3650 23175 3670
rect 23545 3800 23565 3820
rect 23545 3750 23565 3770
rect 23545 3700 23565 3720
rect 23545 3650 23565 3670
rect 21595 3420 21615 3440
rect 21595 3370 21615 3390
rect 21595 3320 21615 3340
rect 21595 3270 21615 3290
rect 22045 3420 22065 3440
rect 22045 3370 22065 3390
rect 22045 3320 22065 3340
rect 22045 3270 22065 3290
rect 22495 3420 22515 3440
rect 22495 3370 22515 3390
rect 22495 3320 22515 3340
rect 22495 3270 22515 3290
rect 22565 3420 22585 3440
rect 22565 3370 22585 3390
rect 22565 3320 22585 3340
rect 22565 3270 22585 3290
rect 22785 3420 22805 3440
rect 22785 3370 22805 3390
rect 22785 3320 22805 3340
rect 22785 3270 22805 3290
rect 22950 3420 22970 3440
rect 22950 3370 22970 3390
rect 22950 3320 22970 3340
rect 22950 3270 22970 3290
rect 23155 3420 23175 3440
rect 23155 3370 23175 3390
rect 23155 3320 23175 3340
rect 23155 3270 23175 3290
rect 23350 3420 23370 3440
rect 23350 3370 23370 3390
rect 23350 3320 23370 3340
rect 23350 3270 23370 3290
rect 23545 3420 23565 3440
rect 23545 3370 23565 3390
rect 23545 3320 23565 3340
rect 23545 3270 23565 3290
rect 23885 3420 23905 3440
rect 23885 3370 23905 3390
rect 23885 3320 23905 3340
rect 23885 3270 23905 3290
rect 24730 3435 24750 3455
rect 24730 3385 24750 3405
rect 24730 3335 24750 3355
rect 24730 3285 24750 3305
rect 25490 3435 25510 3455
rect 25490 3385 25510 3405
rect 25490 3335 25510 3355
rect 25490 3285 25510 3305
rect 26250 3435 26270 3455
rect 26250 3385 26270 3405
rect 26250 3335 26270 3355
rect 26250 3285 26270 3305
<< poly >>
rect 21925 4085 22130 4100
rect 21665 4045 21680 4060
rect 21720 4045 21735 4060
rect 21925 4045 21940 4085
rect 21980 4045 21995 4060
rect 22115 4045 22130 4085
rect 23435 4090 23490 4100
rect 23435 4070 23460 4090
rect 23480 4070 23490 4090
rect 23435 4060 23490 4070
rect 23765 4090 23805 4100
rect 23765 4070 23775 4090
rect 23795 4070 23805 4090
rect 23765 4060 23805 4070
rect 24670 4065 24710 4075
rect 22170 4045 22185 4060
rect 22375 4045 22390 4060
rect 22430 4045 22445 4060
rect 22630 4045 22645 4060
rect 22795 4045 22810 4060
rect 22960 4045 22975 4060
rect 23240 4045 23255 4060
rect 23435 4045 23450 4060
rect 23630 4045 23645 4060
rect 23775 4045 23790 4060
rect 23970 4045 23985 4060
rect 24670 4045 24680 4065
rect 24700 4050 24710 4065
rect 24935 4060 25425 4075
rect 24935 4050 24995 4060
rect 24700 4045 24775 4050
rect 24670 4035 24775 4045
rect 24715 4020 24775 4035
rect 24825 4030 24995 4050
rect 25365 4050 25425 4060
rect 26190 4065 26230 4075
rect 26190 4050 26200 4065
rect 24825 4020 24885 4030
rect 24935 4020 24995 4030
rect 25045 4020 25105 4035
rect 25255 4020 25315 4035
rect 25365 4030 25535 4050
rect 25365 4020 25425 4030
rect 25475 4020 25535 4030
rect 25585 4020 25645 4035
rect 25795 4020 25855 4035
rect 25905 4030 26075 4050
rect 25905 4020 25965 4030
rect 26015 4020 26075 4030
rect 26125 4045 26200 4050
rect 26220 4045 26230 4065
rect 26125 4035 26230 4045
rect 26125 4020 26185 4035
rect 21665 3910 21680 3945
rect 21565 3900 21680 3910
rect 21565 3880 21575 3900
rect 21595 3895 21680 3900
rect 21595 3880 21605 3895
rect 21565 3870 21605 3880
rect 21665 3835 21680 3895
rect 21720 3930 21735 3945
rect 21720 3920 21770 3930
rect 21925 3925 21940 3945
rect 21720 3900 21740 3920
rect 21760 3900 21770 3920
rect 21720 3890 21770 3900
rect 21815 3910 21940 3925
rect 21720 3835 21735 3890
rect 21815 3680 21830 3910
rect 21925 3835 21940 3910
rect 21980 3890 21995 3945
rect 21980 3880 22030 3890
rect 21980 3860 22000 3880
rect 22020 3860 22030 3880
rect 21980 3850 22030 3860
rect 21980 3835 21995 3850
rect 22115 3835 22130 3945
rect 22170 3930 22185 3945
rect 22170 3920 22220 3930
rect 22375 3925 22390 3945
rect 22170 3900 22190 3920
rect 22210 3900 22220 3920
rect 22170 3890 22220 3900
rect 22265 3910 22390 3925
rect 22170 3835 22185 3890
rect 21790 3670 21830 3680
rect 21790 3650 21800 3670
rect 21820 3650 21830 3670
rect 21790 3640 21830 3650
rect 22265 3680 22280 3910
rect 22375 3835 22390 3910
rect 22430 3880 22445 3945
rect 22525 3895 22605 3905
rect 22525 3880 22535 3895
rect 22430 3875 22535 3880
rect 22555 3875 22575 3895
rect 22595 3875 22605 3895
rect 22430 3865 22605 3875
rect 22630 3895 22645 3945
rect 22730 3895 22770 3905
rect 22630 3880 22740 3895
rect 22430 3835 22445 3865
rect 22630 3835 22645 3880
rect 22730 3875 22740 3880
rect 22760 3875 22770 3895
rect 22730 3865 22770 3875
rect 22795 3895 22810 3945
rect 22895 3895 22935 3905
rect 22795 3880 22905 3895
rect 22795 3835 22810 3880
rect 22895 3875 22905 3880
rect 22925 3875 22935 3895
rect 22895 3865 22935 3875
rect 22960 3895 22975 3945
rect 23240 3910 23255 3945
rect 23435 3930 23450 3945
rect 23040 3895 23080 3905
rect 22960 3880 23050 3895
rect 22960 3835 22975 3880
rect 23040 3875 23050 3880
rect 23070 3875 23080 3895
rect 23040 3865 23080 3875
rect 23115 3900 23255 3910
rect 23115 3880 23125 3900
rect 23145 3895 23255 3900
rect 23145 3880 23155 3895
rect 23115 3870 23155 3880
rect 23240 3835 23255 3895
rect 23475 3885 23515 3895
rect 23475 3865 23485 3885
rect 23505 3870 23515 3885
rect 23630 3870 23645 3945
rect 23775 3935 23790 3945
rect 23670 3925 23790 3935
rect 23670 3905 23680 3925
rect 23700 3920 23790 3925
rect 23700 3905 23710 3920
rect 23670 3900 23710 3905
rect 23970 3870 23985 3945
rect 23505 3865 23985 3870
rect 23475 3855 23985 3865
rect 23435 3835 23450 3850
rect 23630 3835 23645 3855
rect 23775 3835 23790 3855
rect 22240 3670 22280 3680
rect 22240 3650 22250 3670
rect 22270 3650 22280 3670
rect 22240 3640 22280 3650
rect 24715 3805 24775 3820
rect 24825 3810 24885 3820
rect 24935 3810 24995 3820
rect 24825 3800 24995 3810
rect 24825 3795 24900 3800
rect 24890 3780 24900 3795
rect 24920 3795 24995 3800
rect 25045 3810 25105 3820
rect 25255 3810 25315 3820
rect 25045 3795 25315 3810
rect 25365 3810 25425 3820
rect 25475 3810 25535 3820
rect 25365 3795 25535 3810
rect 25585 3810 25645 3820
rect 25795 3810 25855 3820
rect 25585 3795 25855 3810
rect 25905 3805 25965 3820
rect 26015 3805 26075 3820
rect 26125 3805 26185 3820
rect 24920 3780 24930 3795
rect 24890 3770 24930 3780
rect 25160 3775 25170 3795
rect 25190 3775 25200 3795
rect 25160 3765 25200 3775
rect 25700 3775 25710 3795
rect 25730 3775 25740 3795
rect 25700 3765 25740 3775
rect 25905 3790 26075 3805
rect 25905 3780 25945 3790
rect 25905 3760 25915 3780
rect 25935 3760 25945 3780
rect 25905 3750 25945 3760
rect 26035 3780 26075 3790
rect 26035 3760 26045 3780
rect 26065 3760 26075 3780
rect 26035 3750 26075 3760
rect 21665 3620 21680 3635
rect 21720 3620 21735 3635
rect 21925 3620 21940 3635
rect 21980 3620 21995 3635
rect 22115 3620 22130 3635
rect 22170 3620 22185 3635
rect 22375 3620 22390 3635
rect 22430 3620 22445 3635
rect 22630 3620 22645 3635
rect 22795 3620 22810 3635
rect 22960 3620 22975 3635
rect 23240 3620 23255 3635
rect 23435 3620 23450 3635
rect 23630 3620 23645 3635
rect 23775 3620 23790 3635
rect 21850 3610 21890 3620
rect 21850 3590 21860 3610
rect 21880 3590 21890 3610
rect 21850 3580 21890 3590
rect 23410 3610 23450 3620
rect 23410 3590 23420 3610
rect 23440 3590 23450 3610
rect 23410 3585 23450 3590
rect 25685 3530 25725 3540
rect 25100 3515 25140 3525
rect 22625 3500 22665 3505
rect 25100 3500 25110 3515
rect 22625 3480 22635 3500
rect 22655 3480 22665 3500
rect 24925 3495 25110 3500
rect 25130 3500 25140 3515
rect 25480 3515 25520 3525
rect 25130 3495 25315 3500
rect 25480 3495 25490 3515
rect 25510 3495 25520 3515
rect 25685 3510 25695 3530
rect 25715 3510 25725 3530
rect 25685 3500 25725 3510
rect 26035 3530 26075 3540
rect 26035 3510 26045 3530
rect 26065 3510 26075 3530
rect 26035 3500 26075 3510
rect 22625 3470 22665 3480
rect 24815 3470 24875 3485
rect 24925 3480 25315 3495
rect 24925 3470 24985 3480
rect 25035 3470 25095 3480
rect 25145 3470 25205 3480
rect 25255 3470 25315 3480
rect 25365 3480 25635 3495
rect 25365 3470 25425 3480
rect 25575 3470 25635 3480
rect 25685 3485 26075 3500
rect 25685 3470 25745 3485
rect 25795 3470 25855 3485
rect 25905 3470 25965 3485
rect 26015 3470 26075 3485
rect 26125 3470 26185 3485
rect 21665 3455 21680 3470
rect 21720 3455 21735 3470
rect 21925 3455 21940 3470
rect 21980 3455 21995 3470
rect 22115 3455 22130 3470
rect 22170 3455 22185 3470
rect 22375 3455 22390 3470
rect 22430 3455 22445 3470
rect 22635 3455 22650 3470
rect 22690 3455 22705 3470
rect 22855 3455 22870 3470
rect 23020 3455 23035 3470
rect 23240 3455 23255 3470
rect 23435 3455 23450 3470
rect 23630 3455 23645 3470
rect 23775 3455 23790 3470
rect 23970 3455 23985 3470
rect 21790 3440 21830 3450
rect 21790 3420 21800 3440
rect 21820 3420 21830 3440
rect 21790 3410 21830 3420
rect 21565 3210 21605 3220
rect 21565 3190 21575 3210
rect 21595 3195 21605 3210
rect 21665 3195 21680 3255
rect 21595 3190 21680 3195
rect 21565 3180 21680 3190
rect 21665 3145 21680 3180
rect 21720 3200 21735 3255
rect 21720 3190 21770 3200
rect 21720 3170 21740 3190
rect 21760 3170 21770 3190
rect 21720 3160 21770 3170
rect 21815 3180 21830 3410
rect 22240 3440 22280 3450
rect 22240 3420 22250 3440
rect 22270 3420 22280 3440
rect 22240 3410 22280 3420
rect 21925 3180 21940 3255
rect 21815 3165 21940 3180
rect 21720 3145 21735 3160
rect 21925 3145 21940 3165
rect 21980 3240 21995 3255
rect 21980 3230 22030 3240
rect 21980 3210 22000 3230
rect 22020 3210 22030 3230
rect 21980 3200 22030 3210
rect 21980 3145 21995 3200
rect 22115 3145 22130 3255
rect 22170 3200 22185 3255
rect 22170 3190 22220 3200
rect 22170 3170 22190 3190
rect 22210 3170 22220 3190
rect 22170 3160 22220 3170
rect 22265 3180 22280 3410
rect 24815 3255 24875 3270
rect 22375 3180 22390 3255
rect 22265 3165 22390 3180
rect 22170 3145 22185 3160
rect 22375 3145 22390 3165
rect 22430 3180 22445 3255
rect 22515 3195 22555 3205
rect 22515 3180 22525 3195
rect 22430 3175 22525 3180
rect 22545 3175 22555 3195
rect 22430 3165 22555 3175
rect 22430 3145 22445 3165
rect 22635 3145 22650 3255
rect 22690 3145 22705 3255
rect 22730 3215 22770 3225
rect 22730 3195 22740 3215
rect 22760 3210 22770 3215
rect 22855 3210 22870 3255
rect 22760 3195 22870 3210
rect 22730 3185 22770 3195
rect 22855 3145 22870 3195
rect 22895 3215 22935 3225
rect 22895 3195 22905 3215
rect 22925 3210 22935 3215
rect 23020 3210 23035 3255
rect 22925 3195 23035 3210
rect 22895 3185 22935 3195
rect 23020 3145 23035 3195
rect 23060 3215 23100 3225
rect 23060 3195 23070 3215
rect 23090 3195 23100 3215
rect 23240 3210 23255 3255
rect 23435 3225 23450 3255
rect 23060 3185 23100 3195
rect 23125 3200 23255 3210
rect 23125 3180 23135 3200
rect 23155 3195 23255 3200
rect 23155 3180 23165 3195
rect 23125 3170 23165 3180
rect 23240 3145 23255 3195
rect 23410 3215 23450 3225
rect 23410 3195 23420 3215
rect 23440 3195 23450 3215
rect 23630 3200 23645 3255
rect 23775 3240 23790 3255
rect 23670 3230 23885 3240
rect 23670 3210 23680 3230
rect 23700 3225 23855 3230
rect 23700 3210 23710 3225
rect 23670 3200 23710 3210
rect 23845 3210 23855 3225
rect 23875 3210 23885 3230
rect 23845 3200 23885 3210
rect 23410 3185 23450 3195
rect 23435 3145 23450 3185
rect 23605 3190 23645 3200
rect 23605 3170 23615 3190
rect 23635 3175 23645 3190
rect 23970 3175 23985 3255
rect 24770 3245 24875 3255
rect 24770 3225 24780 3245
rect 24800 3240 24875 3245
rect 24925 3260 24985 3270
rect 25035 3260 25095 3270
rect 25145 3260 25205 3270
rect 25255 3260 25315 3270
rect 24925 3240 25315 3260
rect 25365 3255 25425 3270
rect 25575 3255 25635 3270
rect 25685 3260 25745 3270
rect 25795 3260 25855 3270
rect 25905 3260 25965 3270
rect 26015 3260 26075 3270
rect 25685 3240 26075 3260
rect 26125 3255 26185 3270
rect 26125 3245 26230 3255
rect 26125 3240 26200 3245
rect 24800 3225 24810 3240
rect 24770 3215 24810 3225
rect 26190 3225 26200 3240
rect 26220 3225 26230 3245
rect 26190 3215 26230 3225
rect 23635 3170 23985 3175
rect 23605 3160 23985 3170
rect 23630 3145 23645 3160
rect 23775 3145 23790 3160
rect 21665 3030 21680 3045
rect 21720 3030 21735 3045
rect 21925 3005 21940 3045
rect 21980 3030 21995 3045
rect 22115 3005 22130 3045
rect 22170 3030 22185 3045
rect 22375 3030 22390 3045
rect 22430 3030 22445 3045
rect 22635 3030 22650 3045
rect 22690 3030 22705 3045
rect 22855 3030 22870 3045
rect 23020 3030 23035 3045
rect 23240 3030 23255 3045
rect 23435 3030 23450 3045
rect 23630 3030 23645 3045
rect 23775 3030 23790 3045
rect 21925 2990 22130 3005
rect 22690 3020 22730 3030
rect 22690 3000 22700 3020
rect 22720 3000 22730 3020
rect 22690 2990 22730 3000
<< polycont >>
rect 23460 4070 23480 4090
rect 23775 4070 23795 4090
rect 24680 4045 24700 4065
rect 26200 4045 26220 4065
rect 21575 3880 21595 3900
rect 21740 3900 21760 3920
rect 22000 3860 22020 3880
rect 22190 3900 22210 3920
rect 21800 3650 21820 3670
rect 22535 3875 22555 3895
rect 22575 3875 22595 3895
rect 22740 3875 22760 3895
rect 22905 3875 22925 3895
rect 23050 3875 23070 3895
rect 23125 3880 23145 3900
rect 23485 3865 23505 3885
rect 23680 3905 23700 3925
rect 22250 3650 22270 3670
rect 24900 3780 24920 3800
rect 25170 3775 25190 3795
rect 25710 3775 25730 3795
rect 25915 3760 25935 3780
rect 26045 3760 26065 3780
rect 21860 3590 21880 3610
rect 23420 3590 23440 3610
rect 22635 3480 22655 3500
rect 25110 3495 25130 3515
rect 25490 3495 25510 3515
rect 25695 3510 25715 3530
rect 26045 3510 26065 3530
rect 21800 3420 21820 3440
rect 21575 3190 21595 3210
rect 21740 3170 21760 3190
rect 22250 3420 22270 3440
rect 22000 3210 22020 3230
rect 22190 3170 22210 3190
rect 22525 3175 22545 3195
rect 22740 3195 22760 3215
rect 22905 3195 22925 3215
rect 23070 3195 23090 3215
rect 23135 3180 23155 3200
rect 23420 3195 23440 3215
rect 23680 3210 23700 3230
rect 23855 3210 23875 3230
rect 23615 3170 23635 3190
rect 24780 3225 24800 3245
rect 26200 3225 26220 3245
rect 22700 3000 22720 3020
<< locali >>
rect 26545 4190 26600 4200
rect 26545 4155 26555 4190
rect 26590 4155 26600 4190
rect 21625 4145 21665 4155
rect 21625 4125 21635 4145
rect 21655 4125 21665 4145
rect 21625 4115 21665 4125
rect 21735 4145 21775 4155
rect 21735 4125 21745 4145
rect 21765 4125 21775 4145
rect 21735 4115 21775 4125
rect 21885 4145 21925 4155
rect 21885 4125 21895 4145
rect 21915 4125 21925 4145
rect 21885 4115 21925 4125
rect 22000 4145 22040 4155
rect 22000 4125 22010 4145
rect 22030 4125 22040 4145
rect 22000 4115 22040 4125
rect 22075 4145 22115 4155
rect 22075 4125 22085 4145
rect 22105 4125 22115 4145
rect 22075 4115 22115 4125
rect 22185 4145 22225 4155
rect 22185 4125 22195 4145
rect 22215 4125 22225 4145
rect 22185 4115 22225 4125
rect 22335 4145 22375 4155
rect 22335 4125 22345 4145
rect 22365 4125 22375 4145
rect 22335 4115 22375 4125
rect 22445 4145 22485 4155
rect 22445 4125 22455 4145
rect 22475 4125 22485 4145
rect 22445 4115 22485 4125
rect 22645 4145 22685 4155
rect 22645 4125 22655 4145
rect 22675 4125 22685 4145
rect 22645 4115 22685 4125
rect 22810 4145 22850 4155
rect 22810 4125 22820 4145
rect 22840 4125 22850 4145
rect 22810 4115 22850 4125
rect 22975 4145 23015 4155
rect 22975 4125 22985 4145
rect 23005 4125 23015 4145
rect 22975 4115 23015 4125
rect 23195 4145 23235 4155
rect 23195 4125 23205 4145
rect 23225 4125 23235 4145
rect 23195 4115 23235 4125
rect 23585 4145 23625 4155
rect 23585 4125 23595 4145
rect 23615 4125 23625 4145
rect 23585 4115 23625 4125
rect 23925 4145 23965 4155
rect 26545 4145 26600 4155
rect 23925 4125 23935 4145
rect 23955 4125 23965 4145
rect 23925 4115 23965 4125
rect 21635 4040 21655 4115
rect 21745 4040 21765 4115
rect 21895 4040 21915 4115
rect 22010 4040 22030 4115
rect 22085 4040 22105 4115
rect 22195 4040 22215 4115
rect 22345 4040 22365 4115
rect 22455 4040 22475 4115
rect 22655 4040 22675 4115
rect 22820 4040 22840 4115
rect 22985 4040 23005 4115
rect 23205 4040 23225 4115
rect 23450 4090 23490 4100
rect 23450 4070 23460 4090
rect 23480 4070 23490 4090
rect 23450 4060 23490 4070
rect 23595 4040 23615 4115
rect 23765 4090 23805 4100
rect 23765 4070 23775 4090
rect 23795 4070 23805 4090
rect 23765 4060 23805 4070
rect 23935 4040 23955 4115
rect 24670 4065 24710 4075
rect 24670 4045 24680 4065
rect 24700 4045 24710 4065
rect 21590 4030 21660 4040
rect 21590 4010 21595 4030
rect 21615 4010 21635 4030
rect 21655 4010 21660 4030
rect 21590 3980 21660 4010
rect 21590 3960 21595 3980
rect 21615 3960 21635 3980
rect 21655 3960 21660 3980
rect 21590 3950 21660 3960
rect 21685 4030 21715 4040
rect 21685 4010 21690 4030
rect 21710 4010 21715 4030
rect 21685 3980 21715 4010
rect 21685 3960 21690 3980
rect 21710 3960 21715 3980
rect 21685 3950 21715 3960
rect 21740 4030 21770 4040
rect 21740 4010 21745 4030
rect 21765 4010 21770 4030
rect 21740 3980 21770 4010
rect 21740 3960 21745 3980
rect 21765 3960 21770 3980
rect 21740 3950 21770 3960
rect 21890 4030 21920 4040
rect 21890 4010 21895 4030
rect 21915 4010 21920 4030
rect 21890 3980 21920 4010
rect 21890 3960 21895 3980
rect 21915 3960 21920 3980
rect 21890 3950 21920 3960
rect 21945 4030 21975 4040
rect 21945 4010 21950 4030
rect 21970 4010 21975 4030
rect 21945 3980 21975 4010
rect 21945 3960 21950 3980
rect 21970 3960 21975 3980
rect 21945 3950 21975 3960
rect 22000 4030 22110 4040
rect 22000 4010 22005 4030
rect 22025 4010 22045 4030
rect 22065 4010 22085 4030
rect 22105 4010 22110 4030
rect 22000 3980 22110 4010
rect 22000 3960 22005 3980
rect 22025 3960 22045 3980
rect 22065 3960 22085 3980
rect 22105 3960 22110 3980
rect 22000 3950 22110 3960
rect 22135 4030 22165 4040
rect 22135 4010 22140 4030
rect 22160 4010 22165 4030
rect 22135 3980 22165 4010
rect 22135 3960 22140 3980
rect 22160 3960 22165 3980
rect 22135 3950 22165 3960
rect 22190 4030 22220 4040
rect 22190 4010 22195 4030
rect 22215 4010 22220 4030
rect 22190 3980 22220 4010
rect 22190 3960 22195 3980
rect 22215 3960 22220 3980
rect 22190 3950 22220 3960
rect 22340 4030 22370 4040
rect 22340 4010 22345 4030
rect 22365 4010 22370 4030
rect 22340 3980 22370 4010
rect 22340 3960 22345 3980
rect 22365 3960 22370 3980
rect 22340 3950 22370 3960
rect 22395 4030 22425 4040
rect 22395 4010 22400 4030
rect 22420 4010 22425 4030
rect 22395 3980 22425 4010
rect 22395 3960 22400 3980
rect 22420 3960 22425 3980
rect 22395 3950 22425 3960
rect 22450 4030 22520 4040
rect 22450 4010 22455 4030
rect 22475 4010 22495 4030
rect 22515 4010 22520 4030
rect 22450 3980 22520 4010
rect 22450 3960 22455 3980
rect 22475 3960 22495 3980
rect 22515 3960 22520 3980
rect 22450 3950 22520 3960
rect 22595 4030 22625 4040
rect 22595 4010 22600 4030
rect 22620 4010 22625 4030
rect 22595 3980 22625 4010
rect 22595 3960 22600 3980
rect 22620 3960 22625 3980
rect 22595 3950 22625 3960
rect 22650 4030 22720 4040
rect 22650 4010 22655 4030
rect 22675 4010 22695 4030
rect 22715 4010 22720 4030
rect 22650 3980 22720 4010
rect 22650 3960 22655 3980
rect 22675 3960 22695 3980
rect 22715 3960 22720 3980
rect 22650 3950 22720 3960
rect 22760 4030 22790 4040
rect 22760 4010 22765 4030
rect 22785 4010 22790 4030
rect 22760 3980 22790 4010
rect 22760 3960 22765 3980
rect 22785 3960 22790 3980
rect 22760 3950 22790 3960
rect 22815 4030 22885 4040
rect 22815 4010 22820 4030
rect 22840 4010 22860 4030
rect 22880 4010 22885 4030
rect 22815 3980 22885 4010
rect 22815 3960 22820 3980
rect 22840 3960 22860 3980
rect 22880 3960 22885 3980
rect 22815 3950 22885 3960
rect 22925 4030 22955 4040
rect 22925 4010 22930 4030
rect 22950 4010 22955 4030
rect 22925 3980 22955 4010
rect 22925 3960 22930 3980
rect 22950 3960 22955 3980
rect 22925 3950 22955 3960
rect 22980 4030 23050 4040
rect 22980 4010 22985 4030
rect 23005 4010 23025 4030
rect 23045 4010 23050 4030
rect 22980 3980 23050 4010
rect 22980 3960 22985 3980
rect 23005 3960 23025 3980
rect 23045 3960 23050 3980
rect 22980 3950 23050 3960
rect 23145 4030 23235 4040
rect 23145 4010 23155 4030
rect 23175 4010 23205 4030
rect 23225 4010 23235 4030
rect 23145 3980 23235 4010
rect 23145 3960 23155 3980
rect 23175 3960 23205 3980
rect 23225 3960 23235 3980
rect 23145 3950 23235 3960
rect 23260 4030 23300 4040
rect 23260 4010 23270 4030
rect 23290 4010 23300 4030
rect 23260 3980 23300 4010
rect 23260 3960 23270 3980
rect 23290 3960 23300 3980
rect 23260 3950 23300 3960
rect 23390 4030 23430 4040
rect 23390 4010 23400 4030
rect 23420 4010 23430 4030
rect 23390 3980 23430 4010
rect 23390 3960 23400 3980
rect 23420 3960 23430 3980
rect 23390 3950 23430 3960
rect 23455 4030 23495 4040
rect 23455 4010 23465 4030
rect 23485 4010 23495 4030
rect 23455 3980 23495 4010
rect 23455 3960 23465 3980
rect 23485 3960 23495 3980
rect 23455 3950 23495 3960
rect 23535 4030 23625 4040
rect 23535 4010 23545 4030
rect 23565 4010 23595 4030
rect 23615 4010 23625 4030
rect 23535 3980 23625 4010
rect 23535 3960 23545 3980
rect 23565 3960 23595 3980
rect 23615 3960 23625 3980
rect 23535 3950 23625 3960
rect 23650 4030 23690 4040
rect 23650 4010 23660 4030
rect 23680 4010 23690 4030
rect 23650 3980 23690 4010
rect 23650 3960 23660 3980
rect 23680 3960 23690 3980
rect 23650 3950 23690 3960
rect 23730 4030 23770 4040
rect 23730 4010 23740 4030
rect 23760 4010 23770 4030
rect 23730 3980 23770 4010
rect 23730 3960 23740 3980
rect 23760 3960 23770 3980
rect 23730 3950 23770 3960
rect 23795 4030 23835 4040
rect 23795 4010 23805 4030
rect 23825 4010 23835 4030
rect 23795 3980 23835 4010
rect 23795 3960 23805 3980
rect 23825 3960 23835 3980
rect 23795 3950 23835 3960
rect 23875 4030 23965 4040
rect 23875 4010 23885 4030
rect 23905 4010 23935 4030
rect 23955 4010 23965 4030
rect 23875 3980 23965 4010
rect 23875 3960 23885 3980
rect 23905 3960 23935 3980
rect 23955 3960 23965 3980
rect 23875 3950 23965 3960
rect 23990 4030 24030 4040
rect 24670 4035 24710 4045
rect 26190 4065 26230 4075
rect 26190 4045 26200 4065
rect 26220 4045 26230 4065
rect 26190 4035 26230 4045
rect 23990 4010 24000 4030
rect 24020 4010 24030 4030
rect 23990 3980 24030 4010
rect 23990 3960 24000 3980
rect 24020 3960 24030 3980
rect 23990 3950 24030 3960
rect 24620 4005 24710 4015
rect 24620 3985 24630 4005
rect 24650 3985 24680 4005
rect 24700 3985 24710 4005
rect 24620 3955 24710 3985
rect 21565 3900 21605 3910
rect 21565 3880 21575 3900
rect 21595 3880 21605 3900
rect 21565 3870 21605 3880
rect 21685 3870 21705 3950
rect 21730 3920 21770 3930
rect 21730 3900 21740 3920
rect 21760 3910 21770 3920
rect 21760 3900 21870 3910
rect 21730 3890 21870 3900
rect 21685 3850 21765 3870
rect 21745 3830 21765 3850
rect 21590 3820 21660 3830
rect 21590 3800 21595 3820
rect 21615 3800 21635 3820
rect 21655 3800 21660 3820
rect 21590 3770 21660 3800
rect 21590 3750 21595 3770
rect 21615 3750 21635 3770
rect 21655 3750 21660 3770
rect 21590 3720 21660 3750
rect 21590 3700 21595 3720
rect 21615 3700 21635 3720
rect 21655 3700 21660 3720
rect 21590 3670 21660 3700
rect 21590 3650 21595 3670
rect 21615 3650 21635 3670
rect 21655 3650 21660 3670
rect 21590 3640 21660 3650
rect 21685 3820 21715 3830
rect 21685 3800 21690 3820
rect 21710 3800 21715 3820
rect 21685 3770 21715 3800
rect 21685 3750 21690 3770
rect 21710 3750 21715 3770
rect 21685 3720 21715 3750
rect 21685 3700 21690 3720
rect 21710 3700 21715 3720
rect 21685 3670 21715 3700
rect 21685 3650 21690 3670
rect 21710 3650 21715 3670
rect 21685 3640 21715 3650
rect 21740 3820 21770 3830
rect 21740 3800 21745 3820
rect 21765 3800 21770 3820
rect 21740 3770 21770 3800
rect 21740 3750 21745 3770
rect 21765 3750 21770 3770
rect 21740 3720 21770 3750
rect 21740 3700 21745 3720
rect 21765 3700 21770 3720
rect 21740 3670 21770 3700
rect 21740 3650 21745 3670
rect 21765 3665 21770 3670
rect 21790 3670 21830 3680
rect 21790 3665 21800 3670
rect 21765 3650 21800 3665
rect 21820 3650 21830 3670
rect 21740 3640 21830 3650
rect 21850 3660 21870 3890
rect 21950 3870 21970 3950
rect 21895 3850 21970 3870
rect 21990 3880 22030 3890
rect 21990 3860 22000 3880
rect 22020 3870 22030 3880
rect 22135 3870 22155 3950
rect 22180 3920 22220 3930
rect 22180 3900 22190 3920
rect 22210 3910 22220 3920
rect 22210 3900 22320 3910
rect 22180 3890 22320 3900
rect 22020 3860 22215 3870
rect 21990 3850 22215 3860
rect 21895 3830 21915 3850
rect 22195 3830 22215 3850
rect 21890 3820 21920 3830
rect 21890 3800 21895 3820
rect 21915 3800 21920 3820
rect 21890 3770 21920 3800
rect 21890 3750 21895 3770
rect 21915 3750 21920 3770
rect 21890 3720 21920 3750
rect 21890 3700 21895 3720
rect 21915 3700 21920 3720
rect 21890 3670 21920 3700
rect 21890 3660 21895 3670
rect 21850 3650 21895 3660
rect 21915 3650 21920 3670
rect 21850 3640 21920 3650
rect 21945 3820 21975 3830
rect 21945 3800 21950 3820
rect 21970 3800 21975 3820
rect 21945 3770 21975 3800
rect 21945 3750 21950 3770
rect 21970 3750 21975 3770
rect 21945 3720 21975 3750
rect 21945 3700 21950 3720
rect 21970 3700 21975 3720
rect 21945 3670 21975 3700
rect 21945 3650 21950 3670
rect 21970 3650 21975 3670
rect 21945 3640 21975 3650
rect 22000 3820 22110 3830
rect 22000 3800 22005 3820
rect 22025 3800 22045 3820
rect 22065 3800 22085 3820
rect 22105 3800 22110 3820
rect 22000 3770 22110 3800
rect 22000 3750 22005 3770
rect 22025 3750 22045 3770
rect 22065 3750 22085 3770
rect 22105 3750 22110 3770
rect 22000 3720 22110 3750
rect 22000 3700 22005 3720
rect 22025 3700 22045 3720
rect 22065 3700 22085 3720
rect 22105 3700 22110 3720
rect 22000 3670 22110 3700
rect 22000 3650 22005 3670
rect 22025 3650 22045 3670
rect 22065 3650 22085 3670
rect 22105 3650 22110 3670
rect 22000 3640 22110 3650
rect 22135 3820 22165 3830
rect 22135 3800 22140 3820
rect 22160 3800 22165 3820
rect 22135 3770 22165 3800
rect 22135 3750 22140 3770
rect 22160 3750 22165 3770
rect 22135 3720 22165 3750
rect 22135 3700 22140 3720
rect 22160 3700 22165 3720
rect 22135 3670 22165 3700
rect 22135 3650 22140 3670
rect 22160 3650 22165 3670
rect 22135 3640 22165 3650
rect 22190 3820 22220 3830
rect 22190 3800 22195 3820
rect 22215 3800 22220 3820
rect 22190 3770 22220 3800
rect 22190 3750 22195 3770
rect 22215 3750 22220 3770
rect 22190 3720 22220 3750
rect 22190 3700 22195 3720
rect 22215 3700 22220 3720
rect 22190 3670 22220 3700
rect 22190 3650 22195 3670
rect 22215 3665 22220 3670
rect 22240 3670 22280 3680
rect 22240 3665 22250 3670
rect 22215 3650 22250 3665
rect 22270 3650 22280 3670
rect 22190 3640 22280 3650
rect 22300 3660 22320 3890
rect 22400 3870 22420 3950
rect 22595 3905 22615 3950
rect 22760 3905 22780 3950
rect 22925 3905 22945 3950
rect 22345 3850 22420 3870
rect 22525 3895 22615 3905
rect 22525 3875 22535 3895
rect 22555 3875 22575 3895
rect 22595 3875 22615 3895
rect 22525 3865 22615 3875
rect 22730 3895 22780 3905
rect 22730 3875 22740 3895
rect 22760 3875 22780 3895
rect 22730 3865 22780 3875
rect 22895 3895 22945 3905
rect 22895 3875 22905 3895
rect 22925 3875 22945 3895
rect 22895 3865 22945 3875
rect 23040 3895 23080 3905
rect 23040 3875 23050 3895
rect 23070 3875 23080 3895
rect 23040 3865 23080 3875
rect 23115 3900 23155 3910
rect 23115 3880 23125 3900
rect 23145 3880 23155 3900
rect 23115 3870 23155 3880
rect 23270 3870 23290 3950
rect 23400 3870 23420 3950
rect 22345 3830 22365 3850
rect 22595 3830 22615 3865
rect 22760 3830 22780 3865
rect 22925 3830 22945 3865
rect 23270 3850 23420 3870
rect 23270 3830 23290 3850
rect 23400 3830 23420 3850
rect 23465 3895 23485 3950
rect 23670 3935 23690 3950
rect 23670 3925 23710 3935
rect 23670 3905 23680 3925
rect 23700 3905 23710 3925
rect 23670 3900 23710 3905
rect 23465 3885 23515 3895
rect 23465 3865 23485 3885
rect 23505 3865 23515 3885
rect 23465 3855 23515 3865
rect 23465 3830 23485 3855
rect 23670 3830 23690 3900
rect 23740 3830 23760 3950
rect 23805 3910 23825 3950
rect 24000 3930 24020 3950
rect 24620 3935 24630 3955
rect 24650 3935 24680 3955
rect 24700 3935 24710 3955
rect 24000 3920 24040 3930
rect 24000 3910 24010 3920
rect 23805 3900 24010 3910
rect 24030 3900 24040 3920
rect 23805 3890 24040 3900
rect 24620 3905 24710 3935
rect 23805 3830 23825 3890
rect 24620 3885 24630 3905
rect 24650 3885 24680 3905
rect 24700 3885 24710 3905
rect 24620 3855 24710 3885
rect 24620 3835 24630 3855
rect 24650 3835 24680 3855
rect 24700 3835 24710 3855
rect 22340 3820 22370 3830
rect 22340 3800 22345 3820
rect 22365 3800 22370 3820
rect 22340 3770 22370 3800
rect 22340 3750 22345 3770
rect 22365 3750 22370 3770
rect 22340 3720 22370 3750
rect 22340 3700 22345 3720
rect 22365 3700 22370 3720
rect 22340 3670 22370 3700
rect 22340 3660 22345 3670
rect 22300 3650 22345 3660
rect 22365 3650 22370 3670
rect 22300 3640 22370 3650
rect 22395 3820 22425 3830
rect 22395 3800 22400 3820
rect 22420 3800 22425 3820
rect 22395 3770 22425 3800
rect 22395 3750 22400 3770
rect 22420 3750 22425 3770
rect 22395 3720 22425 3750
rect 22395 3700 22400 3720
rect 22420 3700 22425 3720
rect 22395 3670 22425 3700
rect 22395 3650 22400 3670
rect 22420 3650 22425 3670
rect 22395 3640 22425 3650
rect 22450 3820 22520 3830
rect 22450 3800 22455 3820
rect 22475 3800 22495 3820
rect 22515 3800 22520 3820
rect 22450 3770 22520 3800
rect 22450 3750 22455 3770
rect 22475 3750 22495 3770
rect 22515 3750 22520 3770
rect 22450 3720 22520 3750
rect 22450 3700 22455 3720
rect 22475 3700 22495 3720
rect 22515 3700 22520 3720
rect 22450 3670 22520 3700
rect 22450 3650 22455 3670
rect 22475 3650 22495 3670
rect 22515 3650 22520 3670
rect 22450 3640 22520 3650
rect 22595 3820 22625 3830
rect 22595 3800 22600 3820
rect 22620 3800 22625 3820
rect 22595 3770 22625 3800
rect 22595 3750 22600 3770
rect 22620 3750 22625 3770
rect 22595 3720 22625 3750
rect 22595 3700 22600 3720
rect 22620 3700 22625 3720
rect 22595 3670 22625 3700
rect 22595 3650 22600 3670
rect 22620 3650 22625 3670
rect 22595 3640 22625 3650
rect 22650 3820 22720 3830
rect 22650 3800 22655 3820
rect 22675 3800 22695 3820
rect 22715 3800 22720 3820
rect 22650 3770 22720 3800
rect 22650 3750 22655 3770
rect 22675 3750 22695 3770
rect 22715 3750 22720 3770
rect 22650 3720 22720 3750
rect 22650 3700 22655 3720
rect 22675 3700 22695 3720
rect 22715 3700 22720 3720
rect 22650 3670 22720 3700
rect 22650 3650 22655 3670
rect 22675 3650 22695 3670
rect 22715 3650 22720 3670
rect 22650 3640 22720 3650
rect 22760 3820 22790 3830
rect 22760 3800 22765 3820
rect 22785 3800 22790 3820
rect 22760 3770 22790 3800
rect 22760 3750 22765 3770
rect 22785 3750 22790 3770
rect 22760 3720 22790 3750
rect 22760 3700 22765 3720
rect 22785 3700 22790 3720
rect 22760 3670 22790 3700
rect 22760 3650 22765 3670
rect 22785 3650 22790 3670
rect 22760 3640 22790 3650
rect 22815 3820 22885 3830
rect 22815 3800 22820 3820
rect 22840 3800 22860 3820
rect 22880 3800 22885 3820
rect 22815 3770 22885 3800
rect 22815 3750 22820 3770
rect 22840 3750 22860 3770
rect 22880 3750 22885 3770
rect 22815 3720 22885 3750
rect 22815 3700 22820 3720
rect 22840 3700 22860 3720
rect 22880 3700 22885 3720
rect 22815 3670 22885 3700
rect 22815 3650 22820 3670
rect 22840 3650 22860 3670
rect 22880 3650 22885 3670
rect 22815 3640 22885 3650
rect 22925 3820 22955 3830
rect 22925 3800 22930 3820
rect 22950 3800 22955 3820
rect 22925 3770 22955 3800
rect 22925 3750 22930 3770
rect 22950 3750 22955 3770
rect 22925 3720 22955 3750
rect 22925 3700 22930 3720
rect 22950 3700 22955 3720
rect 22925 3670 22955 3700
rect 22925 3650 22930 3670
rect 22950 3650 22955 3670
rect 22925 3640 22955 3650
rect 22980 3820 23050 3830
rect 22980 3800 22985 3820
rect 23005 3800 23025 3820
rect 23045 3800 23050 3820
rect 22980 3770 23050 3800
rect 22980 3750 22985 3770
rect 23005 3750 23025 3770
rect 23045 3750 23050 3770
rect 22980 3720 23050 3750
rect 22980 3700 22985 3720
rect 23005 3700 23025 3720
rect 23045 3700 23050 3720
rect 22980 3670 23050 3700
rect 22980 3650 22985 3670
rect 23005 3650 23025 3670
rect 23045 3650 23050 3670
rect 22980 3640 23050 3650
rect 23145 3820 23235 3830
rect 23145 3800 23155 3820
rect 23175 3800 23205 3820
rect 23225 3800 23235 3820
rect 23145 3770 23235 3800
rect 23145 3750 23155 3770
rect 23175 3750 23205 3770
rect 23225 3750 23235 3770
rect 23145 3720 23235 3750
rect 23145 3700 23155 3720
rect 23175 3700 23205 3720
rect 23225 3700 23235 3720
rect 23145 3670 23235 3700
rect 23145 3650 23155 3670
rect 23175 3650 23205 3670
rect 23225 3650 23235 3670
rect 23145 3640 23235 3650
rect 23260 3820 23300 3830
rect 23260 3800 23270 3820
rect 23290 3800 23300 3820
rect 23260 3770 23300 3800
rect 23260 3750 23270 3770
rect 23290 3750 23300 3770
rect 23260 3720 23300 3750
rect 23260 3700 23270 3720
rect 23290 3700 23300 3720
rect 23260 3670 23300 3700
rect 23260 3650 23270 3670
rect 23290 3650 23300 3670
rect 23260 3640 23300 3650
rect 23390 3820 23430 3830
rect 23390 3800 23400 3820
rect 23420 3800 23430 3820
rect 23390 3770 23430 3800
rect 23390 3750 23400 3770
rect 23420 3750 23430 3770
rect 23390 3720 23430 3750
rect 23390 3700 23400 3720
rect 23420 3700 23430 3720
rect 23390 3670 23430 3700
rect 23390 3650 23400 3670
rect 23420 3650 23430 3670
rect 23390 3640 23430 3650
rect 23455 3820 23495 3830
rect 23455 3800 23465 3820
rect 23485 3800 23495 3820
rect 23455 3770 23495 3800
rect 23455 3750 23465 3770
rect 23485 3750 23495 3770
rect 23455 3720 23495 3750
rect 23455 3700 23465 3720
rect 23485 3700 23495 3720
rect 23455 3670 23495 3700
rect 23455 3650 23465 3670
rect 23485 3650 23495 3670
rect 23455 3640 23495 3650
rect 23535 3820 23625 3830
rect 23535 3800 23545 3820
rect 23565 3800 23595 3820
rect 23615 3800 23625 3820
rect 23535 3770 23625 3800
rect 23535 3750 23545 3770
rect 23565 3750 23595 3770
rect 23615 3750 23625 3770
rect 23535 3720 23625 3750
rect 23535 3700 23545 3720
rect 23565 3700 23595 3720
rect 23615 3700 23625 3720
rect 23535 3670 23625 3700
rect 23535 3650 23545 3670
rect 23565 3650 23595 3670
rect 23615 3650 23625 3670
rect 23535 3640 23625 3650
rect 23650 3820 23690 3830
rect 23650 3800 23660 3820
rect 23680 3800 23690 3820
rect 23650 3770 23690 3800
rect 23650 3750 23660 3770
rect 23680 3750 23690 3770
rect 23650 3720 23690 3750
rect 23650 3700 23660 3720
rect 23680 3700 23690 3720
rect 23650 3670 23690 3700
rect 23650 3650 23660 3670
rect 23680 3650 23690 3670
rect 23650 3640 23690 3650
rect 23730 3820 23770 3830
rect 23730 3800 23740 3820
rect 23760 3800 23770 3820
rect 23730 3770 23770 3800
rect 23730 3750 23740 3770
rect 23760 3750 23770 3770
rect 23730 3720 23770 3750
rect 23730 3700 23740 3720
rect 23760 3700 23770 3720
rect 23730 3670 23770 3700
rect 23730 3650 23740 3670
rect 23760 3650 23770 3670
rect 23730 3640 23770 3650
rect 23795 3820 23835 3830
rect 24620 3825 24710 3835
rect 24780 4005 24820 4015
rect 24780 3985 24790 4005
rect 24810 3985 24820 4005
rect 24780 3955 24820 3985
rect 24780 3935 24790 3955
rect 24810 3935 24820 3955
rect 24780 3905 24820 3935
rect 24780 3885 24790 3905
rect 24810 3885 24820 3905
rect 24780 3855 24820 3885
rect 24780 3835 24790 3855
rect 24810 3835 24820 3855
rect 24780 3825 24820 3835
rect 24890 4005 24930 4015
rect 24890 3985 24900 4005
rect 24920 3985 24930 4005
rect 24890 3955 24930 3985
rect 24890 3935 24900 3955
rect 24920 3935 24930 3955
rect 24890 3905 24930 3935
rect 24890 3885 24900 3905
rect 24920 3885 24930 3905
rect 24890 3855 24930 3885
rect 24890 3835 24900 3855
rect 24920 3835 24930 3855
rect 23795 3800 23805 3820
rect 23825 3800 23835 3820
rect 23795 3770 23835 3800
rect 24890 3800 24930 3835
rect 25000 4005 25040 4015
rect 25000 3985 25010 4005
rect 25030 3985 25040 4005
rect 25000 3955 25040 3985
rect 25000 3935 25010 3955
rect 25030 3935 25040 3955
rect 25000 3905 25040 3935
rect 25000 3885 25010 3905
rect 25030 3885 25040 3905
rect 25000 3855 25040 3885
rect 25000 3835 25010 3855
rect 25030 3835 25040 3855
rect 25000 3825 25040 3835
rect 25110 4005 25250 4015
rect 25110 3985 25120 4005
rect 25140 3985 25170 4005
rect 25190 3985 25220 4005
rect 25240 3985 25250 4005
rect 25110 3955 25250 3985
rect 25110 3935 25120 3955
rect 25140 3935 25170 3955
rect 25190 3935 25220 3955
rect 25240 3935 25250 3955
rect 25110 3905 25250 3935
rect 25110 3885 25120 3905
rect 25140 3885 25170 3905
rect 25190 3885 25220 3905
rect 25240 3885 25250 3905
rect 25110 3855 25250 3885
rect 25110 3835 25120 3855
rect 25140 3835 25170 3855
rect 25190 3835 25220 3855
rect 25240 3835 25250 3855
rect 25110 3825 25250 3835
rect 25320 4005 25360 4015
rect 25320 3985 25330 4005
rect 25350 3985 25360 4005
rect 25320 3955 25360 3985
rect 25320 3935 25330 3955
rect 25350 3935 25360 3955
rect 25320 3905 25360 3935
rect 25320 3885 25330 3905
rect 25350 3885 25360 3905
rect 25320 3855 25360 3885
rect 25320 3835 25330 3855
rect 25350 3835 25360 3855
rect 25320 3825 25360 3835
rect 25430 4005 25470 4015
rect 25430 3985 25440 4005
rect 25460 3985 25470 4005
rect 25430 3955 25470 3985
rect 25430 3935 25440 3955
rect 25460 3935 25470 3955
rect 25430 3905 25470 3935
rect 25430 3885 25440 3905
rect 25460 3885 25470 3905
rect 25430 3855 25470 3885
rect 25430 3835 25440 3855
rect 25460 3835 25470 3855
rect 25430 3825 25470 3835
rect 25540 4005 25580 4015
rect 25540 3985 25550 4005
rect 25570 3985 25580 4005
rect 25540 3955 25580 3985
rect 25540 3935 25550 3955
rect 25570 3935 25580 3955
rect 25540 3905 25580 3935
rect 25540 3885 25550 3905
rect 25570 3885 25580 3905
rect 25540 3855 25580 3885
rect 25540 3835 25550 3855
rect 25570 3835 25580 3855
rect 25540 3825 25580 3835
rect 25650 4005 25790 4015
rect 25650 3985 25660 4005
rect 25680 3985 25710 4005
rect 25730 3985 25760 4005
rect 25780 3985 25790 4005
rect 25650 3955 25790 3985
rect 25650 3935 25660 3955
rect 25680 3935 25710 3955
rect 25730 3935 25760 3955
rect 25780 3935 25790 3955
rect 25650 3905 25790 3935
rect 25650 3885 25660 3905
rect 25680 3885 25710 3905
rect 25730 3885 25760 3905
rect 25780 3885 25790 3905
rect 25650 3855 25790 3885
rect 25650 3835 25660 3855
rect 25680 3835 25710 3855
rect 25730 3835 25760 3855
rect 25780 3835 25790 3855
rect 25650 3825 25790 3835
rect 25860 4005 25900 4015
rect 25860 3985 25870 4005
rect 25890 3985 25900 4005
rect 25860 3955 25900 3985
rect 25860 3935 25870 3955
rect 25890 3935 25900 3955
rect 25860 3905 25900 3935
rect 25860 3885 25870 3905
rect 25890 3885 25900 3905
rect 25860 3855 25900 3885
rect 25860 3835 25870 3855
rect 25890 3835 25900 3855
rect 25860 3825 25900 3835
rect 25970 4005 26010 4015
rect 25970 3985 25980 4005
rect 26000 3985 26010 4005
rect 25970 3955 26010 3985
rect 25970 3935 25980 3955
rect 26000 3935 26010 3955
rect 25970 3905 26010 3935
rect 25970 3885 25980 3905
rect 26000 3885 26010 3905
rect 25970 3855 26010 3885
rect 25970 3835 25980 3855
rect 26000 3835 26010 3855
rect 25970 3825 26010 3835
rect 26080 4005 26120 4015
rect 26080 3985 26090 4005
rect 26110 3985 26120 4005
rect 26080 3955 26120 3985
rect 26080 3935 26090 3955
rect 26110 3935 26120 3955
rect 26080 3905 26120 3935
rect 26080 3885 26090 3905
rect 26110 3885 26120 3905
rect 26080 3855 26120 3885
rect 26080 3835 26090 3855
rect 26110 3835 26120 3855
rect 26080 3825 26120 3835
rect 26190 4005 26280 4015
rect 26190 3985 26200 4005
rect 26220 3985 26250 4005
rect 26270 3985 26280 4005
rect 26190 3955 26280 3985
rect 26190 3935 26200 3955
rect 26220 3935 26250 3955
rect 26270 3935 26280 3955
rect 26190 3905 26280 3935
rect 26190 3885 26200 3905
rect 26220 3885 26250 3905
rect 26270 3885 26280 3905
rect 26190 3855 26280 3885
rect 26190 3835 26200 3855
rect 26220 3835 26250 3855
rect 26270 3835 26280 3855
rect 26190 3825 26280 3835
rect 24890 3780 24900 3800
rect 24920 3780 24930 3800
rect 24890 3770 24930 3780
rect 25160 3795 25200 3825
rect 25160 3775 25170 3795
rect 25190 3775 25200 3795
rect 23795 3750 23805 3770
rect 23825 3750 23835 3770
rect 25160 3765 25200 3775
rect 25700 3795 25740 3825
rect 25700 3775 25710 3795
rect 25730 3775 25740 3795
rect 26370 3795 26425 3805
rect 25700 3765 25740 3775
rect 25905 3780 25945 3790
rect 25905 3760 25915 3780
rect 25935 3760 25945 3780
rect 25905 3750 25945 3760
rect 26035 3780 26075 3790
rect 26035 3760 26045 3780
rect 26065 3760 26075 3780
rect 26035 3750 26075 3760
rect 26370 3760 26380 3795
rect 26415 3760 26425 3795
rect 26370 3750 26425 3760
rect 23795 3720 23835 3750
rect 23795 3700 23805 3720
rect 23825 3700 23835 3720
rect 23795 3670 23835 3700
rect 23795 3650 23805 3670
rect 23825 3650 23835 3670
rect 23795 3640 23835 3650
rect 21635 3565 21655 3640
rect 21850 3620 21870 3640
rect 21850 3610 21890 3620
rect 21850 3590 21860 3610
rect 21880 3590 21890 3610
rect 21850 3580 21890 3590
rect 22005 3565 22025 3640
rect 22085 3565 22105 3640
rect 22455 3565 22475 3640
rect 22665 3565 22685 3640
rect 22820 3565 22840 3640
rect 22985 3565 23005 3640
rect 23205 3565 23225 3640
rect 23410 3610 23450 3620
rect 23410 3590 23420 3610
rect 23440 3590 23450 3610
rect 23410 3585 23450 3590
rect 23595 3565 23615 3640
rect 23740 3620 23760 3640
rect 23730 3610 23770 3620
rect 23730 3590 23740 3610
rect 23760 3590 23770 3610
rect 23730 3580 23770 3590
rect 21625 3555 21665 3565
rect 21625 3535 21635 3555
rect 21655 3535 21665 3555
rect 21625 3525 21665 3535
rect 21995 3555 22035 3565
rect 21995 3535 22005 3555
rect 22025 3535 22035 3555
rect 21995 3525 22035 3535
rect 22075 3555 22115 3565
rect 22075 3535 22085 3555
rect 22105 3535 22115 3555
rect 22075 3525 22115 3535
rect 22445 3555 22485 3565
rect 22445 3535 22455 3555
rect 22475 3535 22485 3555
rect 22445 3525 22485 3535
rect 22570 3555 22610 3565
rect 22570 3535 22580 3555
rect 22600 3535 22610 3555
rect 22570 3525 22610 3535
rect 22665 3555 22745 3565
rect 22665 3535 22675 3555
rect 22695 3535 22715 3555
rect 22735 3535 22745 3555
rect 22665 3525 22745 3535
rect 22810 3555 22850 3565
rect 22810 3535 22820 3555
rect 22840 3535 22850 3555
rect 22810 3525 22850 3535
rect 22975 3555 23015 3565
rect 22975 3535 22985 3555
rect 23005 3535 23015 3555
rect 22975 3525 23015 3535
rect 23195 3555 23235 3565
rect 23195 3535 23205 3555
rect 23225 3535 23235 3555
rect 23195 3525 23235 3535
rect 23390 3555 23430 3565
rect 23390 3535 23400 3555
rect 23420 3535 23430 3555
rect 23390 3525 23430 3535
rect 23585 3555 23625 3565
rect 23585 3535 23595 3555
rect 23615 3535 23625 3555
rect 23585 3525 23625 3535
rect 23925 3555 23965 3565
rect 23925 3535 23935 3555
rect 23955 3535 23965 3555
rect 23925 3525 23965 3535
rect 25685 3530 25725 3540
rect 21635 3450 21655 3525
rect 22005 3450 22025 3525
rect 22085 3450 22105 3525
rect 22455 3450 22475 3525
rect 22580 3450 22600 3525
rect 22625 3500 22665 3505
rect 22625 3480 22635 3500
rect 22655 3480 22665 3500
rect 22625 3470 22665 3480
rect 22715 3450 22735 3525
rect 22825 3450 22845 3525
rect 22990 3450 23010 3525
rect 23205 3450 23225 3525
rect 23400 3450 23420 3525
rect 23595 3450 23615 3525
rect 23935 3450 23955 3525
rect 25100 3515 25140 3525
rect 25100 3495 25110 3515
rect 25130 3495 25140 3515
rect 25100 3485 25140 3495
rect 25480 3515 25520 3525
rect 25480 3495 25490 3515
rect 25510 3495 25520 3515
rect 25685 3510 25695 3530
rect 25715 3510 25725 3530
rect 25685 3500 25725 3510
rect 26035 3530 26075 3540
rect 26035 3510 26045 3530
rect 26065 3510 26075 3530
rect 26035 3500 26075 3510
rect 26370 3530 26425 3540
rect 25480 3465 25520 3495
rect 26370 3495 26380 3530
rect 26415 3495 26425 3530
rect 26370 3485 26425 3495
rect 24720 3455 24810 3465
rect 21590 3440 21660 3450
rect 21590 3420 21595 3440
rect 21615 3420 21635 3440
rect 21655 3420 21660 3440
rect 21590 3390 21660 3420
rect 21590 3370 21595 3390
rect 21615 3370 21635 3390
rect 21655 3370 21660 3390
rect 21590 3340 21660 3370
rect 21590 3320 21595 3340
rect 21615 3320 21635 3340
rect 21655 3320 21660 3340
rect 21590 3290 21660 3320
rect 21590 3270 21595 3290
rect 21615 3270 21635 3290
rect 21655 3270 21660 3290
rect 21590 3260 21660 3270
rect 21685 3440 21715 3450
rect 21685 3420 21690 3440
rect 21710 3420 21715 3440
rect 21685 3390 21715 3420
rect 21685 3370 21690 3390
rect 21710 3370 21715 3390
rect 21685 3340 21715 3370
rect 21685 3320 21690 3340
rect 21710 3320 21715 3340
rect 21685 3290 21715 3320
rect 21685 3270 21690 3290
rect 21710 3270 21715 3290
rect 21685 3260 21715 3270
rect 21740 3440 21830 3450
rect 21740 3420 21745 3440
rect 21765 3425 21800 3440
rect 21765 3420 21770 3425
rect 21740 3390 21770 3420
rect 21790 3420 21800 3425
rect 21820 3420 21830 3440
rect 21790 3410 21830 3420
rect 21850 3440 21920 3450
rect 21850 3430 21895 3440
rect 21740 3370 21745 3390
rect 21765 3370 21770 3390
rect 21740 3340 21770 3370
rect 21740 3320 21745 3340
rect 21765 3320 21770 3340
rect 21740 3290 21770 3320
rect 21740 3270 21745 3290
rect 21765 3270 21770 3290
rect 21740 3260 21770 3270
rect 21745 3240 21765 3260
rect 21685 3220 21765 3240
rect 21565 3210 21605 3220
rect 21565 3190 21575 3210
rect 21595 3190 21605 3210
rect 21565 3180 21605 3190
rect 21685 3140 21705 3220
rect 21850 3200 21870 3430
rect 21890 3420 21895 3430
rect 21915 3420 21920 3440
rect 21890 3390 21920 3420
rect 21890 3370 21895 3390
rect 21915 3370 21920 3390
rect 21890 3340 21920 3370
rect 21890 3320 21895 3340
rect 21915 3320 21920 3340
rect 21890 3290 21920 3320
rect 21890 3270 21895 3290
rect 21915 3270 21920 3290
rect 21890 3260 21920 3270
rect 21945 3440 21975 3450
rect 21945 3420 21950 3440
rect 21970 3420 21975 3440
rect 21945 3390 21975 3420
rect 21945 3370 21950 3390
rect 21970 3370 21975 3390
rect 21945 3340 21975 3370
rect 21945 3320 21950 3340
rect 21970 3320 21975 3340
rect 21945 3290 21975 3320
rect 21945 3270 21950 3290
rect 21970 3270 21975 3290
rect 21945 3260 21975 3270
rect 22000 3440 22110 3450
rect 22000 3420 22005 3440
rect 22025 3420 22045 3440
rect 22065 3420 22085 3440
rect 22105 3420 22110 3440
rect 22000 3390 22110 3420
rect 22000 3370 22005 3390
rect 22025 3370 22045 3390
rect 22065 3370 22085 3390
rect 22105 3370 22110 3390
rect 22000 3340 22110 3370
rect 22000 3320 22005 3340
rect 22025 3320 22045 3340
rect 22065 3320 22085 3340
rect 22105 3320 22110 3340
rect 22000 3290 22110 3320
rect 22000 3270 22005 3290
rect 22025 3270 22045 3290
rect 22065 3270 22085 3290
rect 22105 3270 22110 3290
rect 22000 3260 22110 3270
rect 22135 3440 22165 3450
rect 22135 3420 22140 3440
rect 22160 3420 22165 3440
rect 22135 3390 22165 3420
rect 22135 3370 22140 3390
rect 22160 3370 22165 3390
rect 22135 3340 22165 3370
rect 22135 3320 22140 3340
rect 22160 3320 22165 3340
rect 22135 3290 22165 3320
rect 22135 3270 22140 3290
rect 22160 3270 22165 3290
rect 22135 3260 22165 3270
rect 22190 3440 22280 3450
rect 22190 3420 22195 3440
rect 22215 3425 22250 3440
rect 22215 3420 22220 3425
rect 22190 3390 22220 3420
rect 22240 3420 22250 3425
rect 22270 3420 22280 3440
rect 22240 3410 22280 3420
rect 22300 3440 22370 3450
rect 22300 3430 22345 3440
rect 22190 3370 22195 3390
rect 22215 3370 22220 3390
rect 22190 3340 22220 3370
rect 22190 3320 22195 3340
rect 22215 3320 22220 3340
rect 22190 3290 22220 3320
rect 22190 3270 22195 3290
rect 22215 3270 22220 3290
rect 22190 3260 22220 3270
rect 21895 3240 21915 3260
rect 22195 3240 22215 3260
rect 21895 3220 21970 3240
rect 21730 3190 21870 3200
rect 21730 3170 21740 3190
rect 21760 3180 21870 3190
rect 21760 3170 21770 3180
rect 21730 3160 21770 3170
rect 21590 3130 21660 3140
rect 21590 3110 21595 3130
rect 21615 3110 21635 3130
rect 21655 3110 21660 3130
rect 21590 3080 21660 3110
rect 21590 3060 21595 3080
rect 21615 3060 21635 3080
rect 21655 3060 21660 3080
rect 21590 3050 21660 3060
rect 21685 3130 21715 3140
rect 21685 3110 21690 3130
rect 21710 3110 21715 3130
rect 21685 3080 21715 3110
rect 21685 3060 21690 3080
rect 21710 3060 21715 3080
rect 21685 3050 21715 3060
rect 21740 3130 21770 3140
rect 21740 3110 21745 3130
rect 21765 3110 21770 3130
rect 21740 3080 21770 3110
rect 21740 3060 21745 3080
rect 21765 3060 21770 3080
rect 21740 3050 21770 3060
rect 21635 2975 21655 3050
rect 21745 2975 21765 3050
rect 21850 3030 21870 3180
rect 21950 3140 21970 3220
rect 21990 3230 22215 3240
rect 21990 3210 22000 3230
rect 22020 3220 22215 3230
rect 22020 3210 22030 3220
rect 21990 3200 22030 3210
rect 22135 3140 22155 3220
rect 22300 3200 22320 3430
rect 22340 3420 22345 3430
rect 22365 3420 22370 3440
rect 22340 3390 22370 3420
rect 22340 3370 22345 3390
rect 22365 3370 22370 3390
rect 22340 3340 22370 3370
rect 22340 3320 22345 3340
rect 22365 3320 22370 3340
rect 22340 3290 22370 3320
rect 22340 3270 22345 3290
rect 22365 3270 22370 3290
rect 22340 3260 22370 3270
rect 22395 3440 22425 3450
rect 22395 3420 22400 3440
rect 22420 3420 22425 3440
rect 22395 3390 22425 3420
rect 22395 3370 22400 3390
rect 22420 3370 22425 3390
rect 22395 3340 22425 3370
rect 22395 3320 22400 3340
rect 22420 3320 22425 3340
rect 22395 3290 22425 3320
rect 22395 3270 22400 3290
rect 22420 3270 22425 3290
rect 22395 3260 22425 3270
rect 22450 3440 22520 3450
rect 22450 3420 22455 3440
rect 22475 3420 22495 3440
rect 22515 3420 22520 3440
rect 22450 3390 22520 3420
rect 22450 3370 22455 3390
rect 22475 3370 22495 3390
rect 22515 3370 22520 3390
rect 22450 3340 22520 3370
rect 22450 3320 22455 3340
rect 22475 3320 22495 3340
rect 22515 3320 22520 3340
rect 22450 3290 22520 3320
rect 22450 3270 22455 3290
rect 22475 3270 22495 3290
rect 22515 3270 22520 3290
rect 22450 3260 22520 3270
rect 22560 3440 22630 3450
rect 22560 3420 22565 3440
rect 22585 3420 22605 3440
rect 22625 3420 22630 3440
rect 22560 3390 22630 3420
rect 22560 3370 22565 3390
rect 22585 3370 22605 3390
rect 22625 3370 22630 3390
rect 22560 3340 22630 3370
rect 22560 3320 22565 3340
rect 22585 3320 22605 3340
rect 22625 3320 22630 3340
rect 22560 3290 22630 3320
rect 22560 3270 22565 3290
rect 22585 3270 22605 3290
rect 22625 3270 22630 3290
rect 22560 3260 22630 3270
rect 22655 3440 22685 3450
rect 22655 3420 22660 3440
rect 22680 3420 22685 3440
rect 22655 3390 22685 3420
rect 22655 3370 22660 3390
rect 22680 3370 22685 3390
rect 22655 3340 22685 3370
rect 22655 3320 22660 3340
rect 22680 3320 22685 3340
rect 22655 3290 22685 3320
rect 22655 3270 22660 3290
rect 22680 3270 22685 3290
rect 22655 3260 22685 3270
rect 22710 3440 22740 3450
rect 22710 3420 22715 3440
rect 22735 3420 22740 3440
rect 22710 3390 22740 3420
rect 22710 3370 22715 3390
rect 22735 3370 22740 3390
rect 22710 3340 22740 3370
rect 22710 3320 22715 3340
rect 22735 3320 22740 3340
rect 22710 3290 22740 3320
rect 22710 3270 22715 3290
rect 22735 3270 22740 3290
rect 22710 3260 22740 3270
rect 22780 3440 22850 3450
rect 22780 3420 22785 3440
rect 22805 3420 22825 3440
rect 22845 3420 22850 3440
rect 22780 3390 22850 3420
rect 22780 3370 22785 3390
rect 22805 3370 22825 3390
rect 22845 3370 22850 3390
rect 22780 3340 22850 3370
rect 22780 3320 22785 3340
rect 22805 3320 22825 3340
rect 22845 3320 22850 3340
rect 22780 3290 22850 3320
rect 22780 3270 22785 3290
rect 22805 3270 22825 3290
rect 22845 3270 22850 3290
rect 22780 3260 22850 3270
rect 22875 3440 22905 3450
rect 22875 3420 22880 3440
rect 22900 3420 22905 3440
rect 22875 3390 22905 3420
rect 22875 3370 22880 3390
rect 22900 3370 22905 3390
rect 22875 3340 22905 3370
rect 22875 3320 22880 3340
rect 22900 3320 22905 3340
rect 22875 3290 22905 3320
rect 22875 3270 22880 3290
rect 22900 3270 22905 3290
rect 22875 3260 22905 3270
rect 22945 3440 23015 3450
rect 22945 3420 22950 3440
rect 22970 3420 22990 3440
rect 23010 3420 23015 3440
rect 22945 3390 23015 3420
rect 22945 3370 22950 3390
rect 22970 3370 22990 3390
rect 23010 3370 23015 3390
rect 22945 3340 23015 3370
rect 22945 3320 22950 3340
rect 22970 3320 22990 3340
rect 23010 3320 23015 3340
rect 22945 3290 23015 3320
rect 22945 3270 22950 3290
rect 22970 3270 22990 3290
rect 23010 3270 23015 3290
rect 22945 3260 23015 3270
rect 23040 3440 23070 3450
rect 23040 3420 23045 3440
rect 23065 3420 23070 3440
rect 23040 3390 23070 3420
rect 23040 3370 23045 3390
rect 23065 3370 23070 3390
rect 23040 3340 23070 3370
rect 23040 3320 23045 3340
rect 23065 3320 23070 3340
rect 23040 3290 23070 3320
rect 23040 3270 23045 3290
rect 23065 3270 23070 3290
rect 23040 3260 23070 3270
rect 23145 3440 23235 3450
rect 23145 3420 23155 3440
rect 23175 3420 23205 3440
rect 23225 3420 23235 3440
rect 23145 3390 23235 3420
rect 23145 3370 23155 3390
rect 23175 3370 23205 3390
rect 23225 3370 23235 3390
rect 23145 3340 23235 3370
rect 23145 3320 23155 3340
rect 23175 3320 23205 3340
rect 23225 3320 23235 3340
rect 23145 3290 23235 3320
rect 23145 3270 23155 3290
rect 23175 3270 23205 3290
rect 23225 3270 23235 3290
rect 23145 3260 23235 3270
rect 23260 3440 23300 3450
rect 23260 3420 23270 3440
rect 23290 3420 23300 3440
rect 23260 3390 23300 3420
rect 23260 3370 23270 3390
rect 23290 3370 23300 3390
rect 23260 3340 23300 3370
rect 23260 3320 23270 3340
rect 23290 3320 23300 3340
rect 23260 3290 23300 3320
rect 23260 3270 23270 3290
rect 23290 3270 23300 3290
rect 23260 3260 23300 3270
rect 23340 3440 23430 3450
rect 23340 3420 23350 3440
rect 23370 3420 23400 3440
rect 23420 3420 23430 3440
rect 23340 3390 23430 3420
rect 23340 3370 23350 3390
rect 23370 3370 23400 3390
rect 23420 3370 23430 3390
rect 23340 3340 23430 3370
rect 23340 3320 23350 3340
rect 23370 3320 23400 3340
rect 23420 3320 23430 3340
rect 23340 3290 23430 3320
rect 23340 3270 23350 3290
rect 23370 3270 23400 3290
rect 23420 3270 23430 3290
rect 23340 3260 23430 3270
rect 23455 3440 23495 3450
rect 23455 3420 23465 3440
rect 23485 3420 23495 3440
rect 23455 3390 23495 3420
rect 23455 3370 23465 3390
rect 23485 3370 23495 3390
rect 23455 3340 23495 3370
rect 23455 3320 23465 3340
rect 23485 3320 23495 3340
rect 23455 3290 23495 3320
rect 23455 3270 23465 3290
rect 23485 3270 23495 3290
rect 23455 3260 23495 3270
rect 23535 3440 23625 3450
rect 23535 3420 23545 3440
rect 23565 3420 23595 3440
rect 23615 3420 23625 3440
rect 23535 3390 23625 3420
rect 23535 3370 23545 3390
rect 23565 3370 23595 3390
rect 23615 3370 23625 3390
rect 23535 3340 23625 3370
rect 23535 3320 23545 3340
rect 23565 3320 23595 3340
rect 23615 3320 23625 3340
rect 23535 3290 23625 3320
rect 23535 3270 23545 3290
rect 23565 3270 23595 3290
rect 23615 3270 23625 3290
rect 23535 3260 23625 3270
rect 23650 3440 23690 3450
rect 23650 3420 23660 3440
rect 23680 3420 23690 3440
rect 23650 3390 23690 3420
rect 23650 3370 23660 3390
rect 23680 3370 23690 3390
rect 23650 3340 23690 3370
rect 23650 3320 23660 3340
rect 23680 3320 23690 3340
rect 23650 3290 23690 3320
rect 23650 3270 23660 3290
rect 23680 3270 23690 3290
rect 23650 3260 23690 3270
rect 23730 3440 23770 3450
rect 23730 3420 23740 3440
rect 23760 3420 23770 3440
rect 23730 3390 23770 3420
rect 23730 3370 23740 3390
rect 23760 3370 23770 3390
rect 23730 3340 23770 3370
rect 23730 3320 23740 3340
rect 23760 3320 23770 3340
rect 23730 3290 23770 3320
rect 23730 3270 23740 3290
rect 23760 3270 23770 3290
rect 23730 3260 23770 3270
rect 23795 3440 23835 3450
rect 23795 3420 23805 3440
rect 23825 3420 23835 3440
rect 23795 3390 23835 3420
rect 23795 3370 23805 3390
rect 23825 3370 23835 3390
rect 23795 3340 23835 3370
rect 23795 3320 23805 3340
rect 23825 3320 23835 3340
rect 23795 3290 23835 3320
rect 23795 3270 23805 3290
rect 23825 3270 23835 3290
rect 23795 3260 23835 3270
rect 23875 3440 23965 3450
rect 23875 3420 23885 3440
rect 23905 3420 23935 3440
rect 23955 3420 23965 3440
rect 23875 3390 23965 3420
rect 23875 3370 23885 3390
rect 23905 3370 23935 3390
rect 23955 3370 23965 3390
rect 23875 3340 23965 3370
rect 23875 3320 23885 3340
rect 23905 3320 23935 3340
rect 23955 3320 23965 3340
rect 23875 3290 23965 3320
rect 23875 3270 23885 3290
rect 23905 3270 23935 3290
rect 23955 3270 23965 3290
rect 23875 3260 23965 3270
rect 23990 3440 24030 3450
rect 23990 3420 24000 3440
rect 24020 3420 24030 3440
rect 23990 3390 24030 3420
rect 23990 3370 24000 3390
rect 24020 3370 24030 3390
rect 23990 3340 24030 3370
rect 23990 3320 24000 3340
rect 24020 3320 24030 3340
rect 23990 3290 24030 3320
rect 23990 3270 24000 3290
rect 24020 3270 24030 3290
rect 24720 3435 24730 3455
rect 24750 3435 24780 3455
rect 24800 3435 24810 3455
rect 24720 3405 24810 3435
rect 24720 3385 24730 3405
rect 24750 3385 24780 3405
rect 24800 3385 24810 3405
rect 24720 3355 24810 3385
rect 24720 3335 24730 3355
rect 24750 3335 24780 3355
rect 24800 3335 24810 3355
rect 24720 3305 24810 3335
rect 24720 3285 24730 3305
rect 24750 3285 24780 3305
rect 24800 3285 24810 3305
rect 24720 3275 24810 3285
rect 24880 3455 24920 3465
rect 24880 3435 24890 3455
rect 24910 3435 24920 3455
rect 24880 3405 24920 3435
rect 24880 3385 24890 3405
rect 24910 3385 24920 3405
rect 24880 3355 24920 3385
rect 24880 3335 24890 3355
rect 24910 3335 24920 3355
rect 24880 3305 24920 3335
rect 24880 3285 24890 3305
rect 24910 3285 24920 3305
rect 24880 3275 24920 3285
rect 24990 3455 25030 3465
rect 24990 3435 25000 3455
rect 25020 3435 25030 3455
rect 24990 3405 25030 3435
rect 24990 3385 25000 3405
rect 25020 3385 25030 3405
rect 24990 3355 25030 3385
rect 24990 3335 25000 3355
rect 25020 3335 25030 3355
rect 24990 3305 25030 3335
rect 24990 3285 25000 3305
rect 25020 3285 25030 3305
rect 24990 3275 25030 3285
rect 25100 3455 25140 3465
rect 25100 3435 25110 3455
rect 25130 3435 25140 3455
rect 25100 3405 25140 3435
rect 25100 3385 25110 3405
rect 25130 3385 25140 3405
rect 25100 3355 25140 3385
rect 25100 3335 25110 3355
rect 25130 3335 25140 3355
rect 25100 3305 25140 3335
rect 25100 3285 25110 3305
rect 25130 3285 25140 3305
rect 25100 3275 25140 3285
rect 25210 3455 25250 3465
rect 25210 3435 25220 3455
rect 25240 3435 25250 3455
rect 25210 3405 25250 3435
rect 25210 3385 25220 3405
rect 25240 3385 25250 3405
rect 25210 3355 25250 3385
rect 25210 3335 25220 3355
rect 25240 3335 25250 3355
rect 25210 3305 25250 3335
rect 25210 3285 25220 3305
rect 25240 3285 25250 3305
rect 25210 3275 25250 3285
rect 25320 3455 25360 3465
rect 25320 3435 25330 3455
rect 25350 3435 25360 3455
rect 25320 3405 25360 3435
rect 25320 3385 25330 3405
rect 25350 3385 25360 3405
rect 25320 3355 25360 3385
rect 25320 3335 25330 3355
rect 25350 3335 25360 3355
rect 25320 3305 25360 3335
rect 25320 3285 25330 3305
rect 25350 3285 25360 3305
rect 25320 3275 25360 3285
rect 25430 3455 25570 3465
rect 25430 3435 25440 3455
rect 25460 3435 25490 3455
rect 25510 3435 25540 3455
rect 25560 3435 25570 3455
rect 25430 3405 25570 3435
rect 25430 3385 25440 3405
rect 25460 3385 25490 3405
rect 25510 3385 25540 3405
rect 25560 3385 25570 3405
rect 25430 3355 25570 3385
rect 25430 3335 25440 3355
rect 25460 3335 25490 3355
rect 25510 3335 25540 3355
rect 25560 3335 25570 3355
rect 25430 3305 25570 3335
rect 25430 3285 25440 3305
rect 25460 3285 25490 3305
rect 25510 3285 25540 3305
rect 25560 3285 25570 3305
rect 25430 3275 25570 3285
rect 25640 3455 25680 3465
rect 25640 3435 25650 3455
rect 25670 3435 25680 3455
rect 25640 3405 25680 3435
rect 25640 3385 25650 3405
rect 25670 3385 25680 3405
rect 25640 3355 25680 3385
rect 25640 3335 25650 3355
rect 25670 3335 25680 3355
rect 25640 3305 25680 3335
rect 25640 3285 25650 3305
rect 25670 3285 25680 3305
rect 25640 3275 25680 3285
rect 25750 3455 25790 3465
rect 25750 3435 25760 3455
rect 25780 3435 25790 3455
rect 25750 3405 25790 3435
rect 25750 3385 25760 3405
rect 25780 3385 25790 3405
rect 25750 3355 25790 3385
rect 25750 3335 25760 3355
rect 25780 3335 25790 3355
rect 25750 3305 25790 3335
rect 25750 3285 25760 3305
rect 25780 3285 25790 3305
rect 25750 3275 25790 3285
rect 25860 3455 25900 3465
rect 25860 3435 25870 3455
rect 25890 3435 25900 3455
rect 25860 3405 25900 3435
rect 25860 3385 25870 3405
rect 25890 3385 25900 3405
rect 25860 3355 25900 3385
rect 25860 3335 25870 3355
rect 25890 3335 25900 3355
rect 25860 3305 25900 3335
rect 25860 3285 25870 3305
rect 25890 3285 25900 3305
rect 25860 3275 25900 3285
rect 25970 3455 26010 3465
rect 25970 3435 25980 3455
rect 26000 3435 26010 3455
rect 25970 3405 26010 3435
rect 25970 3385 25980 3405
rect 26000 3385 26010 3405
rect 25970 3355 26010 3385
rect 25970 3335 25980 3355
rect 26000 3335 26010 3355
rect 25970 3305 26010 3335
rect 25970 3285 25980 3305
rect 26000 3285 26010 3305
rect 25970 3275 26010 3285
rect 26080 3455 26120 3465
rect 26080 3435 26090 3455
rect 26110 3435 26120 3455
rect 26080 3405 26120 3435
rect 26080 3385 26090 3405
rect 26110 3385 26120 3405
rect 26080 3355 26120 3385
rect 26080 3335 26090 3355
rect 26110 3335 26120 3355
rect 26080 3305 26120 3335
rect 26080 3285 26090 3305
rect 26110 3285 26120 3305
rect 26080 3275 26120 3285
rect 26190 3455 26280 3465
rect 26190 3435 26200 3455
rect 26220 3435 26250 3455
rect 26270 3435 26280 3455
rect 26190 3405 26280 3435
rect 26190 3385 26200 3405
rect 26220 3385 26250 3405
rect 26270 3385 26280 3405
rect 26190 3355 26280 3385
rect 26190 3335 26200 3355
rect 26220 3335 26250 3355
rect 26270 3335 26280 3355
rect 26190 3305 26280 3335
rect 26190 3285 26200 3305
rect 26220 3285 26250 3305
rect 26270 3285 26280 3305
rect 26190 3275 26280 3285
rect 23990 3260 24030 3270
rect 22345 3240 22365 3260
rect 22345 3220 22420 3240
rect 22180 3190 22320 3200
rect 22180 3170 22190 3190
rect 22210 3180 22320 3190
rect 22210 3170 22220 3180
rect 22180 3160 22220 3170
rect 22400 3140 22420 3220
rect 22660 3225 22680 3260
rect 22885 3225 22905 3260
rect 23050 3225 23070 3260
rect 22660 3215 22770 3225
rect 22660 3205 22740 3215
rect 22515 3195 22555 3205
rect 22515 3175 22525 3195
rect 22545 3175 22555 3195
rect 22515 3165 22555 3175
rect 22715 3195 22740 3205
rect 22760 3195 22770 3215
rect 22715 3185 22770 3195
rect 22885 3215 22935 3225
rect 22885 3195 22905 3215
rect 22925 3195 22935 3215
rect 22885 3185 22935 3195
rect 23050 3215 23100 3225
rect 23050 3195 23070 3215
rect 23090 3195 23100 3215
rect 23280 3215 23300 3260
rect 23410 3215 23450 3225
rect 23050 3185 23100 3195
rect 23125 3200 23165 3210
rect 22715 3140 22735 3185
rect 22885 3140 22905 3185
rect 23050 3140 23070 3185
rect 23125 3180 23135 3200
rect 23155 3180 23165 3200
rect 23125 3170 23165 3180
rect 23280 3195 23420 3215
rect 23440 3195 23450 3215
rect 23280 3140 23300 3195
rect 23410 3185 23450 3195
rect 23475 3200 23495 3260
rect 23670 3240 23690 3260
rect 23670 3230 23710 3240
rect 23670 3210 23680 3230
rect 23700 3210 23710 3230
rect 23670 3200 23710 3210
rect 23475 3190 23645 3200
rect 23475 3180 23615 3190
rect 23475 3140 23495 3180
rect 23605 3170 23615 3180
rect 23635 3170 23645 3190
rect 23605 3160 23645 3170
rect 23670 3140 23690 3200
rect 23740 3140 23760 3260
rect 23805 3180 23825 3260
rect 23845 3230 23885 3240
rect 23845 3210 23855 3230
rect 23875 3210 23885 3230
rect 23845 3200 23885 3210
rect 24000 3200 24020 3260
rect 24770 3245 24810 3255
rect 24770 3225 24780 3245
rect 24800 3225 24810 3245
rect 24770 3215 24810 3225
rect 26190 3245 26230 3255
rect 26190 3225 26200 3245
rect 26220 3225 26230 3245
rect 26190 3215 26230 3225
rect 24000 3190 24040 3200
rect 24000 3180 24010 3190
rect 23805 3170 24010 3180
rect 24030 3170 24040 3190
rect 23805 3160 24040 3170
rect 23805 3140 23825 3160
rect 21890 3130 21920 3140
rect 21890 3110 21895 3130
rect 21915 3110 21920 3130
rect 21890 3080 21920 3110
rect 21890 3060 21895 3080
rect 21915 3060 21920 3080
rect 21890 3050 21920 3060
rect 21945 3130 21975 3140
rect 21945 3110 21950 3130
rect 21970 3110 21975 3130
rect 21945 3080 21975 3110
rect 21945 3060 21950 3080
rect 21970 3060 21975 3080
rect 21945 3050 21975 3060
rect 22000 3130 22110 3140
rect 22000 3110 22005 3130
rect 22025 3110 22045 3130
rect 22065 3110 22085 3130
rect 22105 3110 22110 3130
rect 22000 3080 22110 3110
rect 22000 3060 22005 3080
rect 22025 3060 22045 3080
rect 22065 3060 22085 3080
rect 22105 3060 22110 3080
rect 22000 3050 22110 3060
rect 22135 3130 22165 3140
rect 22135 3110 22140 3130
rect 22160 3110 22165 3130
rect 22135 3080 22165 3110
rect 22135 3060 22140 3080
rect 22160 3060 22165 3080
rect 22135 3050 22165 3060
rect 22190 3130 22220 3140
rect 22190 3110 22195 3130
rect 22215 3110 22220 3130
rect 22190 3080 22220 3110
rect 22190 3060 22195 3080
rect 22215 3060 22220 3080
rect 22190 3050 22220 3060
rect 22340 3130 22370 3140
rect 22340 3110 22345 3130
rect 22365 3110 22370 3130
rect 22340 3080 22370 3110
rect 22340 3060 22345 3080
rect 22365 3060 22370 3080
rect 22340 3050 22370 3060
rect 22395 3130 22425 3140
rect 22395 3110 22400 3130
rect 22420 3110 22425 3130
rect 22395 3080 22425 3110
rect 22395 3060 22400 3080
rect 22420 3060 22425 3080
rect 22395 3050 22425 3060
rect 22450 3130 22520 3140
rect 22450 3110 22455 3130
rect 22475 3110 22495 3130
rect 22515 3110 22520 3130
rect 22450 3080 22520 3110
rect 22450 3060 22455 3080
rect 22475 3060 22495 3080
rect 22515 3060 22520 3080
rect 22450 3050 22520 3060
rect 22560 3130 22630 3140
rect 22560 3110 22565 3130
rect 22585 3110 22605 3130
rect 22625 3110 22630 3130
rect 22560 3080 22630 3110
rect 22560 3060 22565 3080
rect 22585 3060 22605 3080
rect 22625 3060 22630 3080
rect 22560 3050 22630 3060
rect 22655 3130 22685 3140
rect 22655 3110 22660 3130
rect 22680 3110 22685 3130
rect 22655 3080 22685 3110
rect 22655 3060 22660 3080
rect 22680 3060 22685 3080
rect 22655 3050 22685 3060
rect 22710 3130 22740 3140
rect 22710 3110 22715 3130
rect 22735 3110 22740 3130
rect 22710 3080 22740 3110
rect 22710 3060 22715 3080
rect 22735 3060 22740 3080
rect 22710 3050 22740 3060
rect 22780 3130 22850 3140
rect 22780 3110 22785 3130
rect 22805 3110 22825 3130
rect 22845 3110 22850 3130
rect 22780 3080 22850 3110
rect 22780 3060 22785 3080
rect 22805 3060 22825 3080
rect 22845 3060 22850 3080
rect 22780 3050 22850 3060
rect 22875 3130 22905 3140
rect 22875 3110 22880 3130
rect 22900 3110 22905 3130
rect 22875 3080 22905 3110
rect 22875 3060 22880 3080
rect 22900 3060 22905 3080
rect 22875 3050 22905 3060
rect 22945 3130 23015 3140
rect 22945 3110 22950 3130
rect 22970 3110 22990 3130
rect 23010 3110 23015 3130
rect 22945 3080 23015 3110
rect 22945 3060 22950 3080
rect 22970 3060 22990 3080
rect 23010 3060 23015 3080
rect 22945 3050 23015 3060
rect 23040 3130 23070 3140
rect 23040 3110 23045 3130
rect 23065 3110 23070 3130
rect 23040 3080 23070 3110
rect 23040 3060 23045 3080
rect 23065 3060 23070 3080
rect 23040 3050 23070 3060
rect 23155 3130 23235 3140
rect 23155 3110 23160 3130
rect 23180 3110 23205 3130
rect 23225 3110 23235 3130
rect 23155 3080 23235 3110
rect 23155 3060 23160 3080
rect 23180 3060 23205 3080
rect 23225 3060 23235 3080
rect 23155 3050 23235 3060
rect 23260 3130 23300 3140
rect 23260 3110 23270 3130
rect 23290 3110 23300 3130
rect 23260 3080 23300 3110
rect 23260 3060 23270 3080
rect 23290 3060 23300 3080
rect 23260 3050 23300 3060
rect 23350 3130 23430 3140
rect 23350 3110 23355 3130
rect 23375 3110 23400 3130
rect 23420 3110 23430 3130
rect 23350 3080 23430 3110
rect 23350 3060 23355 3080
rect 23375 3060 23400 3080
rect 23420 3060 23430 3080
rect 23350 3050 23430 3060
rect 23455 3130 23495 3140
rect 23455 3110 23465 3130
rect 23485 3110 23495 3130
rect 23455 3080 23495 3110
rect 23455 3060 23465 3080
rect 23485 3060 23495 3080
rect 23455 3050 23495 3060
rect 23545 3130 23625 3140
rect 23545 3110 23550 3130
rect 23570 3110 23595 3130
rect 23615 3110 23625 3130
rect 23545 3080 23625 3110
rect 23545 3060 23550 3080
rect 23570 3060 23595 3080
rect 23615 3060 23625 3080
rect 23545 3050 23625 3060
rect 23650 3130 23690 3140
rect 23650 3110 23660 3130
rect 23680 3110 23690 3130
rect 23650 3080 23690 3110
rect 23650 3060 23660 3080
rect 23680 3060 23690 3080
rect 23650 3050 23690 3060
rect 23730 3130 23770 3140
rect 23730 3110 23740 3130
rect 23760 3110 23770 3130
rect 23730 3080 23770 3110
rect 23730 3060 23740 3080
rect 23760 3060 23770 3080
rect 23730 3050 23770 3060
rect 23795 3130 23835 3140
rect 23795 3110 23805 3130
rect 23825 3110 23835 3130
rect 23795 3080 23835 3110
rect 23795 3060 23805 3080
rect 23825 3060 23835 3080
rect 23795 3050 23835 3060
rect 21830 3020 21870 3030
rect 21830 3000 21840 3020
rect 21860 3000 21870 3020
rect 21830 2990 21870 3000
rect 21895 2975 21915 3050
rect 22005 2975 22025 3050
rect 22085 2975 22105 3050
rect 22195 2975 22215 3050
rect 22345 2975 22365 3050
rect 22455 2975 22475 3050
rect 22605 2975 22625 3050
rect 22690 3020 22730 3030
rect 22690 3000 22700 3020
rect 22720 3000 22730 3020
rect 22690 2990 22730 3000
rect 22825 2975 22845 3050
rect 22990 2975 23010 3050
rect 23205 2975 23225 3050
rect 23400 2975 23420 3050
rect 23595 2975 23615 3050
rect 23740 3030 23760 3050
rect 23730 3020 23770 3030
rect 23730 3000 23740 3020
rect 23760 3000 23770 3020
rect 23730 2990 23770 3000
rect 21625 2965 21665 2975
rect 21625 2945 21635 2965
rect 21655 2945 21665 2965
rect 21625 2935 21665 2945
rect 21735 2965 21775 2975
rect 21735 2945 21745 2965
rect 21765 2945 21775 2965
rect 21735 2935 21775 2945
rect 21885 2965 21925 2975
rect 21885 2945 21895 2965
rect 21915 2945 21925 2965
rect 21885 2935 21925 2945
rect 21995 2965 22035 2975
rect 21995 2945 22005 2965
rect 22025 2945 22035 2965
rect 21995 2935 22035 2945
rect 22075 2965 22115 2975
rect 22075 2945 22085 2965
rect 22105 2945 22115 2965
rect 22075 2935 22115 2945
rect 22185 2965 22225 2975
rect 22185 2945 22195 2965
rect 22215 2945 22225 2965
rect 22185 2935 22225 2945
rect 22335 2965 22375 2975
rect 22335 2945 22345 2965
rect 22365 2945 22375 2965
rect 22335 2935 22375 2945
rect 22445 2965 22485 2975
rect 22445 2945 22455 2965
rect 22475 2945 22485 2965
rect 22445 2935 22485 2945
rect 22595 2965 22635 2975
rect 22595 2945 22605 2965
rect 22625 2945 22635 2965
rect 22595 2935 22635 2945
rect 22815 2965 22855 2975
rect 22815 2945 22825 2965
rect 22845 2945 22855 2965
rect 22815 2935 22855 2945
rect 22980 2965 23020 2975
rect 22980 2945 22990 2965
rect 23010 2945 23020 2965
rect 22980 2935 23020 2945
rect 23195 2965 23235 2975
rect 23195 2945 23205 2965
rect 23225 2945 23235 2965
rect 23195 2935 23235 2945
rect 23390 2965 23430 2975
rect 23390 2945 23400 2965
rect 23420 2945 23430 2965
rect 23390 2935 23430 2945
rect 23585 2965 23625 2975
rect 23585 2945 23595 2965
rect 23615 2945 23625 2965
rect 23585 2935 23625 2945
rect 26490 2940 26545 2950
rect 26490 2905 26500 2940
rect 26535 2905 26545 2940
rect 26490 2895 26545 2905
<< viali >>
rect 26555 4155 26590 4190
rect 21635 4125 21655 4145
rect 21745 4125 21765 4145
rect 21895 4125 21915 4145
rect 22010 4125 22030 4145
rect 22085 4125 22105 4145
rect 22195 4125 22215 4145
rect 22345 4125 22365 4145
rect 22455 4125 22475 4145
rect 22655 4125 22675 4145
rect 22820 4125 22840 4145
rect 22985 4125 23005 4145
rect 23205 4125 23225 4145
rect 23595 4125 23615 4145
rect 23935 4125 23955 4145
rect 23460 4070 23480 4090
rect 23775 4070 23795 4090
rect 24680 4045 24700 4065
rect 26200 4045 26220 4065
rect 24680 3985 24700 4005
rect 21575 3880 21595 3900
rect 22535 3875 22555 3895
rect 23050 3875 23070 3895
rect 23125 3880 23145 3900
rect 24680 3935 24700 3955
rect 24010 3900 24030 3920
rect 24680 3885 24700 3905
rect 24680 3835 24700 3855
rect 24790 3985 24810 4005
rect 24790 3935 24810 3955
rect 24790 3885 24810 3905
rect 24790 3835 24810 3855
rect 24900 3985 24920 4005
rect 24900 3935 24920 3955
rect 24900 3885 24920 3905
rect 24900 3835 24920 3855
rect 25010 3985 25030 4005
rect 25010 3935 25030 3955
rect 25010 3885 25030 3905
rect 25010 3835 25030 3855
rect 25120 3985 25140 4005
rect 25170 3985 25190 4005
rect 25220 3985 25240 4005
rect 25120 3935 25140 3955
rect 25170 3935 25190 3955
rect 25220 3935 25240 3955
rect 25120 3885 25140 3905
rect 25170 3885 25190 3905
rect 25220 3885 25240 3905
rect 25120 3835 25140 3855
rect 25170 3835 25190 3855
rect 25220 3835 25240 3855
rect 25330 3985 25350 4005
rect 25330 3935 25350 3955
rect 25330 3885 25350 3905
rect 25330 3835 25350 3855
rect 25440 3985 25460 4005
rect 25440 3935 25460 3955
rect 25440 3885 25460 3905
rect 25440 3835 25460 3855
rect 25550 3985 25570 4005
rect 25550 3935 25570 3955
rect 25550 3885 25570 3905
rect 25550 3835 25570 3855
rect 25660 3985 25680 4005
rect 25710 3985 25730 4005
rect 25760 3985 25780 4005
rect 25660 3935 25680 3955
rect 25710 3935 25730 3955
rect 25760 3935 25780 3955
rect 25660 3885 25680 3905
rect 25710 3885 25730 3905
rect 25760 3885 25780 3905
rect 25660 3835 25680 3855
rect 25710 3835 25730 3855
rect 25760 3835 25780 3855
rect 25870 3985 25890 4005
rect 25870 3935 25890 3955
rect 25870 3885 25890 3905
rect 25870 3835 25890 3855
rect 25980 3985 26000 4005
rect 25980 3935 26000 3955
rect 25980 3885 26000 3905
rect 25980 3835 26000 3855
rect 26090 3985 26110 4005
rect 26090 3935 26110 3955
rect 26090 3885 26110 3905
rect 26090 3835 26110 3855
rect 26200 3985 26220 4005
rect 26200 3935 26220 3955
rect 26200 3885 26220 3905
rect 26200 3835 26220 3855
rect 24900 3780 24920 3800
rect 25915 3760 25935 3780
rect 26045 3760 26065 3780
rect 26380 3760 26415 3795
rect 21860 3590 21880 3610
rect 23420 3590 23440 3610
rect 23740 3590 23760 3610
rect 21635 3535 21655 3555
rect 22005 3535 22025 3555
rect 22085 3535 22105 3555
rect 22455 3535 22475 3555
rect 22580 3535 22600 3555
rect 22675 3535 22695 3555
rect 22715 3535 22735 3555
rect 22820 3535 22840 3555
rect 22985 3535 23005 3555
rect 23205 3535 23225 3555
rect 23400 3535 23420 3555
rect 23595 3535 23615 3555
rect 23935 3535 23955 3555
rect 22635 3480 22655 3500
rect 25110 3495 25130 3515
rect 25695 3510 25715 3530
rect 26045 3510 26065 3530
rect 26380 3495 26415 3530
rect 21575 3190 21595 3210
rect 24780 3435 24800 3455
rect 24780 3385 24800 3405
rect 24780 3335 24800 3355
rect 24780 3285 24800 3305
rect 24890 3435 24910 3455
rect 24890 3385 24910 3405
rect 24890 3335 24910 3355
rect 24890 3285 24910 3305
rect 25000 3435 25020 3455
rect 25000 3385 25020 3405
rect 25000 3335 25020 3355
rect 25000 3285 25020 3305
rect 25110 3435 25130 3455
rect 25110 3385 25130 3405
rect 25110 3335 25130 3355
rect 25110 3285 25130 3305
rect 25220 3435 25240 3455
rect 25220 3385 25240 3405
rect 25220 3335 25240 3355
rect 25220 3285 25240 3305
rect 25330 3435 25350 3455
rect 25330 3385 25350 3405
rect 25330 3335 25350 3355
rect 25330 3285 25350 3305
rect 25440 3435 25460 3455
rect 25490 3435 25510 3455
rect 25540 3435 25560 3455
rect 25440 3385 25460 3405
rect 25490 3385 25510 3405
rect 25540 3385 25560 3405
rect 25440 3335 25460 3355
rect 25490 3335 25510 3355
rect 25540 3335 25560 3355
rect 25440 3285 25460 3305
rect 25490 3285 25510 3305
rect 25540 3285 25560 3305
rect 25650 3435 25670 3455
rect 25650 3385 25670 3405
rect 25650 3335 25670 3355
rect 25650 3285 25670 3305
rect 25760 3435 25780 3455
rect 25760 3385 25780 3405
rect 25760 3335 25780 3355
rect 25760 3285 25780 3305
rect 25870 3435 25890 3455
rect 25870 3385 25890 3405
rect 25870 3335 25890 3355
rect 25870 3285 25890 3305
rect 25980 3435 26000 3455
rect 25980 3385 26000 3405
rect 25980 3335 26000 3355
rect 25980 3285 26000 3305
rect 26090 3435 26110 3455
rect 26090 3385 26110 3405
rect 26090 3335 26110 3355
rect 26090 3285 26110 3305
rect 26200 3435 26220 3455
rect 26200 3385 26220 3405
rect 26200 3335 26220 3355
rect 26200 3285 26220 3305
rect 22525 3175 22545 3195
rect 23070 3195 23090 3215
rect 23135 3180 23155 3200
rect 23855 3210 23875 3230
rect 24780 3225 24800 3245
rect 26200 3225 26220 3245
rect 24010 3170 24030 3190
rect 21840 3000 21860 3020
rect 22700 3000 22720 3020
rect 23740 3000 23760 3020
rect 21635 2945 21655 2965
rect 21745 2945 21765 2965
rect 21895 2945 21915 2965
rect 22005 2945 22025 2965
rect 22085 2945 22105 2965
rect 22195 2945 22215 2965
rect 22345 2945 22365 2965
rect 22455 2945 22475 2965
rect 22605 2945 22625 2965
rect 22825 2945 22845 2965
rect 22990 2945 23010 2965
rect 23205 2945 23225 2965
rect 23400 2945 23420 2965
rect 23595 2945 23615 2965
rect 26500 2905 26535 2940
<< metal1 >>
rect 26545 4190 26600 4200
rect 24050 4185 24090 4190
rect 24050 4155 24055 4185
rect 24085 4155 24090 4185
rect 21625 4150 21665 4155
rect 21625 4120 21630 4150
rect 21660 4120 21665 4150
rect 21625 4115 21665 4120
rect 21735 4150 21775 4155
rect 21735 4120 21740 4150
rect 21770 4120 21775 4150
rect 21735 4115 21775 4120
rect 21885 4150 21925 4155
rect 21885 4120 21890 4150
rect 21920 4120 21925 4150
rect 21885 4115 21925 4120
rect 22000 4150 22040 4155
rect 22000 4120 22005 4150
rect 22035 4120 22040 4150
rect 22000 4115 22040 4120
rect 22075 4150 22115 4155
rect 22075 4120 22080 4150
rect 22110 4120 22115 4150
rect 22075 4115 22115 4120
rect 22185 4150 22225 4155
rect 22185 4120 22190 4150
rect 22220 4120 22225 4150
rect 22185 4115 22225 4120
rect 22335 4150 22375 4155
rect 22335 4120 22340 4150
rect 22370 4120 22375 4150
rect 22335 4115 22375 4120
rect 22445 4150 22485 4155
rect 22445 4120 22450 4150
rect 22480 4120 22485 4150
rect 22445 4115 22485 4120
rect 22645 4150 22685 4155
rect 22645 4120 22650 4150
rect 22680 4120 22685 4150
rect 22645 4115 22685 4120
rect 22810 4150 22850 4155
rect 22810 4120 22815 4150
rect 22845 4120 22850 4150
rect 22810 4115 22850 4120
rect 22975 4150 23015 4155
rect 22975 4120 22980 4150
rect 23010 4120 23015 4150
rect 22975 4115 23015 4120
rect 23195 4150 23235 4155
rect 23195 4120 23200 4150
rect 23230 4120 23235 4150
rect 23195 4115 23235 4120
rect 23325 4150 23365 4155
rect 23325 4120 23330 4150
rect 23360 4120 23365 4150
rect 23325 4115 23365 4120
rect 23585 4150 23625 4155
rect 23585 4120 23590 4150
rect 23620 4120 23625 4150
rect 23585 4115 23625 4120
rect 23925 4150 23965 4155
rect 23925 4120 23930 4150
rect 23960 4120 23965 4150
rect 23925 4115 23965 4120
rect 21565 3905 21605 3910
rect 21565 3875 21570 3905
rect 21600 3875 21605 3905
rect 21565 3870 21605 3875
rect 22525 3900 22565 3905
rect 22525 3870 22530 3900
rect 22560 3870 22565 3900
rect 22525 3865 22565 3870
rect 23040 3900 23100 3905
rect 23040 3870 23045 3900
rect 23075 3870 23100 3900
rect 23040 3865 23100 3870
rect 21850 3615 21890 3620
rect 21850 3585 21855 3615
rect 21885 3585 21890 3615
rect 21850 3580 21890 3585
rect 21625 3560 21665 3565
rect 21625 3530 21630 3560
rect 21660 3530 21665 3560
rect 21625 3525 21665 3530
rect 21995 3560 22035 3565
rect 21995 3530 22000 3560
rect 22030 3530 22035 3560
rect 21995 3525 22035 3530
rect 22075 3560 22115 3565
rect 22075 3530 22080 3560
rect 22110 3530 22115 3560
rect 22075 3525 22115 3530
rect 22445 3560 22485 3565
rect 22445 3530 22450 3560
rect 22480 3530 22485 3560
rect 22445 3525 22485 3530
rect 21565 3215 21605 3220
rect 21565 3185 21570 3215
rect 21600 3185 21605 3215
rect 22535 3205 22555 3865
rect 22615 3615 22655 3620
rect 22615 3585 22620 3615
rect 22650 3585 22655 3615
rect 22615 3580 22655 3585
rect 22570 3560 22610 3565
rect 22570 3530 22575 3560
rect 22605 3530 22610 3560
rect 22570 3525 22610 3530
rect 22625 3505 22645 3580
rect 22665 3560 22745 3565
rect 22665 3530 22670 3560
rect 22700 3530 22710 3560
rect 22740 3530 22745 3560
rect 22665 3525 22745 3530
rect 22810 3560 22850 3565
rect 22810 3530 22815 3560
rect 22845 3530 22850 3560
rect 22810 3525 22850 3530
rect 22975 3560 23015 3565
rect 22975 3530 22980 3560
rect 23010 3530 23015 3560
rect 22975 3525 23015 3530
rect 22625 3475 22630 3505
rect 22660 3475 22665 3505
rect 22625 3470 22665 3475
rect 23080 3225 23100 3865
rect 23115 3900 23155 3910
rect 23115 3880 23125 3900
rect 23145 3880 23155 3900
rect 23115 3870 23155 3880
rect 23115 3625 23135 3870
rect 23115 3620 23155 3625
rect 23115 3590 23120 3620
rect 23150 3590 23155 3620
rect 23335 3615 23355 4115
rect 23450 4095 23525 4100
rect 23450 4065 23455 4095
rect 23485 4065 23525 4095
rect 23450 4060 23525 4065
rect 23765 4095 23805 4100
rect 23765 4065 23770 4095
rect 23800 4065 23805 4095
rect 23765 4060 23805 4065
rect 24050 4095 24090 4155
rect 26545 4155 26555 4190
rect 26590 4155 26600 4190
rect 26545 4145 26600 4155
rect 24050 4065 24055 4095
rect 24085 4065 24090 4095
rect 24050 4060 24090 4065
rect 24670 4115 24710 4120
rect 24670 4085 24675 4115
rect 24705 4085 24710 4115
rect 24670 4065 24710 4085
rect 23410 3615 23450 3620
rect 23115 3585 23155 3590
rect 23325 3585 23330 3615
rect 23360 3585 23365 3615
rect 23410 3585 23415 3615
rect 23445 3585 23450 3615
rect 23505 3565 23525 4060
rect 24670 4045 24680 4065
rect 24700 4045 24710 4065
rect 24670 4005 24710 4045
rect 24670 3985 24680 4005
rect 24700 3985 24710 4005
rect 24670 3955 24710 3985
rect 24670 3935 24680 3955
rect 24700 3935 24710 3955
rect 24000 3925 24040 3930
rect 24000 3895 24005 3925
rect 24035 3895 24040 3925
rect 24000 3890 24040 3895
rect 24090 3925 24130 3930
rect 24090 3895 24095 3925
rect 24125 3895 24130 3925
rect 24090 3745 24130 3895
rect 24670 3905 24710 3935
rect 24670 3885 24680 3905
rect 24700 3885 24710 3905
rect 24670 3855 24710 3885
rect 24670 3835 24680 3855
rect 24700 3835 24710 3855
rect 24670 3825 24710 3835
rect 24780 4115 24820 4120
rect 24780 4085 24785 4115
rect 24815 4085 24820 4115
rect 24780 4005 24820 4085
rect 25000 4115 25040 4120
rect 25000 4085 25005 4115
rect 25035 4085 25040 4115
rect 24780 3985 24790 4005
rect 24810 3985 24820 4005
rect 24780 3955 24820 3985
rect 24780 3935 24790 3955
rect 24810 3935 24820 3955
rect 24780 3905 24820 3935
rect 24780 3885 24790 3905
rect 24810 3885 24820 3905
rect 24780 3855 24820 3885
rect 24780 3835 24790 3855
rect 24810 3835 24820 3855
rect 24780 3825 24820 3835
rect 24890 4005 24930 4015
rect 24890 3985 24900 4005
rect 24920 3985 24930 4005
rect 24890 3955 24930 3985
rect 24890 3935 24900 3955
rect 24920 3935 24930 3955
rect 24890 3905 24930 3935
rect 24890 3885 24900 3905
rect 24920 3885 24930 3905
rect 24890 3855 24930 3885
rect 24890 3835 24900 3855
rect 24920 3835 24930 3855
rect 24890 3825 24930 3835
rect 25000 4005 25040 4085
rect 25160 4115 25200 4120
rect 25160 4085 25165 4115
rect 25195 4085 25200 4115
rect 25160 4015 25200 4085
rect 25320 4115 25360 4120
rect 25320 4085 25325 4115
rect 25355 4085 25360 4115
rect 25000 3985 25010 4005
rect 25030 3985 25040 4005
rect 25000 3955 25040 3985
rect 25000 3935 25010 3955
rect 25030 3935 25040 3955
rect 25000 3905 25040 3935
rect 25000 3885 25010 3905
rect 25030 3885 25040 3905
rect 25000 3855 25040 3885
rect 25000 3835 25010 3855
rect 25030 3835 25040 3855
rect 25000 3825 25040 3835
rect 25110 4005 25250 4015
rect 25110 3985 25120 4005
rect 25140 3985 25170 4005
rect 25190 3985 25220 4005
rect 25240 3985 25250 4005
rect 25110 3955 25250 3985
rect 25110 3935 25120 3955
rect 25140 3935 25170 3955
rect 25190 3935 25220 3955
rect 25240 3935 25250 3955
rect 25110 3905 25250 3935
rect 25110 3885 25120 3905
rect 25140 3885 25170 3905
rect 25190 3885 25220 3905
rect 25240 3885 25250 3905
rect 25110 3855 25250 3885
rect 25110 3835 25120 3855
rect 25140 3835 25170 3855
rect 25190 3835 25220 3855
rect 25240 3835 25250 3855
rect 25110 3825 25250 3835
rect 25320 4005 25360 4085
rect 25540 4115 25580 4120
rect 25540 4085 25545 4115
rect 25575 4085 25580 4115
rect 25320 3985 25330 4005
rect 25350 3985 25360 4005
rect 25320 3955 25360 3985
rect 25320 3935 25330 3955
rect 25350 3935 25360 3955
rect 25320 3905 25360 3935
rect 25320 3885 25330 3905
rect 25350 3885 25360 3905
rect 25320 3855 25360 3885
rect 25320 3835 25330 3855
rect 25350 3835 25360 3855
rect 25320 3825 25360 3835
rect 25430 4005 25470 4015
rect 25430 3985 25440 4005
rect 25460 3985 25470 4005
rect 25430 3955 25470 3985
rect 25430 3935 25440 3955
rect 25460 3935 25470 3955
rect 25430 3905 25470 3935
rect 25430 3885 25440 3905
rect 25460 3885 25470 3905
rect 25430 3855 25470 3885
rect 25430 3835 25440 3855
rect 25460 3835 25470 3855
rect 24090 3715 24095 3745
rect 24125 3715 24130 3745
rect 24090 3710 24130 3715
rect 24890 3800 24930 3810
rect 24890 3780 24900 3800
rect 24920 3780 24930 3800
rect 24090 3690 24130 3695
rect 24090 3660 24095 3690
rect 24125 3660 24130 3690
rect 23730 3615 23770 3620
rect 23730 3585 23735 3615
rect 23765 3585 23770 3615
rect 23730 3580 23770 3585
rect 24090 3615 24130 3660
rect 24890 3690 24930 3780
rect 24890 3660 24895 3690
rect 24925 3660 24930 3690
rect 24890 3655 24930 3660
rect 24090 3585 24095 3615
rect 24125 3585 24130 3615
rect 24090 3580 24130 3585
rect 24145 3635 24185 3640
rect 24145 3605 24150 3635
rect 24180 3605 24185 3635
rect 23195 3560 23235 3565
rect 23195 3530 23200 3560
rect 23230 3530 23235 3560
rect 23195 3525 23235 3530
rect 23390 3560 23430 3565
rect 23390 3530 23395 3560
rect 23425 3530 23430 3560
rect 23390 3525 23430 3530
rect 23495 3560 23535 3565
rect 23495 3530 23500 3560
rect 23530 3530 23535 3560
rect 23495 3525 23535 3530
rect 23585 3560 23625 3565
rect 23585 3530 23590 3560
rect 23620 3530 23625 3560
rect 23585 3525 23625 3530
rect 23925 3560 23965 3565
rect 23925 3530 23930 3560
rect 23960 3530 23965 3560
rect 23925 3525 23965 3530
rect 21565 3180 21605 3185
rect 22515 3200 22555 3205
rect 22515 3170 22520 3200
rect 22550 3170 22555 3200
rect 23060 3220 23100 3225
rect 23060 3190 23065 3220
rect 23095 3190 23100 3220
rect 23845 3235 23885 3240
rect 23060 3185 23100 3190
rect 23125 3200 23165 3210
rect 22515 3165 22555 3170
rect 23125 3180 23135 3200
rect 23155 3180 23165 3200
rect 23125 3170 23165 3180
rect 23845 3205 23850 3235
rect 23880 3205 23885 3235
rect 23125 3040 23145 3170
rect 23115 3035 23155 3040
rect 21830 3025 21870 3030
rect 21830 2995 21835 3025
rect 21865 2995 21870 3025
rect 21830 2990 21870 2995
rect 22690 3025 22730 3030
rect 22690 2995 22695 3025
rect 22725 2995 22730 3025
rect 23115 3005 23120 3035
rect 23150 3005 23155 3035
rect 23115 3000 23155 3005
rect 23730 3025 23770 3030
rect 22690 2990 22730 2995
rect 23730 2995 23735 3025
rect 23765 2995 23770 3025
rect 23730 2990 23770 2995
rect 21625 2970 21665 2975
rect 21625 2940 21630 2970
rect 21660 2940 21665 2970
rect 21625 2935 21665 2940
rect 21735 2970 21775 2975
rect 21735 2940 21740 2970
rect 21770 2940 21775 2970
rect 21735 2935 21775 2940
rect 21885 2970 21925 2975
rect 21885 2940 21890 2970
rect 21920 2940 21925 2970
rect 21885 2935 21925 2940
rect 21995 2970 22035 2975
rect 21995 2940 22000 2970
rect 22030 2940 22035 2970
rect 21995 2935 22035 2940
rect 22075 2970 22115 2975
rect 22075 2940 22080 2970
rect 22110 2940 22115 2970
rect 22075 2935 22115 2940
rect 22185 2970 22225 2975
rect 22185 2940 22190 2970
rect 22220 2940 22225 2970
rect 22185 2935 22225 2940
rect 22335 2970 22375 2975
rect 22335 2940 22340 2970
rect 22370 2940 22375 2970
rect 22335 2935 22375 2940
rect 22445 2970 22485 2975
rect 22445 2940 22450 2970
rect 22480 2940 22485 2970
rect 22445 2935 22485 2940
rect 22595 2970 22635 2975
rect 22595 2940 22600 2970
rect 22630 2940 22635 2970
rect 22595 2935 22635 2940
rect 22815 2970 22855 2975
rect 22815 2940 22820 2970
rect 22850 2940 22855 2970
rect 22815 2935 22855 2940
rect 22980 2970 23020 2975
rect 22980 2940 22985 2970
rect 23015 2940 23020 2970
rect 22980 2935 23020 2940
rect 23195 2970 23235 2975
rect 23195 2940 23200 2970
rect 23230 2940 23235 2970
rect 23195 2935 23235 2940
rect 23390 2970 23430 2975
rect 23390 2940 23395 2970
rect 23425 2940 23430 2970
rect 23390 2935 23430 2940
rect 23585 2970 23625 2975
rect 23585 2940 23590 2970
rect 23620 2940 23625 2970
rect 23585 2935 23625 2940
rect 23845 2940 23885 3205
rect 24000 3195 24040 3200
rect 24000 3165 24005 3195
rect 24035 3165 24040 3195
rect 24000 3160 24040 3165
rect 24145 3195 24185 3605
rect 24145 3165 24150 3195
rect 24180 3165 24185 3195
rect 24145 3160 24185 3165
rect 24200 3580 24240 3585
rect 24200 3550 24205 3580
rect 24235 3550 24240 3580
rect 24200 3025 24240 3550
rect 25100 3580 25140 3585
rect 25100 3550 25105 3580
rect 25135 3550 25140 3580
rect 24990 3520 25030 3525
rect 24990 3490 24995 3520
rect 25025 3490 25030 3520
rect 24770 3455 24810 3465
rect 24770 3435 24780 3455
rect 24800 3435 24810 3455
rect 24770 3405 24810 3435
rect 24770 3385 24780 3405
rect 24800 3385 24810 3405
rect 24770 3355 24810 3385
rect 24770 3335 24780 3355
rect 24800 3335 24810 3355
rect 24770 3305 24810 3335
rect 24770 3285 24780 3305
rect 24800 3285 24810 3305
rect 24770 3245 24810 3285
rect 24770 3225 24780 3245
rect 24800 3225 24810 3245
rect 24770 3195 24810 3225
rect 24770 3165 24775 3195
rect 24805 3165 24810 3195
rect 24770 3160 24810 3165
rect 24880 3455 24920 3465
rect 24880 3435 24890 3455
rect 24910 3435 24920 3455
rect 24880 3405 24920 3435
rect 24880 3385 24890 3405
rect 24910 3385 24920 3405
rect 24880 3355 24920 3385
rect 24880 3335 24890 3355
rect 24910 3335 24920 3355
rect 24880 3305 24920 3335
rect 24880 3285 24890 3305
rect 24910 3285 24920 3305
rect 24880 3195 24920 3285
rect 24990 3455 25030 3490
rect 25100 3515 25140 3550
rect 25100 3495 25110 3515
rect 25130 3495 25140 3515
rect 25100 3485 25140 3495
rect 25210 3520 25250 3525
rect 25210 3490 25215 3520
rect 25245 3490 25250 3520
rect 24990 3435 25000 3455
rect 25020 3435 25030 3455
rect 24990 3405 25030 3435
rect 24990 3385 25000 3405
rect 25020 3385 25030 3405
rect 24990 3355 25030 3385
rect 24990 3335 25000 3355
rect 25020 3335 25030 3355
rect 24990 3305 25030 3335
rect 24990 3285 25000 3305
rect 25020 3285 25030 3305
rect 24990 3275 25030 3285
rect 25100 3455 25140 3465
rect 25100 3435 25110 3455
rect 25130 3435 25140 3455
rect 25100 3405 25140 3435
rect 25100 3385 25110 3405
rect 25130 3385 25140 3405
rect 25100 3355 25140 3385
rect 25100 3335 25110 3355
rect 25130 3335 25140 3355
rect 25100 3305 25140 3335
rect 25100 3285 25110 3305
rect 25130 3285 25140 3305
rect 24880 3165 24885 3195
rect 24915 3165 24920 3195
rect 24880 3160 24920 3165
rect 25100 3195 25140 3285
rect 25210 3455 25250 3490
rect 25430 3520 25470 3835
rect 25540 4005 25580 4085
rect 25700 4115 25740 4120
rect 25700 4085 25705 4115
rect 25735 4085 25740 4115
rect 25700 4015 25740 4085
rect 25860 4115 25900 4120
rect 25860 4085 25865 4115
rect 25895 4085 25900 4115
rect 25540 3985 25550 4005
rect 25570 3985 25580 4005
rect 25540 3955 25580 3985
rect 25540 3935 25550 3955
rect 25570 3935 25580 3955
rect 25540 3905 25580 3935
rect 25540 3885 25550 3905
rect 25570 3885 25580 3905
rect 25540 3855 25580 3885
rect 25540 3835 25550 3855
rect 25570 3835 25580 3855
rect 25540 3825 25580 3835
rect 25650 4005 25790 4015
rect 25650 3985 25660 4005
rect 25680 3985 25710 4005
rect 25730 3985 25760 4005
rect 25780 3985 25790 4005
rect 25650 3955 25790 3985
rect 25650 3935 25660 3955
rect 25680 3935 25710 3955
rect 25730 3935 25760 3955
rect 25780 3935 25790 3955
rect 25650 3905 25790 3935
rect 25650 3885 25660 3905
rect 25680 3885 25710 3905
rect 25730 3885 25760 3905
rect 25780 3885 25790 3905
rect 25650 3855 25790 3885
rect 25650 3835 25660 3855
rect 25680 3835 25710 3855
rect 25730 3835 25760 3855
rect 25780 3835 25790 3855
rect 25650 3825 25790 3835
rect 25860 4005 25900 4085
rect 26080 4115 26120 4120
rect 26080 4085 26085 4115
rect 26115 4085 26120 4115
rect 25860 3985 25870 4005
rect 25890 3985 25900 4005
rect 25860 3955 25900 3985
rect 25860 3935 25870 3955
rect 25890 3935 25900 3955
rect 25860 3905 25900 3935
rect 25860 3885 25870 3905
rect 25890 3885 25900 3905
rect 25860 3855 25900 3885
rect 25860 3835 25870 3855
rect 25890 3835 25900 3855
rect 25860 3825 25900 3835
rect 25970 4005 26010 4015
rect 25970 3985 25980 4005
rect 26000 3985 26010 4005
rect 25970 3955 26010 3985
rect 25970 3935 25980 3955
rect 26000 3935 26010 3955
rect 25970 3905 26010 3935
rect 25970 3885 25980 3905
rect 26000 3885 26010 3905
rect 25970 3855 26010 3885
rect 25970 3835 25980 3855
rect 26000 3835 26010 3855
rect 25905 3785 25945 3790
rect 25905 3755 25910 3785
rect 25940 3755 25945 3785
rect 25905 3750 25945 3755
rect 25970 3660 26010 3835
rect 26080 4005 26120 4085
rect 26080 3985 26090 4005
rect 26110 3985 26120 4005
rect 26080 3955 26120 3985
rect 26080 3935 26090 3955
rect 26110 3935 26120 3955
rect 26080 3905 26120 3935
rect 26080 3885 26090 3905
rect 26110 3885 26120 3905
rect 26080 3855 26120 3885
rect 26080 3835 26090 3855
rect 26110 3835 26120 3855
rect 26080 3825 26120 3835
rect 26190 4115 26230 4120
rect 26190 4085 26195 4115
rect 26225 4085 26230 4115
rect 26190 4065 26230 4085
rect 26190 4045 26200 4065
rect 26220 4045 26230 4065
rect 26190 4005 26230 4045
rect 26190 3985 26200 4005
rect 26220 3985 26230 4005
rect 26190 3955 26230 3985
rect 26190 3935 26200 3955
rect 26220 3935 26230 3955
rect 26190 3905 26230 3935
rect 26190 3885 26200 3905
rect 26220 3885 26230 3905
rect 26190 3855 26230 3885
rect 26190 3835 26200 3855
rect 26220 3835 26230 3855
rect 26190 3825 26230 3835
rect 26370 3795 26425 3805
rect 26035 3785 26075 3790
rect 26035 3755 26040 3785
rect 26070 3755 26075 3785
rect 26035 3750 26075 3755
rect 26370 3760 26380 3795
rect 26415 3760 26425 3795
rect 26370 3750 26425 3760
rect 25430 3490 25435 3520
rect 25465 3490 25470 3520
rect 25685 3635 25725 3640
rect 25685 3605 25690 3635
rect 25720 3605 25725 3635
rect 25685 3535 25725 3605
rect 25685 3505 25690 3535
rect 25720 3505 25725 3535
rect 25970 3630 25975 3660
rect 26005 3630 26010 3660
rect 25685 3500 25725 3505
rect 25750 3520 25790 3525
rect 25430 3485 25470 3490
rect 25750 3490 25755 3520
rect 25785 3490 25790 3520
rect 25210 3435 25220 3455
rect 25240 3435 25250 3455
rect 25210 3405 25250 3435
rect 25210 3385 25220 3405
rect 25240 3385 25250 3405
rect 25210 3355 25250 3385
rect 25210 3335 25220 3355
rect 25240 3335 25250 3355
rect 25210 3305 25250 3335
rect 25210 3285 25220 3305
rect 25240 3285 25250 3305
rect 25210 3275 25250 3285
rect 25320 3455 25360 3465
rect 25320 3435 25330 3455
rect 25350 3435 25360 3455
rect 25320 3405 25360 3435
rect 25320 3385 25330 3405
rect 25350 3385 25360 3405
rect 25320 3355 25360 3385
rect 25320 3335 25330 3355
rect 25350 3335 25360 3355
rect 25320 3305 25360 3335
rect 25320 3285 25330 3305
rect 25350 3285 25360 3305
rect 25100 3165 25105 3195
rect 25135 3165 25140 3195
rect 25100 3160 25140 3165
rect 25320 3195 25360 3285
rect 25430 3455 25570 3465
rect 25430 3435 25440 3455
rect 25460 3435 25490 3455
rect 25510 3435 25540 3455
rect 25560 3435 25570 3455
rect 25430 3405 25570 3435
rect 25430 3385 25440 3405
rect 25460 3385 25490 3405
rect 25510 3385 25540 3405
rect 25560 3385 25570 3405
rect 25430 3355 25570 3385
rect 25430 3335 25440 3355
rect 25460 3335 25490 3355
rect 25510 3335 25540 3355
rect 25560 3335 25570 3355
rect 25430 3305 25570 3335
rect 25430 3285 25440 3305
rect 25460 3285 25490 3305
rect 25510 3285 25540 3305
rect 25560 3285 25570 3305
rect 25430 3275 25570 3285
rect 25640 3455 25680 3465
rect 25640 3435 25650 3455
rect 25670 3435 25680 3455
rect 25640 3405 25680 3435
rect 25640 3385 25650 3405
rect 25670 3385 25680 3405
rect 25640 3355 25680 3385
rect 25640 3335 25650 3355
rect 25670 3335 25680 3355
rect 25640 3305 25680 3335
rect 25640 3285 25650 3305
rect 25670 3285 25680 3305
rect 25320 3165 25325 3195
rect 25355 3165 25360 3195
rect 25320 3160 25360 3165
rect 25480 3195 25520 3275
rect 25480 3165 25485 3195
rect 25515 3165 25520 3195
rect 25480 3160 25520 3165
rect 25640 3195 25680 3285
rect 25750 3455 25790 3490
rect 25970 3520 26010 3630
rect 25970 3490 25975 3520
rect 26005 3490 26010 3520
rect 26035 3535 26075 3540
rect 26035 3505 26040 3535
rect 26070 3505 26075 3535
rect 26035 3500 26075 3505
rect 26370 3530 26425 3540
rect 25750 3435 25760 3455
rect 25780 3435 25790 3455
rect 25750 3405 25790 3435
rect 25750 3385 25760 3405
rect 25780 3385 25790 3405
rect 25750 3355 25790 3385
rect 25750 3335 25760 3355
rect 25780 3335 25790 3355
rect 25750 3305 25790 3335
rect 25750 3285 25760 3305
rect 25780 3285 25790 3305
rect 25750 3275 25790 3285
rect 25860 3455 25900 3465
rect 25860 3435 25870 3455
rect 25890 3435 25900 3455
rect 25860 3405 25900 3435
rect 25860 3385 25870 3405
rect 25890 3385 25900 3405
rect 25860 3355 25900 3385
rect 25860 3335 25870 3355
rect 25890 3335 25900 3355
rect 25860 3305 25900 3335
rect 25860 3285 25870 3305
rect 25890 3285 25900 3305
rect 25640 3165 25645 3195
rect 25675 3165 25680 3195
rect 25640 3160 25680 3165
rect 25860 3195 25900 3285
rect 25970 3455 26010 3490
rect 26370 3495 26380 3530
rect 26415 3495 26425 3530
rect 26370 3485 26425 3495
rect 25970 3435 25980 3455
rect 26000 3435 26010 3455
rect 25970 3405 26010 3435
rect 25970 3385 25980 3405
rect 26000 3385 26010 3405
rect 25970 3355 26010 3385
rect 25970 3335 25980 3355
rect 26000 3335 26010 3355
rect 25970 3305 26010 3335
rect 25970 3285 25980 3305
rect 26000 3285 26010 3305
rect 25970 3275 26010 3285
rect 26080 3455 26120 3465
rect 26080 3435 26090 3455
rect 26110 3435 26120 3455
rect 26080 3405 26120 3435
rect 26080 3385 26090 3405
rect 26110 3385 26120 3405
rect 26080 3355 26120 3385
rect 26080 3335 26090 3355
rect 26110 3335 26120 3355
rect 26080 3305 26120 3335
rect 26080 3285 26090 3305
rect 26110 3285 26120 3305
rect 25860 3165 25865 3195
rect 25895 3165 25900 3195
rect 25860 3160 25900 3165
rect 26080 3195 26120 3285
rect 26080 3165 26085 3195
rect 26115 3165 26120 3195
rect 26080 3160 26120 3165
rect 26190 3455 26230 3465
rect 26190 3435 26200 3455
rect 26220 3435 26230 3455
rect 26190 3405 26230 3435
rect 26190 3385 26200 3405
rect 26220 3385 26230 3405
rect 26190 3355 26230 3385
rect 26190 3335 26200 3355
rect 26220 3335 26230 3355
rect 26190 3305 26230 3335
rect 26190 3285 26200 3305
rect 26220 3285 26230 3305
rect 26190 3245 26230 3285
rect 26190 3225 26200 3245
rect 26220 3225 26230 3245
rect 26190 3195 26230 3225
rect 26190 3165 26195 3195
rect 26225 3165 26230 3195
rect 26190 3160 26230 3165
rect 24200 2995 24205 3025
rect 24235 2995 24240 3025
rect 24200 2990 24240 2995
rect 23845 2910 23850 2940
rect 23880 2910 23885 2940
rect 23845 2905 23885 2910
rect 26490 2940 26545 2950
rect 26490 2905 26500 2940
rect 26535 2905 26545 2940
rect 26490 2895 26545 2905
<< via1 >>
rect 24055 4155 24085 4185
rect 21630 4145 21660 4150
rect 21630 4125 21635 4145
rect 21635 4125 21655 4145
rect 21655 4125 21660 4145
rect 21630 4120 21660 4125
rect 21740 4145 21770 4150
rect 21740 4125 21745 4145
rect 21745 4125 21765 4145
rect 21765 4125 21770 4145
rect 21740 4120 21770 4125
rect 21890 4145 21920 4150
rect 21890 4125 21895 4145
rect 21895 4125 21915 4145
rect 21915 4125 21920 4145
rect 21890 4120 21920 4125
rect 22005 4145 22035 4150
rect 22005 4125 22010 4145
rect 22010 4125 22030 4145
rect 22030 4125 22035 4145
rect 22005 4120 22035 4125
rect 22080 4145 22110 4150
rect 22080 4125 22085 4145
rect 22085 4125 22105 4145
rect 22105 4125 22110 4145
rect 22080 4120 22110 4125
rect 22190 4145 22220 4150
rect 22190 4125 22195 4145
rect 22195 4125 22215 4145
rect 22215 4125 22220 4145
rect 22190 4120 22220 4125
rect 22340 4145 22370 4150
rect 22340 4125 22345 4145
rect 22345 4125 22365 4145
rect 22365 4125 22370 4145
rect 22340 4120 22370 4125
rect 22450 4145 22480 4150
rect 22450 4125 22455 4145
rect 22455 4125 22475 4145
rect 22475 4125 22480 4145
rect 22450 4120 22480 4125
rect 22650 4145 22680 4150
rect 22650 4125 22655 4145
rect 22655 4125 22675 4145
rect 22675 4125 22680 4145
rect 22650 4120 22680 4125
rect 22815 4145 22845 4150
rect 22815 4125 22820 4145
rect 22820 4125 22840 4145
rect 22840 4125 22845 4145
rect 22815 4120 22845 4125
rect 22980 4145 23010 4150
rect 22980 4125 22985 4145
rect 22985 4125 23005 4145
rect 23005 4125 23010 4145
rect 22980 4120 23010 4125
rect 23200 4145 23230 4150
rect 23200 4125 23205 4145
rect 23205 4125 23225 4145
rect 23225 4125 23230 4145
rect 23200 4120 23230 4125
rect 23330 4120 23360 4150
rect 23590 4145 23620 4150
rect 23590 4125 23595 4145
rect 23595 4125 23615 4145
rect 23615 4125 23620 4145
rect 23590 4120 23620 4125
rect 23930 4145 23960 4150
rect 23930 4125 23935 4145
rect 23935 4125 23955 4145
rect 23955 4125 23960 4145
rect 23930 4120 23960 4125
rect 21570 3900 21600 3905
rect 21570 3880 21575 3900
rect 21575 3880 21595 3900
rect 21595 3880 21600 3900
rect 21570 3875 21600 3880
rect 22530 3895 22560 3900
rect 22530 3875 22535 3895
rect 22535 3875 22555 3895
rect 22555 3875 22560 3895
rect 22530 3870 22560 3875
rect 23045 3895 23075 3900
rect 23045 3875 23050 3895
rect 23050 3875 23070 3895
rect 23070 3875 23075 3895
rect 23045 3870 23075 3875
rect 21855 3610 21885 3615
rect 21855 3590 21860 3610
rect 21860 3590 21880 3610
rect 21880 3590 21885 3610
rect 21855 3585 21885 3590
rect 21630 3555 21660 3560
rect 21630 3535 21635 3555
rect 21635 3535 21655 3555
rect 21655 3535 21660 3555
rect 21630 3530 21660 3535
rect 22000 3555 22030 3560
rect 22000 3535 22005 3555
rect 22005 3535 22025 3555
rect 22025 3535 22030 3555
rect 22000 3530 22030 3535
rect 22080 3555 22110 3560
rect 22080 3535 22085 3555
rect 22085 3535 22105 3555
rect 22105 3535 22110 3555
rect 22080 3530 22110 3535
rect 22450 3555 22480 3560
rect 22450 3535 22455 3555
rect 22455 3535 22475 3555
rect 22475 3535 22480 3555
rect 22450 3530 22480 3535
rect 21570 3210 21600 3215
rect 21570 3190 21575 3210
rect 21575 3190 21595 3210
rect 21595 3190 21600 3210
rect 21570 3185 21600 3190
rect 22620 3585 22650 3615
rect 22575 3555 22605 3560
rect 22575 3535 22580 3555
rect 22580 3535 22600 3555
rect 22600 3535 22605 3555
rect 22575 3530 22605 3535
rect 22670 3555 22700 3560
rect 22670 3535 22675 3555
rect 22675 3535 22695 3555
rect 22695 3535 22700 3555
rect 22670 3530 22700 3535
rect 22710 3555 22740 3560
rect 22710 3535 22715 3555
rect 22715 3535 22735 3555
rect 22735 3535 22740 3555
rect 22710 3530 22740 3535
rect 22815 3555 22845 3560
rect 22815 3535 22820 3555
rect 22820 3535 22840 3555
rect 22840 3535 22845 3555
rect 22815 3530 22845 3535
rect 22980 3555 23010 3560
rect 22980 3535 22985 3555
rect 22985 3535 23005 3555
rect 23005 3535 23010 3555
rect 22980 3530 23010 3535
rect 22630 3500 22660 3505
rect 22630 3480 22635 3500
rect 22635 3480 22655 3500
rect 22655 3480 22660 3500
rect 22630 3475 22660 3480
rect 23120 3590 23150 3620
rect 23455 4090 23485 4095
rect 23455 4070 23460 4090
rect 23460 4070 23480 4090
rect 23480 4070 23485 4090
rect 23455 4065 23485 4070
rect 23770 4090 23800 4095
rect 23770 4070 23775 4090
rect 23775 4070 23795 4090
rect 23795 4070 23800 4090
rect 23770 4065 23800 4070
rect 26555 4155 26590 4190
rect 24055 4065 24085 4095
rect 24675 4085 24705 4115
rect 23330 3585 23360 3615
rect 23415 3610 23445 3615
rect 23415 3590 23420 3610
rect 23420 3590 23440 3610
rect 23440 3590 23445 3610
rect 23415 3585 23445 3590
rect 24005 3920 24035 3925
rect 24005 3900 24010 3920
rect 24010 3900 24030 3920
rect 24030 3900 24035 3920
rect 24005 3895 24035 3900
rect 24095 3895 24125 3925
rect 24785 4085 24815 4115
rect 25005 4085 25035 4115
rect 25165 4085 25195 4115
rect 25325 4085 25355 4115
rect 25545 4085 25575 4115
rect 24095 3715 24125 3745
rect 24095 3660 24125 3690
rect 23735 3610 23765 3615
rect 23735 3590 23740 3610
rect 23740 3590 23760 3610
rect 23760 3590 23765 3610
rect 23735 3585 23765 3590
rect 24895 3660 24925 3690
rect 24095 3585 24125 3615
rect 24150 3605 24180 3635
rect 23200 3555 23230 3560
rect 23200 3535 23205 3555
rect 23205 3535 23225 3555
rect 23225 3535 23230 3555
rect 23200 3530 23230 3535
rect 23395 3555 23425 3560
rect 23395 3535 23400 3555
rect 23400 3535 23420 3555
rect 23420 3535 23425 3555
rect 23395 3530 23425 3535
rect 23500 3530 23530 3560
rect 23590 3555 23620 3560
rect 23590 3535 23595 3555
rect 23595 3535 23615 3555
rect 23615 3535 23620 3555
rect 23590 3530 23620 3535
rect 23930 3555 23960 3560
rect 23930 3535 23935 3555
rect 23935 3535 23955 3555
rect 23955 3535 23960 3555
rect 23930 3530 23960 3535
rect 22520 3195 22550 3200
rect 22520 3175 22525 3195
rect 22525 3175 22545 3195
rect 22545 3175 22550 3195
rect 22520 3170 22550 3175
rect 23065 3215 23095 3220
rect 23065 3195 23070 3215
rect 23070 3195 23090 3215
rect 23090 3195 23095 3215
rect 23065 3190 23095 3195
rect 23850 3230 23880 3235
rect 23850 3210 23855 3230
rect 23855 3210 23875 3230
rect 23875 3210 23880 3230
rect 23850 3205 23880 3210
rect 21835 3020 21865 3025
rect 21835 3000 21840 3020
rect 21840 3000 21860 3020
rect 21860 3000 21865 3020
rect 21835 2995 21865 3000
rect 22695 3020 22725 3025
rect 22695 3000 22700 3020
rect 22700 3000 22720 3020
rect 22720 3000 22725 3020
rect 22695 2995 22725 3000
rect 23120 3005 23150 3035
rect 23735 3020 23765 3025
rect 23735 3000 23740 3020
rect 23740 3000 23760 3020
rect 23760 3000 23765 3020
rect 23735 2995 23765 3000
rect 21630 2965 21660 2970
rect 21630 2945 21635 2965
rect 21635 2945 21655 2965
rect 21655 2945 21660 2965
rect 21630 2940 21660 2945
rect 21740 2965 21770 2970
rect 21740 2945 21745 2965
rect 21745 2945 21765 2965
rect 21765 2945 21770 2965
rect 21740 2940 21770 2945
rect 21890 2965 21920 2970
rect 21890 2945 21895 2965
rect 21895 2945 21915 2965
rect 21915 2945 21920 2965
rect 21890 2940 21920 2945
rect 22000 2965 22030 2970
rect 22000 2945 22005 2965
rect 22005 2945 22025 2965
rect 22025 2945 22030 2965
rect 22000 2940 22030 2945
rect 22080 2965 22110 2970
rect 22080 2945 22085 2965
rect 22085 2945 22105 2965
rect 22105 2945 22110 2965
rect 22080 2940 22110 2945
rect 22190 2965 22220 2970
rect 22190 2945 22195 2965
rect 22195 2945 22215 2965
rect 22215 2945 22220 2965
rect 22190 2940 22220 2945
rect 22340 2965 22370 2970
rect 22340 2945 22345 2965
rect 22345 2945 22365 2965
rect 22365 2945 22370 2965
rect 22340 2940 22370 2945
rect 22450 2965 22480 2970
rect 22450 2945 22455 2965
rect 22455 2945 22475 2965
rect 22475 2945 22480 2965
rect 22450 2940 22480 2945
rect 22600 2965 22630 2970
rect 22600 2945 22605 2965
rect 22605 2945 22625 2965
rect 22625 2945 22630 2965
rect 22600 2940 22630 2945
rect 22820 2965 22850 2970
rect 22820 2945 22825 2965
rect 22825 2945 22845 2965
rect 22845 2945 22850 2965
rect 22820 2940 22850 2945
rect 22985 2965 23015 2970
rect 22985 2945 22990 2965
rect 22990 2945 23010 2965
rect 23010 2945 23015 2965
rect 22985 2940 23015 2945
rect 23200 2965 23230 2970
rect 23200 2945 23205 2965
rect 23205 2945 23225 2965
rect 23225 2945 23230 2965
rect 23200 2940 23230 2945
rect 23395 2965 23425 2970
rect 23395 2945 23400 2965
rect 23400 2945 23420 2965
rect 23420 2945 23425 2965
rect 23395 2940 23425 2945
rect 23590 2965 23620 2970
rect 23590 2945 23595 2965
rect 23595 2945 23615 2965
rect 23615 2945 23620 2965
rect 23590 2940 23620 2945
rect 24005 3190 24035 3195
rect 24005 3170 24010 3190
rect 24010 3170 24030 3190
rect 24030 3170 24035 3190
rect 24005 3165 24035 3170
rect 24150 3165 24180 3195
rect 24205 3550 24235 3580
rect 25105 3550 25135 3580
rect 24995 3490 25025 3520
rect 24775 3165 24805 3195
rect 25215 3490 25245 3520
rect 24885 3165 24915 3195
rect 25705 4085 25735 4115
rect 25865 4085 25895 4115
rect 26085 4085 26115 4115
rect 25910 3780 25940 3785
rect 25910 3760 25915 3780
rect 25915 3760 25935 3780
rect 25935 3760 25940 3780
rect 25910 3755 25940 3760
rect 26195 4085 26225 4115
rect 26040 3780 26070 3785
rect 26040 3760 26045 3780
rect 26045 3760 26065 3780
rect 26065 3760 26070 3780
rect 26040 3755 26070 3760
rect 26380 3760 26415 3795
rect 25435 3490 25465 3520
rect 25690 3605 25720 3635
rect 25690 3530 25720 3535
rect 25690 3510 25695 3530
rect 25695 3510 25715 3530
rect 25715 3510 25720 3530
rect 25690 3505 25720 3510
rect 25975 3630 26005 3660
rect 25755 3490 25785 3520
rect 25105 3165 25135 3195
rect 25325 3165 25355 3195
rect 25485 3165 25515 3195
rect 25975 3490 26005 3520
rect 26040 3530 26070 3535
rect 26040 3510 26045 3530
rect 26045 3510 26065 3530
rect 26065 3510 26070 3530
rect 26040 3505 26070 3510
rect 25645 3165 25675 3195
rect 26380 3495 26415 3530
rect 25865 3165 25895 3195
rect 26085 3165 26115 3195
rect 26195 3165 26225 3195
rect 24205 2995 24235 3025
rect 23850 2910 23880 2940
rect 26500 2905 26535 2940
<< metal2 >>
rect 26545 4190 26600 4200
rect 24050 4185 26555 4190
rect 24050 4155 24055 4185
rect 24085 4155 26555 4185
rect 26590 4155 26600 4190
rect 21505 4150 23965 4155
rect 24050 4150 26600 4155
rect 21505 4120 21630 4150
rect 21660 4120 21740 4150
rect 21770 4120 21890 4150
rect 21920 4120 22005 4150
rect 22035 4120 22080 4150
rect 22110 4120 22190 4150
rect 22220 4120 22340 4150
rect 22370 4120 22450 4150
rect 22480 4120 22650 4150
rect 22680 4120 22815 4150
rect 22845 4120 22980 4150
rect 23010 4120 23200 4150
rect 23230 4120 23330 4150
rect 23360 4120 23590 4150
rect 23620 4120 23930 4150
rect 23960 4120 23965 4150
rect 26545 4145 26600 4150
rect 21505 4115 23965 4120
rect 24670 4115 26230 4120
rect 23450 4095 23490 4100
rect 23450 4065 23455 4095
rect 23485 4065 23490 4095
rect 23450 4060 23490 4065
rect 23765 4095 24090 4100
rect 23765 4065 23770 4095
rect 23800 4065 24055 4095
rect 24085 4065 24090 4095
rect 24670 4085 24675 4115
rect 24705 4085 24785 4115
rect 24815 4085 25005 4115
rect 25035 4085 25165 4115
rect 25195 4085 25325 4115
rect 25355 4085 25545 4115
rect 25575 4085 25705 4115
rect 25735 4085 25865 4115
rect 25895 4085 26085 4115
rect 26115 4085 26195 4115
rect 26225 4085 26230 4115
rect 24670 4080 26230 4085
rect 23765 4060 24090 4065
rect 24000 3925 24130 3930
rect 21505 3905 21605 3910
rect 21505 3875 21570 3905
rect 21600 3875 21605 3905
rect 21505 3870 21605 3875
rect 22525 3900 22565 3905
rect 22525 3870 22530 3900
rect 22560 3870 22565 3900
rect 22525 3865 22565 3870
rect 23040 3900 23080 3905
rect 23040 3870 23045 3900
rect 23075 3870 23080 3900
rect 24000 3895 24005 3925
rect 24035 3895 24095 3925
rect 24125 3895 24130 3925
rect 24000 3890 24130 3895
rect 23040 3865 23080 3870
rect 26370 3795 26425 3805
rect 26370 3790 26380 3795
rect 25905 3785 25945 3790
rect 25905 3755 25910 3785
rect 25940 3755 25945 3785
rect 25905 3750 25945 3755
rect 26035 3785 26380 3790
rect 26035 3755 26040 3785
rect 26070 3760 26380 3785
rect 26415 3760 26425 3795
rect 26070 3755 26425 3760
rect 26035 3750 26425 3755
rect 24090 3745 25945 3750
rect 24090 3715 24095 3745
rect 24125 3715 25945 3745
rect 24090 3710 25945 3715
rect 24090 3690 24930 3695
rect 24090 3660 24095 3690
rect 24125 3660 24895 3690
rect 24925 3660 24930 3690
rect 24090 3655 24930 3660
rect 25970 3660 27095 3665
rect 24145 3635 25725 3640
rect 23115 3620 23155 3625
rect 21850 3615 21890 3620
rect 21850 3585 21855 3615
rect 21885 3610 21890 3615
rect 22615 3615 22655 3620
rect 23115 3615 23120 3620
rect 22615 3610 22620 3615
rect 21885 3590 22620 3610
rect 21885 3585 21890 3590
rect 21850 3580 21890 3585
rect 22615 3585 22620 3590
rect 22650 3595 23120 3615
rect 22650 3585 22655 3595
rect 23115 3590 23120 3595
rect 23150 3590 23155 3620
rect 23410 3615 23450 3620
rect 23115 3585 23155 3590
rect 23325 3585 23330 3615
rect 23360 3610 23365 3615
rect 23410 3610 23415 3615
rect 23360 3590 23415 3610
rect 23360 3585 23365 3590
rect 23410 3585 23415 3590
rect 23445 3585 23450 3615
rect 23730 3615 24130 3620
rect 23730 3585 23735 3615
rect 23765 3585 24095 3615
rect 24125 3585 24130 3615
rect 24145 3605 24150 3635
rect 24180 3605 25690 3635
rect 25720 3605 25725 3635
rect 25970 3630 25975 3660
rect 26005 3630 27095 3660
rect 25970 3625 27095 3630
rect 24145 3600 25725 3605
rect 22615 3580 22655 3585
rect 23730 3580 24130 3585
rect 24200 3580 25140 3585
rect 21505 3560 23965 3565
rect 21505 3530 21630 3560
rect 21660 3530 22000 3560
rect 22030 3530 22080 3560
rect 22110 3530 22450 3560
rect 22480 3530 22575 3560
rect 22605 3530 22670 3560
rect 22700 3530 22710 3560
rect 22740 3530 22815 3560
rect 22845 3530 22980 3560
rect 23010 3530 23200 3560
rect 23230 3530 23395 3560
rect 23425 3530 23500 3560
rect 23530 3530 23590 3560
rect 23620 3530 23930 3560
rect 23960 3530 23965 3560
rect 24200 3550 24205 3580
rect 24235 3550 25105 3580
rect 25135 3550 25140 3580
rect 24200 3545 25140 3550
rect 21505 3525 23965 3530
rect 25685 3535 25725 3540
rect 24990 3520 25470 3525
rect 22625 3475 22630 3505
rect 22660 3475 22665 3505
rect 24990 3490 24995 3520
rect 25025 3490 25215 3520
rect 25245 3490 25435 3520
rect 25465 3490 25470 3520
rect 25685 3505 25690 3535
rect 25720 3505 25725 3535
rect 26035 3535 26425 3540
rect 25685 3500 25725 3505
rect 25750 3520 26010 3525
rect 24990 3485 25470 3490
rect 25750 3490 25755 3520
rect 25785 3490 25975 3520
rect 26005 3490 26010 3520
rect 26035 3505 26040 3535
rect 26070 3530 26425 3535
rect 26070 3505 26380 3530
rect 26035 3500 26380 3505
rect 25750 3485 26010 3490
rect 26370 3495 26380 3500
rect 26415 3495 26425 3530
rect 26370 3485 26425 3495
rect 22625 3470 22665 3475
rect 23845 3235 23885 3240
rect 23060 3220 23100 3225
rect 21505 3215 21605 3220
rect 21505 3185 21570 3215
rect 21600 3185 21605 3215
rect 21505 3180 21605 3185
rect 22515 3200 22555 3205
rect 22515 3170 22520 3200
rect 22550 3170 22555 3200
rect 23060 3190 23065 3220
rect 23095 3190 23100 3220
rect 23845 3205 23850 3235
rect 23880 3205 23885 3235
rect 23845 3200 23885 3205
rect 23060 3185 23100 3190
rect 24000 3195 24185 3200
rect 22515 3165 22555 3170
rect 24000 3165 24005 3195
rect 24035 3165 24150 3195
rect 24180 3165 24185 3195
rect 24000 3160 24185 3165
rect 24770 3195 26230 3200
rect 24770 3165 24775 3195
rect 24805 3165 24885 3195
rect 24915 3165 25105 3195
rect 25135 3165 25325 3195
rect 25355 3165 25485 3195
rect 25515 3165 25645 3195
rect 25675 3165 25865 3195
rect 25895 3165 26085 3195
rect 26115 3165 26195 3195
rect 26225 3165 26230 3195
rect 24770 3160 26230 3165
rect 23115 3035 23155 3040
rect 23115 3030 23120 3035
rect 21830 3025 23120 3030
rect 21830 2995 21835 3025
rect 21865 3010 22695 3025
rect 21865 2995 21870 3010
rect 21830 2990 21870 2995
rect 22690 2995 22695 3010
rect 22725 3010 23120 3025
rect 22725 2995 22730 3010
rect 23115 3005 23120 3010
rect 23150 3005 23155 3035
rect 23115 3000 23155 3005
rect 23730 3025 24240 3030
rect 22690 2990 22730 2995
rect 23730 2995 23735 3025
rect 23765 2995 24205 3025
rect 24235 2995 24240 3025
rect 23730 2990 24240 2995
rect 21505 2970 23625 2975
rect 21505 2940 21630 2970
rect 21660 2940 21740 2970
rect 21770 2940 21890 2970
rect 21920 2940 22000 2970
rect 22030 2940 22080 2970
rect 22110 2940 22190 2970
rect 22220 2940 22340 2970
rect 22370 2940 22450 2970
rect 22480 2940 22600 2970
rect 22630 2940 22820 2970
rect 22850 2940 22985 2970
rect 23015 2940 23200 2970
rect 23230 2940 23395 2970
rect 23425 2940 23590 2970
rect 23620 2940 23625 2970
rect 26490 2945 26545 2950
rect 21505 2935 23625 2940
rect 23845 2940 26545 2945
rect 23845 2910 23850 2940
rect 23880 2910 26500 2940
rect 23845 2905 26500 2910
rect 26535 2905 26545 2940
rect 26490 2895 26545 2905
<< via2 >>
rect 26555 4155 26590 4190
rect 26380 3760 26415 3795
rect 26380 3495 26415 3530
rect 26500 2905 26535 2940
<< metal3 >>
rect 26545 4190 26600 4200
rect 26545 4155 26555 4190
rect 26590 4155 26600 4190
rect 26545 4145 26600 4155
rect 26370 3795 26425 3805
rect 26370 3760 26380 3795
rect 26415 3760 26425 3795
rect 26370 3750 26425 3760
rect 26545 3735 26845 4145
rect 26370 3530 26425 3540
rect 26370 3495 26380 3530
rect 26415 3495 26425 3530
rect 26370 3485 26425 3495
rect 26545 2950 27095 3555
rect 26490 2940 27095 2950
rect 26490 2905 26500 2940
rect 26535 2905 27095 2940
rect 26490 2895 27095 2905
<< via3 >>
rect 26380 3760 26415 3795
rect 26380 3495 26415 3530
<< mimcap >>
rect 26560 3795 26830 4130
rect 26560 3760 26570 3795
rect 26605 3760 26830 3795
rect 26560 3750 26830 3760
rect 26560 3530 27080 3540
rect 26560 3495 26570 3530
rect 26605 3495 27080 3530
rect 26560 2910 27080 3495
<< mimcapcontact >>
rect 26570 3760 26605 3795
rect 26570 3495 26605 3530
<< metal4 >>
rect 26370 3795 26615 3805
rect 26370 3760 26380 3795
rect 26415 3760 26570 3795
rect 26605 3760 26615 3795
rect 26370 3750 26615 3760
rect 26370 3530 26615 3540
rect 26370 3495 26380 3530
rect 26415 3495 26570 3530
rect 26605 3495 26615 3530
rect 26370 3485 26615 3495
<< end >>
