magic
tech sky130A
timestamp 1757103027
<< nwell >>
rect 6565 3235 9055 3855
rect 9695 3250 11305 3540
<< nmos >>
rect 6665 3945 6680 4045
rect 6720 3945 6735 4045
rect 6925 3945 6940 4045
rect 6980 3945 6995 4045
rect 7115 3945 7130 4045
rect 7170 3945 7185 4045
rect 7375 3945 7390 4045
rect 7430 3945 7445 4045
rect 7630 3945 7645 4045
rect 7795 3945 7810 4045
rect 7960 3945 7975 4045
rect 8240 3945 8255 4045
rect 8435 3945 8450 4045
rect 8630 3945 8645 4045
rect 8775 3945 8790 4045
rect 8970 3945 8985 4045
rect 9715 3820 9775 4020
rect 9825 3820 9885 4020
rect 9935 3820 9995 4020
rect 10045 3820 10105 4020
rect 10255 3820 10315 4020
rect 10365 3820 10425 4020
rect 10475 3820 10535 4020
rect 10585 3820 10645 4020
rect 10795 3820 10855 4020
rect 10905 3820 10965 4020
rect 11015 3820 11075 4020
rect 11125 3820 11185 4020
rect 6665 3045 6680 3145
rect 6720 3045 6735 3145
rect 6925 3045 6940 3145
rect 6980 3045 6995 3145
rect 7115 3045 7130 3145
rect 7170 3045 7185 3145
rect 7375 3045 7390 3145
rect 7430 3045 7445 3145
rect 7635 3045 7650 3145
rect 7690 3045 7705 3145
rect 7855 3045 7870 3145
rect 8020 3045 8035 3145
rect 8240 3045 8255 3145
rect 8435 3045 8450 3145
rect 8630 3045 8645 3145
rect 8775 3045 8790 3145
<< pmos >>
rect 6665 3635 6680 3835
rect 6720 3635 6735 3835
rect 6925 3635 6940 3835
rect 6980 3635 6995 3835
rect 7115 3635 7130 3835
rect 7170 3635 7185 3835
rect 7375 3635 7390 3835
rect 7430 3635 7445 3835
rect 7630 3635 7645 3835
rect 7795 3635 7810 3835
rect 7960 3635 7975 3835
rect 8240 3635 8255 3835
rect 8435 3635 8450 3835
rect 8630 3635 8645 3835
rect 8775 3635 8790 3835
rect 6665 3255 6680 3455
rect 6720 3255 6735 3455
rect 6925 3255 6940 3455
rect 6980 3255 6995 3455
rect 7115 3255 7130 3455
rect 7170 3255 7185 3455
rect 7375 3255 7390 3455
rect 7430 3255 7445 3455
rect 7635 3255 7650 3455
rect 7690 3255 7705 3455
rect 7855 3255 7870 3455
rect 8020 3255 8035 3455
rect 8240 3255 8255 3455
rect 8435 3255 8450 3455
rect 8630 3255 8645 3455
rect 8775 3255 8790 3455
rect 8970 3255 8985 3455
rect 9815 3270 9875 3470
rect 9925 3270 9985 3470
rect 10035 3270 10095 3470
rect 10145 3270 10205 3470
rect 10255 3270 10315 3470
rect 10365 3270 10425 3470
rect 10575 3270 10635 3470
rect 10685 3270 10745 3470
rect 10795 3270 10855 3470
rect 10905 3270 10965 3470
rect 11015 3270 11075 3470
rect 11125 3270 11185 3470
<< ndiff >>
rect 6625 4030 6665 4045
rect 6625 4010 6635 4030
rect 6655 4010 6665 4030
rect 6625 3980 6665 4010
rect 6625 3960 6635 3980
rect 6655 3960 6665 3980
rect 6625 3945 6665 3960
rect 6680 4030 6720 4045
rect 6680 4010 6690 4030
rect 6710 4010 6720 4030
rect 6680 3980 6720 4010
rect 6680 3960 6690 3980
rect 6710 3960 6720 3980
rect 6680 3945 6720 3960
rect 6735 4030 6775 4045
rect 6735 4010 6745 4030
rect 6765 4010 6775 4030
rect 6735 3980 6775 4010
rect 6735 3960 6745 3980
rect 6765 3960 6775 3980
rect 6735 3945 6775 3960
rect 6885 4030 6925 4045
rect 6885 4010 6895 4030
rect 6915 4010 6925 4030
rect 6885 3980 6925 4010
rect 6885 3960 6895 3980
rect 6915 3960 6925 3980
rect 6885 3945 6925 3960
rect 6940 4030 6980 4045
rect 6940 4010 6950 4030
rect 6970 4010 6980 4030
rect 6940 3980 6980 4010
rect 6940 3960 6950 3980
rect 6970 3960 6980 3980
rect 6940 3945 6980 3960
rect 6995 4030 7035 4045
rect 7075 4030 7115 4045
rect 6995 4010 7005 4030
rect 7025 4010 7035 4030
rect 7075 4010 7085 4030
rect 7105 4010 7115 4030
rect 6995 3980 7035 4010
rect 7075 3980 7115 4010
rect 6995 3960 7005 3980
rect 7025 3960 7035 3980
rect 7075 3960 7085 3980
rect 7105 3960 7115 3980
rect 6995 3945 7035 3960
rect 7075 3945 7115 3960
rect 7130 4030 7170 4045
rect 7130 4010 7140 4030
rect 7160 4010 7170 4030
rect 7130 3980 7170 4010
rect 7130 3960 7140 3980
rect 7160 3960 7170 3980
rect 7130 3945 7170 3960
rect 7185 4030 7225 4045
rect 7185 4010 7195 4030
rect 7215 4010 7225 4030
rect 7185 3980 7225 4010
rect 7185 3960 7195 3980
rect 7215 3960 7225 3980
rect 7185 3945 7225 3960
rect 7335 4030 7375 4045
rect 7335 4010 7345 4030
rect 7365 4010 7375 4030
rect 7335 3980 7375 4010
rect 7335 3960 7345 3980
rect 7365 3960 7375 3980
rect 7335 3945 7375 3960
rect 7390 4030 7430 4045
rect 7390 4010 7400 4030
rect 7420 4010 7430 4030
rect 7390 3980 7430 4010
rect 7390 3960 7400 3980
rect 7420 3960 7430 3980
rect 7390 3945 7430 3960
rect 7445 4030 7485 4045
rect 7445 4010 7455 4030
rect 7475 4010 7485 4030
rect 7445 3980 7485 4010
rect 7445 3960 7455 3980
rect 7475 3960 7485 3980
rect 7445 3945 7485 3960
rect 7590 4030 7630 4045
rect 7590 4010 7600 4030
rect 7620 4010 7630 4030
rect 7590 3980 7630 4010
rect 7590 3960 7600 3980
rect 7620 3960 7630 3980
rect 7590 3945 7630 3960
rect 7645 4030 7685 4045
rect 7645 4010 7655 4030
rect 7675 4010 7685 4030
rect 7645 3980 7685 4010
rect 7645 3960 7655 3980
rect 7675 3960 7685 3980
rect 7645 3945 7685 3960
rect 7755 4030 7795 4045
rect 7755 4010 7765 4030
rect 7785 4010 7795 4030
rect 7755 3980 7795 4010
rect 7755 3960 7765 3980
rect 7785 3960 7795 3980
rect 7755 3945 7795 3960
rect 7810 4030 7850 4045
rect 7810 4010 7820 4030
rect 7840 4010 7850 4030
rect 7810 3980 7850 4010
rect 7810 3960 7820 3980
rect 7840 3960 7850 3980
rect 7810 3945 7850 3960
rect 7920 4030 7960 4045
rect 7920 4010 7930 4030
rect 7950 4010 7960 4030
rect 7920 3980 7960 4010
rect 7920 3960 7930 3980
rect 7950 3960 7960 3980
rect 7920 3945 7960 3960
rect 7975 4030 8015 4045
rect 7975 4010 7985 4030
rect 8005 4010 8015 4030
rect 7975 3980 8015 4010
rect 7975 3960 7985 3980
rect 8005 3960 8015 3980
rect 7975 3945 8015 3960
rect 8190 4030 8240 4045
rect 8190 4010 8205 4030
rect 8225 4010 8240 4030
rect 8190 3980 8240 4010
rect 8190 3960 8205 3980
rect 8225 3960 8240 3980
rect 8190 3945 8240 3960
rect 8255 4030 8305 4045
rect 8255 4010 8270 4030
rect 8290 4010 8305 4030
rect 8255 3980 8305 4010
rect 8255 3960 8270 3980
rect 8290 3960 8305 3980
rect 8255 3945 8305 3960
rect 8385 4030 8435 4045
rect 8385 4010 8400 4030
rect 8420 4010 8435 4030
rect 8385 3980 8435 4010
rect 8385 3960 8400 3980
rect 8420 3960 8435 3980
rect 8385 3945 8435 3960
rect 8450 4030 8500 4045
rect 8450 4010 8465 4030
rect 8485 4010 8500 4030
rect 8450 3980 8500 4010
rect 8450 3960 8465 3980
rect 8485 3960 8500 3980
rect 8450 3945 8500 3960
rect 8580 4030 8630 4045
rect 8580 4010 8595 4030
rect 8615 4010 8630 4030
rect 8580 3980 8630 4010
rect 8580 3960 8595 3980
rect 8615 3960 8630 3980
rect 8580 3945 8630 3960
rect 8645 4030 8695 4045
rect 8645 4010 8660 4030
rect 8680 4010 8695 4030
rect 8645 3980 8695 4010
rect 8645 3960 8660 3980
rect 8680 3960 8695 3980
rect 8645 3945 8695 3960
rect 8725 4030 8775 4045
rect 8725 4010 8740 4030
rect 8760 4010 8775 4030
rect 8725 3980 8775 4010
rect 8725 3960 8740 3980
rect 8760 3960 8775 3980
rect 8725 3945 8775 3960
rect 8790 4030 8840 4045
rect 8790 4010 8805 4030
rect 8825 4010 8840 4030
rect 8790 3980 8840 4010
rect 8790 3960 8805 3980
rect 8825 3960 8840 3980
rect 8790 3945 8840 3960
rect 8920 4030 8970 4045
rect 8920 4010 8935 4030
rect 8955 4010 8970 4030
rect 8920 3980 8970 4010
rect 8920 3960 8935 3980
rect 8955 3960 8970 3980
rect 8920 3945 8970 3960
rect 8985 4030 9035 4045
rect 8985 4010 9000 4030
rect 9020 4010 9035 4030
rect 8985 3980 9035 4010
rect 8985 3960 9000 3980
rect 9020 3960 9035 3980
rect 8985 3945 9035 3960
rect 9665 4005 9715 4020
rect 9665 3985 9680 4005
rect 9700 3985 9715 4005
rect 9665 3955 9715 3985
rect 9665 3935 9680 3955
rect 9700 3935 9715 3955
rect 9665 3905 9715 3935
rect 9665 3885 9680 3905
rect 9700 3885 9715 3905
rect 9665 3855 9715 3885
rect 9665 3835 9680 3855
rect 9700 3835 9715 3855
rect 9665 3820 9715 3835
rect 9775 4005 9825 4020
rect 9775 3985 9790 4005
rect 9810 3985 9825 4005
rect 9775 3955 9825 3985
rect 9775 3935 9790 3955
rect 9810 3935 9825 3955
rect 9775 3905 9825 3935
rect 9775 3885 9790 3905
rect 9810 3885 9825 3905
rect 9775 3855 9825 3885
rect 9775 3835 9790 3855
rect 9810 3835 9825 3855
rect 9775 3820 9825 3835
rect 9885 4005 9935 4020
rect 9885 3985 9900 4005
rect 9920 3985 9935 4005
rect 9885 3955 9935 3985
rect 9885 3935 9900 3955
rect 9920 3935 9935 3955
rect 9885 3905 9935 3935
rect 9885 3885 9900 3905
rect 9920 3885 9935 3905
rect 9885 3855 9935 3885
rect 9885 3835 9900 3855
rect 9920 3835 9935 3855
rect 9885 3820 9935 3835
rect 9995 4005 10045 4020
rect 9995 3985 10010 4005
rect 10030 3985 10045 4005
rect 9995 3955 10045 3985
rect 9995 3935 10010 3955
rect 10030 3935 10045 3955
rect 9995 3905 10045 3935
rect 9995 3885 10010 3905
rect 10030 3885 10045 3905
rect 9995 3855 10045 3885
rect 9995 3835 10010 3855
rect 10030 3835 10045 3855
rect 9995 3820 10045 3835
rect 10105 4005 10155 4020
rect 10205 4005 10255 4020
rect 10105 3985 10120 4005
rect 10140 3985 10155 4005
rect 10205 3985 10220 4005
rect 10240 3985 10255 4005
rect 10105 3955 10155 3985
rect 10205 3955 10255 3985
rect 10105 3935 10120 3955
rect 10140 3935 10155 3955
rect 10205 3935 10220 3955
rect 10240 3935 10255 3955
rect 10105 3905 10155 3935
rect 10205 3905 10255 3935
rect 10105 3885 10120 3905
rect 10140 3885 10155 3905
rect 10205 3885 10220 3905
rect 10240 3885 10255 3905
rect 10105 3855 10155 3885
rect 10205 3855 10255 3885
rect 10105 3835 10120 3855
rect 10140 3835 10155 3855
rect 10205 3835 10220 3855
rect 10240 3835 10255 3855
rect 10105 3820 10155 3835
rect 10205 3820 10255 3835
rect 10315 4005 10365 4020
rect 10315 3985 10330 4005
rect 10350 3985 10365 4005
rect 10315 3955 10365 3985
rect 10315 3935 10330 3955
rect 10350 3935 10365 3955
rect 10315 3905 10365 3935
rect 10315 3885 10330 3905
rect 10350 3885 10365 3905
rect 10315 3855 10365 3885
rect 10315 3835 10330 3855
rect 10350 3835 10365 3855
rect 10315 3820 10365 3835
rect 10425 4005 10475 4020
rect 10425 3985 10440 4005
rect 10460 3985 10475 4005
rect 10425 3955 10475 3985
rect 10425 3935 10440 3955
rect 10460 3935 10475 3955
rect 10425 3905 10475 3935
rect 10425 3885 10440 3905
rect 10460 3885 10475 3905
rect 10425 3855 10475 3885
rect 10425 3835 10440 3855
rect 10460 3835 10475 3855
rect 10425 3820 10475 3835
rect 10535 4005 10585 4020
rect 10535 3985 10550 4005
rect 10570 3985 10585 4005
rect 10535 3955 10585 3985
rect 10535 3935 10550 3955
rect 10570 3935 10585 3955
rect 10535 3905 10585 3935
rect 10535 3885 10550 3905
rect 10570 3885 10585 3905
rect 10535 3855 10585 3885
rect 10535 3835 10550 3855
rect 10570 3835 10585 3855
rect 10535 3820 10585 3835
rect 10645 4005 10695 4020
rect 10745 4005 10795 4020
rect 10645 3985 10660 4005
rect 10680 3985 10695 4005
rect 10745 3985 10760 4005
rect 10780 3985 10795 4005
rect 10645 3955 10695 3985
rect 10745 3955 10795 3985
rect 10645 3935 10660 3955
rect 10680 3935 10695 3955
rect 10745 3935 10760 3955
rect 10780 3935 10795 3955
rect 10645 3905 10695 3935
rect 10745 3905 10795 3935
rect 10645 3885 10660 3905
rect 10680 3885 10695 3905
rect 10745 3885 10760 3905
rect 10780 3885 10795 3905
rect 10645 3855 10695 3885
rect 10745 3855 10795 3885
rect 10645 3835 10660 3855
rect 10680 3835 10695 3855
rect 10745 3835 10760 3855
rect 10780 3835 10795 3855
rect 10645 3820 10695 3835
rect 10745 3820 10795 3835
rect 10855 4005 10905 4020
rect 10855 3985 10870 4005
rect 10890 3985 10905 4005
rect 10855 3955 10905 3985
rect 10855 3935 10870 3955
rect 10890 3935 10905 3955
rect 10855 3905 10905 3935
rect 10855 3885 10870 3905
rect 10890 3885 10905 3905
rect 10855 3855 10905 3885
rect 10855 3835 10870 3855
rect 10890 3835 10905 3855
rect 10855 3820 10905 3835
rect 10965 4005 11015 4020
rect 10965 3985 10980 4005
rect 11000 3985 11015 4005
rect 10965 3955 11015 3985
rect 10965 3935 10980 3955
rect 11000 3935 11015 3955
rect 10965 3905 11015 3935
rect 10965 3885 10980 3905
rect 11000 3885 11015 3905
rect 10965 3855 11015 3885
rect 10965 3835 10980 3855
rect 11000 3835 11015 3855
rect 10965 3820 11015 3835
rect 11075 4005 11125 4020
rect 11075 3985 11090 4005
rect 11110 3985 11125 4005
rect 11075 3955 11125 3985
rect 11075 3935 11090 3955
rect 11110 3935 11125 3955
rect 11075 3905 11125 3935
rect 11075 3885 11090 3905
rect 11110 3885 11125 3905
rect 11075 3855 11125 3885
rect 11075 3835 11090 3855
rect 11110 3835 11125 3855
rect 11075 3820 11125 3835
rect 11185 4005 11235 4020
rect 11185 3985 11200 4005
rect 11220 3985 11235 4005
rect 11185 3955 11235 3985
rect 11185 3935 11200 3955
rect 11220 3935 11235 3955
rect 11185 3905 11235 3935
rect 11185 3885 11200 3905
rect 11220 3885 11235 3905
rect 11185 3855 11235 3885
rect 11185 3835 11200 3855
rect 11220 3835 11235 3855
rect 11185 3820 11235 3835
rect 6625 3130 6665 3145
rect 6625 3110 6635 3130
rect 6655 3110 6665 3130
rect 6625 3080 6665 3110
rect 6625 3060 6635 3080
rect 6655 3060 6665 3080
rect 6625 3045 6665 3060
rect 6680 3130 6720 3145
rect 6680 3110 6690 3130
rect 6710 3110 6720 3130
rect 6680 3080 6720 3110
rect 6680 3060 6690 3080
rect 6710 3060 6720 3080
rect 6680 3045 6720 3060
rect 6735 3130 6775 3145
rect 6735 3110 6745 3130
rect 6765 3110 6775 3130
rect 6735 3080 6775 3110
rect 6735 3060 6745 3080
rect 6765 3060 6775 3080
rect 6735 3045 6775 3060
rect 6885 3130 6925 3145
rect 6885 3110 6895 3130
rect 6915 3110 6925 3130
rect 6885 3080 6925 3110
rect 6885 3060 6895 3080
rect 6915 3060 6925 3080
rect 6885 3045 6925 3060
rect 6940 3130 6980 3145
rect 6940 3110 6950 3130
rect 6970 3110 6980 3130
rect 6940 3080 6980 3110
rect 6940 3060 6950 3080
rect 6970 3060 6980 3080
rect 6940 3045 6980 3060
rect 6995 3130 7035 3145
rect 7075 3130 7115 3145
rect 6995 3110 7005 3130
rect 7025 3110 7035 3130
rect 7075 3110 7085 3130
rect 7105 3110 7115 3130
rect 6995 3080 7035 3110
rect 7075 3080 7115 3110
rect 6995 3060 7005 3080
rect 7025 3060 7035 3080
rect 7075 3060 7085 3080
rect 7105 3060 7115 3080
rect 6995 3045 7035 3060
rect 7075 3045 7115 3060
rect 7130 3130 7170 3145
rect 7130 3110 7140 3130
rect 7160 3110 7170 3130
rect 7130 3080 7170 3110
rect 7130 3060 7140 3080
rect 7160 3060 7170 3080
rect 7130 3045 7170 3060
rect 7185 3130 7225 3145
rect 7185 3110 7195 3130
rect 7215 3110 7225 3130
rect 7185 3080 7225 3110
rect 7185 3060 7195 3080
rect 7215 3060 7225 3080
rect 7185 3045 7225 3060
rect 7335 3130 7375 3145
rect 7335 3110 7345 3130
rect 7365 3110 7375 3130
rect 7335 3080 7375 3110
rect 7335 3060 7345 3080
rect 7365 3060 7375 3080
rect 7335 3045 7375 3060
rect 7390 3130 7430 3145
rect 7390 3110 7400 3130
rect 7420 3110 7430 3130
rect 7390 3080 7430 3110
rect 7390 3060 7400 3080
rect 7420 3060 7430 3080
rect 7390 3045 7430 3060
rect 7445 3130 7485 3145
rect 7445 3110 7455 3130
rect 7475 3110 7485 3130
rect 7445 3080 7485 3110
rect 7445 3060 7455 3080
rect 7475 3060 7485 3080
rect 7445 3045 7485 3060
rect 7595 3130 7635 3145
rect 7595 3110 7605 3130
rect 7625 3110 7635 3130
rect 7595 3080 7635 3110
rect 7595 3060 7605 3080
rect 7625 3060 7635 3080
rect 7595 3045 7635 3060
rect 7650 3130 7690 3145
rect 7650 3110 7660 3130
rect 7680 3110 7690 3130
rect 7650 3080 7690 3110
rect 7650 3060 7660 3080
rect 7680 3060 7690 3080
rect 7650 3045 7690 3060
rect 7705 3130 7745 3145
rect 7705 3110 7715 3130
rect 7735 3110 7745 3130
rect 7705 3080 7745 3110
rect 7705 3060 7715 3080
rect 7735 3060 7745 3080
rect 7705 3045 7745 3060
rect 7815 3130 7855 3145
rect 7815 3110 7825 3130
rect 7845 3110 7855 3130
rect 7815 3080 7855 3110
rect 7815 3060 7825 3080
rect 7845 3060 7855 3080
rect 7815 3045 7855 3060
rect 7870 3130 7910 3145
rect 7870 3110 7880 3130
rect 7900 3110 7910 3130
rect 7870 3080 7910 3110
rect 7870 3060 7880 3080
rect 7900 3060 7910 3080
rect 7870 3045 7910 3060
rect 7980 3130 8020 3145
rect 7980 3110 7990 3130
rect 8010 3110 8020 3130
rect 7980 3080 8020 3110
rect 7980 3060 7990 3080
rect 8010 3060 8020 3080
rect 7980 3045 8020 3060
rect 8035 3130 8075 3145
rect 8035 3110 8045 3130
rect 8065 3110 8075 3130
rect 8035 3080 8075 3110
rect 8035 3060 8045 3080
rect 8065 3060 8075 3080
rect 8035 3045 8075 3060
rect 8190 3130 8240 3145
rect 8190 3110 8205 3130
rect 8225 3110 8240 3130
rect 8190 3080 8240 3110
rect 8190 3060 8205 3080
rect 8225 3060 8240 3080
rect 8190 3045 8240 3060
rect 8255 3130 8305 3145
rect 8255 3110 8270 3130
rect 8290 3110 8305 3130
rect 8255 3080 8305 3110
rect 8255 3060 8270 3080
rect 8290 3060 8305 3080
rect 8255 3045 8305 3060
rect 8385 3130 8435 3145
rect 8385 3110 8400 3130
rect 8420 3110 8435 3130
rect 8385 3080 8435 3110
rect 8385 3060 8400 3080
rect 8420 3060 8435 3080
rect 8385 3045 8435 3060
rect 8450 3130 8500 3145
rect 8450 3110 8465 3130
rect 8485 3110 8500 3130
rect 8450 3080 8500 3110
rect 8450 3060 8465 3080
rect 8485 3060 8500 3080
rect 8450 3045 8500 3060
rect 8580 3130 8630 3145
rect 8580 3110 8595 3130
rect 8615 3110 8630 3130
rect 8580 3080 8630 3110
rect 8580 3060 8595 3080
rect 8615 3060 8630 3080
rect 8580 3045 8630 3060
rect 8645 3130 8695 3145
rect 8645 3110 8660 3130
rect 8680 3110 8695 3130
rect 8645 3080 8695 3110
rect 8645 3060 8660 3080
rect 8680 3060 8695 3080
rect 8645 3045 8695 3060
rect 8725 3130 8775 3145
rect 8725 3110 8740 3130
rect 8760 3110 8775 3130
rect 8725 3080 8775 3110
rect 8725 3060 8740 3080
rect 8760 3060 8775 3080
rect 8725 3045 8775 3060
rect 8790 3130 8840 3145
rect 8790 3110 8805 3130
rect 8825 3110 8840 3130
rect 8790 3080 8840 3110
rect 8790 3060 8805 3080
rect 8825 3060 8840 3080
rect 8790 3045 8840 3060
<< pdiff >>
rect 6625 3820 6665 3835
rect 6625 3800 6635 3820
rect 6655 3800 6665 3820
rect 6625 3770 6665 3800
rect 6625 3750 6635 3770
rect 6655 3750 6665 3770
rect 6625 3720 6665 3750
rect 6625 3700 6635 3720
rect 6655 3700 6665 3720
rect 6625 3670 6665 3700
rect 6625 3650 6635 3670
rect 6655 3650 6665 3670
rect 6625 3635 6665 3650
rect 6680 3820 6720 3835
rect 6680 3800 6690 3820
rect 6710 3800 6720 3820
rect 6680 3770 6720 3800
rect 6680 3750 6690 3770
rect 6710 3750 6720 3770
rect 6680 3720 6720 3750
rect 6680 3700 6690 3720
rect 6710 3700 6720 3720
rect 6680 3670 6720 3700
rect 6680 3650 6690 3670
rect 6710 3650 6720 3670
rect 6680 3635 6720 3650
rect 6735 3820 6775 3835
rect 6735 3800 6745 3820
rect 6765 3800 6775 3820
rect 6735 3770 6775 3800
rect 6735 3750 6745 3770
rect 6765 3750 6775 3770
rect 6735 3720 6775 3750
rect 6735 3700 6745 3720
rect 6765 3700 6775 3720
rect 6735 3670 6775 3700
rect 6735 3650 6745 3670
rect 6765 3650 6775 3670
rect 6735 3635 6775 3650
rect 6885 3820 6925 3835
rect 6885 3800 6895 3820
rect 6915 3800 6925 3820
rect 6885 3770 6925 3800
rect 6885 3750 6895 3770
rect 6915 3750 6925 3770
rect 6885 3720 6925 3750
rect 6885 3700 6895 3720
rect 6915 3700 6925 3720
rect 6885 3670 6925 3700
rect 6885 3650 6895 3670
rect 6915 3650 6925 3670
rect 6885 3635 6925 3650
rect 6940 3820 6980 3835
rect 6940 3800 6950 3820
rect 6970 3800 6980 3820
rect 6940 3770 6980 3800
rect 6940 3750 6950 3770
rect 6970 3750 6980 3770
rect 6940 3720 6980 3750
rect 6940 3700 6950 3720
rect 6970 3700 6980 3720
rect 6940 3670 6980 3700
rect 6940 3650 6950 3670
rect 6970 3650 6980 3670
rect 6940 3635 6980 3650
rect 6995 3820 7035 3835
rect 7075 3820 7115 3835
rect 6995 3800 7005 3820
rect 7025 3800 7035 3820
rect 7075 3800 7085 3820
rect 7105 3800 7115 3820
rect 6995 3770 7035 3800
rect 7075 3770 7115 3800
rect 6995 3750 7005 3770
rect 7025 3750 7035 3770
rect 7075 3750 7085 3770
rect 7105 3750 7115 3770
rect 6995 3720 7035 3750
rect 7075 3720 7115 3750
rect 6995 3700 7005 3720
rect 7025 3700 7035 3720
rect 7075 3700 7085 3720
rect 7105 3700 7115 3720
rect 6995 3670 7035 3700
rect 7075 3670 7115 3700
rect 6995 3650 7005 3670
rect 7025 3650 7035 3670
rect 7075 3650 7085 3670
rect 7105 3650 7115 3670
rect 6995 3635 7035 3650
rect 7075 3635 7115 3650
rect 7130 3820 7170 3835
rect 7130 3800 7140 3820
rect 7160 3800 7170 3820
rect 7130 3770 7170 3800
rect 7130 3750 7140 3770
rect 7160 3750 7170 3770
rect 7130 3720 7170 3750
rect 7130 3700 7140 3720
rect 7160 3700 7170 3720
rect 7130 3670 7170 3700
rect 7130 3650 7140 3670
rect 7160 3650 7170 3670
rect 7130 3635 7170 3650
rect 7185 3820 7225 3835
rect 7185 3800 7195 3820
rect 7215 3800 7225 3820
rect 7185 3770 7225 3800
rect 7185 3750 7195 3770
rect 7215 3750 7225 3770
rect 7185 3720 7225 3750
rect 7185 3700 7195 3720
rect 7215 3700 7225 3720
rect 7185 3670 7225 3700
rect 7185 3650 7195 3670
rect 7215 3650 7225 3670
rect 7185 3635 7225 3650
rect 7335 3820 7375 3835
rect 7335 3800 7345 3820
rect 7365 3800 7375 3820
rect 7335 3770 7375 3800
rect 7335 3750 7345 3770
rect 7365 3750 7375 3770
rect 7335 3720 7375 3750
rect 7335 3700 7345 3720
rect 7365 3700 7375 3720
rect 7335 3670 7375 3700
rect 7335 3650 7345 3670
rect 7365 3650 7375 3670
rect 7335 3635 7375 3650
rect 7390 3820 7430 3835
rect 7390 3800 7400 3820
rect 7420 3800 7430 3820
rect 7390 3770 7430 3800
rect 7390 3750 7400 3770
rect 7420 3750 7430 3770
rect 7390 3720 7430 3750
rect 7390 3700 7400 3720
rect 7420 3700 7430 3720
rect 7390 3670 7430 3700
rect 7390 3650 7400 3670
rect 7420 3650 7430 3670
rect 7390 3635 7430 3650
rect 7445 3820 7485 3835
rect 7445 3800 7455 3820
rect 7475 3800 7485 3820
rect 7445 3770 7485 3800
rect 7445 3750 7455 3770
rect 7475 3750 7485 3770
rect 7445 3720 7485 3750
rect 7445 3700 7455 3720
rect 7475 3700 7485 3720
rect 7445 3670 7485 3700
rect 7445 3650 7455 3670
rect 7475 3650 7485 3670
rect 7445 3635 7485 3650
rect 7590 3820 7630 3835
rect 7590 3800 7600 3820
rect 7620 3800 7630 3820
rect 7590 3770 7630 3800
rect 7590 3750 7600 3770
rect 7620 3750 7630 3770
rect 7590 3720 7630 3750
rect 7590 3700 7600 3720
rect 7620 3700 7630 3720
rect 7590 3670 7630 3700
rect 7590 3650 7600 3670
rect 7620 3650 7630 3670
rect 7590 3635 7630 3650
rect 7645 3820 7685 3835
rect 7645 3800 7655 3820
rect 7675 3800 7685 3820
rect 7645 3770 7685 3800
rect 7645 3750 7655 3770
rect 7675 3750 7685 3770
rect 7645 3720 7685 3750
rect 7645 3700 7655 3720
rect 7675 3700 7685 3720
rect 7645 3670 7685 3700
rect 7645 3650 7655 3670
rect 7675 3650 7685 3670
rect 7645 3635 7685 3650
rect 7755 3820 7795 3835
rect 7755 3800 7765 3820
rect 7785 3800 7795 3820
rect 7755 3770 7795 3800
rect 7755 3750 7765 3770
rect 7785 3750 7795 3770
rect 7755 3720 7795 3750
rect 7755 3700 7765 3720
rect 7785 3700 7795 3720
rect 7755 3670 7795 3700
rect 7755 3650 7765 3670
rect 7785 3650 7795 3670
rect 7755 3635 7795 3650
rect 7810 3820 7850 3835
rect 7810 3800 7820 3820
rect 7840 3800 7850 3820
rect 7810 3770 7850 3800
rect 7810 3750 7820 3770
rect 7840 3750 7850 3770
rect 7810 3720 7850 3750
rect 7810 3700 7820 3720
rect 7840 3700 7850 3720
rect 7810 3670 7850 3700
rect 7810 3650 7820 3670
rect 7840 3650 7850 3670
rect 7810 3635 7850 3650
rect 7920 3820 7960 3835
rect 7920 3800 7930 3820
rect 7950 3800 7960 3820
rect 7920 3770 7960 3800
rect 7920 3750 7930 3770
rect 7950 3750 7960 3770
rect 7920 3720 7960 3750
rect 7920 3700 7930 3720
rect 7950 3700 7960 3720
rect 7920 3670 7960 3700
rect 7920 3650 7930 3670
rect 7950 3650 7960 3670
rect 7920 3635 7960 3650
rect 7975 3820 8015 3835
rect 7975 3800 7985 3820
rect 8005 3800 8015 3820
rect 7975 3770 8015 3800
rect 7975 3750 7985 3770
rect 8005 3750 8015 3770
rect 7975 3720 8015 3750
rect 7975 3700 7985 3720
rect 8005 3700 8015 3720
rect 7975 3670 8015 3700
rect 7975 3650 7985 3670
rect 8005 3650 8015 3670
rect 7975 3635 8015 3650
rect 8190 3820 8240 3835
rect 8190 3800 8205 3820
rect 8225 3800 8240 3820
rect 8190 3770 8240 3800
rect 8190 3750 8205 3770
rect 8225 3750 8240 3770
rect 8190 3720 8240 3750
rect 8190 3700 8205 3720
rect 8225 3700 8240 3720
rect 8190 3670 8240 3700
rect 8190 3650 8205 3670
rect 8225 3650 8240 3670
rect 8190 3635 8240 3650
rect 8255 3820 8305 3835
rect 8255 3800 8270 3820
rect 8290 3800 8305 3820
rect 8255 3770 8305 3800
rect 8255 3750 8270 3770
rect 8290 3750 8305 3770
rect 8255 3720 8305 3750
rect 8255 3700 8270 3720
rect 8290 3700 8305 3720
rect 8255 3670 8305 3700
rect 8255 3650 8270 3670
rect 8290 3650 8305 3670
rect 8255 3635 8305 3650
rect 8385 3820 8435 3835
rect 8385 3800 8400 3820
rect 8420 3800 8435 3820
rect 8385 3770 8435 3800
rect 8385 3750 8400 3770
rect 8420 3750 8435 3770
rect 8385 3720 8435 3750
rect 8385 3700 8400 3720
rect 8420 3700 8435 3720
rect 8385 3670 8435 3700
rect 8385 3650 8400 3670
rect 8420 3650 8435 3670
rect 8385 3635 8435 3650
rect 8450 3820 8500 3835
rect 8450 3800 8465 3820
rect 8485 3800 8500 3820
rect 8450 3770 8500 3800
rect 8450 3750 8465 3770
rect 8485 3750 8500 3770
rect 8450 3720 8500 3750
rect 8450 3700 8465 3720
rect 8485 3700 8500 3720
rect 8450 3670 8500 3700
rect 8450 3650 8465 3670
rect 8485 3650 8500 3670
rect 8450 3635 8500 3650
rect 8580 3820 8630 3835
rect 8580 3800 8595 3820
rect 8615 3800 8630 3820
rect 8580 3770 8630 3800
rect 8580 3750 8595 3770
rect 8615 3750 8630 3770
rect 8580 3720 8630 3750
rect 8580 3700 8595 3720
rect 8615 3700 8630 3720
rect 8580 3670 8630 3700
rect 8580 3650 8595 3670
rect 8615 3650 8630 3670
rect 8580 3635 8630 3650
rect 8645 3820 8695 3835
rect 8645 3800 8660 3820
rect 8680 3800 8695 3820
rect 8645 3770 8695 3800
rect 8645 3750 8660 3770
rect 8680 3750 8695 3770
rect 8645 3720 8695 3750
rect 8645 3700 8660 3720
rect 8680 3700 8695 3720
rect 8645 3670 8695 3700
rect 8645 3650 8660 3670
rect 8680 3650 8695 3670
rect 8645 3635 8695 3650
rect 8725 3820 8775 3835
rect 8725 3800 8740 3820
rect 8760 3800 8775 3820
rect 8725 3770 8775 3800
rect 8725 3750 8740 3770
rect 8760 3750 8775 3770
rect 8725 3720 8775 3750
rect 8725 3700 8740 3720
rect 8760 3700 8775 3720
rect 8725 3670 8775 3700
rect 8725 3650 8740 3670
rect 8760 3650 8775 3670
rect 8725 3635 8775 3650
rect 8790 3820 8840 3835
rect 8790 3800 8805 3820
rect 8825 3800 8840 3820
rect 8790 3770 8840 3800
rect 8790 3750 8805 3770
rect 8825 3750 8840 3770
rect 8790 3720 8840 3750
rect 8790 3700 8805 3720
rect 8825 3700 8840 3720
rect 8790 3670 8840 3700
rect 8790 3650 8805 3670
rect 8825 3650 8840 3670
rect 8790 3635 8840 3650
rect 9765 3455 9815 3470
rect 6625 3440 6665 3455
rect 6625 3420 6635 3440
rect 6655 3420 6665 3440
rect 6625 3390 6665 3420
rect 6625 3370 6635 3390
rect 6655 3370 6665 3390
rect 6625 3340 6665 3370
rect 6625 3320 6635 3340
rect 6655 3320 6665 3340
rect 6625 3290 6665 3320
rect 6625 3270 6635 3290
rect 6655 3270 6665 3290
rect 6625 3255 6665 3270
rect 6680 3440 6720 3455
rect 6680 3420 6690 3440
rect 6710 3420 6720 3440
rect 6680 3390 6720 3420
rect 6680 3370 6690 3390
rect 6710 3370 6720 3390
rect 6680 3340 6720 3370
rect 6680 3320 6690 3340
rect 6710 3320 6720 3340
rect 6680 3290 6720 3320
rect 6680 3270 6690 3290
rect 6710 3270 6720 3290
rect 6680 3255 6720 3270
rect 6735 3440 6775 3455
rect 6735 3420 6745 3440
rect 6765 3420 6775 3440
rect 6735 3390 6775 3420
rect 6735 3370 6745 3390
rect 6765 3370 6775 3390
rect 6735 3340 6775 3370
rect 6735 3320 6745 3340
rect 6765 3320 6775 3340
rect 6735 3290 6775 3320
rect 6735 3270 6745 3290
rect 6765 3270 6775 3290
rect 6735 3255 6775 3270
rect 6885 3440 6925 3455
rect 6885 3420 6895 3440
rect 6915 3420 6925 3440
rect 6885 3390 6925 3420
rect 6885 3370 6895 3390
rect 6915 3370 6925 3390
rect 6885 3340 6925 3370
rect 6885 3320 6895 3340
rect 6915 3320 6925 3340
rect 6885 3290 6925 3320
rect 6885 3270 6895 3290
rect 6915 3270 6925 3290
rect 6885 3255 6925 3270
rect 6940 3440 6980 3455
rect 6940 3420 6950 3440
rect 6970 3420 6980 3440
rect 6940 3390 6980 3420
rect 6940 3370 6950 3390
rect 6970 3370 6980 3390
rect 6940 3340 6980 3370
rect 6940 3320 6950 3340
rect 6970 3320 6980 3340
rect 6940 3290 6980 3320
rect 6940 3270 6950 3290
rect 6970 3270 6980 3290
rect 6940 3255 6980 3270
rect 6995 3440 7035 3455
rect 7075 3440 7115 3455
rect 6995 3420 7005 3440
rect 7025 3420 7035 3440
rect 7075 3420 7085 3440
rect 7105 3420 7115 3440
rect 6995 3390 7035 3420
rect 7075 3390 7115 3420
rect 6995 3370 7005 3390
rect 7025 3370 7035 3390
rect 7075 3370 7085 3390
rect 7105 3370 7115 3390
rect 6995 3340 7035 3370
rect 7075 3340 7115 3370
rect 6995 3320 7005 3340
rect 7025 3320 7035 3340
rect 7075 3320 7085 3340
rect 7105 3320 7115 3340
rect 6995 3290 7035 3320
rect 7075 3290 7115 3320
rect 6995 3270 7005 3290
rect 7025 3270 7035 3290
rect 7075 3270 7085 3290
rect 7105 3270 7115 3290
rect 6995 3255 7035 3270
rect 7075 3255 7115 3270
rect 7130 3440 7170 3455
rect 7130 3420 7140 3440
rect 7160 3420 7170 3440
rect 7130 3390 7170 3420
rect 7130 3370 7140 3390
rect 7160 3370 7170 3390
rect 7130 3340 7170 3370
rect 7130 3320 7140 3340
rect 7160 3320 7170 3340
rect 7130 3290 7170 3320
rect 7130 3270 7140 3290
rect 7160 3270 7170 3290
rect 7130 3255 7170 3270
rect 7185 3440 7225 3455
rect 7185 3420 7195 3440
rect 7215 3420 7225 3440
rect 7185 3390 7225 3420
rect 7185 3370 7195 3390
rect 7215 3370 7225 3390
rect 7185 3340 7225 3370
rect 7185 3320 7195 3340
rect 7215 3320 7225 3340
rect 7185 3290 7225 3320
rect 7185 3270 7195 3290
rect 7215 3270 7225 3290
rect 7185 3255 7225 3270
rect 7335 3440 7375 3455
rect 7335 3420 7345 3440
rect 7365 3420 7375 3440
rect 7335 3390 7375 3420
rect 7335 3370 7345 3390
rect 7365 3370 7375 3390
rect 7335 3340 7375 3370
rect 7335 3320 7345 3340
rect 7365 3320 7375 3340
rect 7335 3290 7375 3320
rect 7335 3270 7345 3290
rect 7365 3270 7375 3290
rect 7335 3255 7375 3270
rect 7390 3440 7430 3455
rect 7390 3420 7400 3440
rect 7420 3420 7430 3440
rect 7390 3390 7430 3420
rect 7390 3370 7400 3390
rect 7420 3370 7430 3390
rect 7390 3340 7430 3370
rect 7390 3320 7400 3340
rect 7420 3320 7430 3340
rect 7390 3290 7430 3320
rect 7390 3270 7400 3290
rect 7420 3270 7430 3290
rect 7390 3255 7430 3270
rect 7445 3440 7485 3455
rect 7445 3420 7455 3440
rect 7475 3420 7485 3440
rect 7445 3390 7485 3420
rect 7445 3370 7455 3390
rect 7475 3370 7485 3390
rect 7445 3340 7485 3370
rect 7445 3320 7455 3340
rect 7475 3320 7485 3340
rect 7445 3290 7485 3320
rect 7445 3270 7455 3290
rect 7475 3270 7485 3290
rect 7445 3255 7485 3270
rect 7595 3440 7635 3455
rect 7595 3420 7605 3440
rect 7625 3420 7635 3440
rect 7595 3390 7635 3420
rect 7595 3370 7605 3390
rect 7625 3370 7635 3390
rect 7595 3340 7635 3370
rect 7595 3320 7605 3340
rect 7625 3320 7635 3340
rect 7595 3290 7635 3320
rect 7595 3270 7605 3290
rect 7625 3270 7635 3290
rect 7595 3255 7635 3270
rect 7650 3440 7690 3455
rect 7650 3420 7660 3440
rect 7680 3420 7690 3440
rect 7650 3390 7690 3420
rect 7650 3370 7660 3390
rect 7680 3370 7690 3390
rect 7650 3340 7690 3370
rect 7650 3320 7660 3340
rect 7680 3320 7690 3340
rect 7650 3290 7690 3320
rect 7650 3270 7660 3290
rect 7680 3270 7690 3290
rect 7650 3255 7690 3270
rect 7705 3440 7745 3455
rect 7705 3420 7715 3440
rect 7735 3420 7745 3440
rect 7705 3390 7745 3420
rect 7705 3370 7715 3390
rect 7735 3370 7745 3390
rect 7705 3340 7745 3370
rect 7705 3320 7715 3340
rect 7735 3320 7745 3340
rect 7705 3290 7745 3320
rect 7705 3270 7715 3290
rect 7735 3270 7745 3290
rect 7705 3255 7745 3270
rect 7815 3440 7855 3455
rect 7815 3420 7825 3440
rect 7845 3420 7855 3440
rect 7815 3390 7855 3420
rect 7815 3370 7825 3390
rect 7845 3370 7855 3390
rect 7815 3340 7855 3370
rect 7815 3320 7825 3340
rect 7845 3320 7855 3340
rect 7815 3290 7855 3320
rect 7815 3270 7825 3290
rect 7845 3270 7855 3290
rect 7815 3255 7855 3270
rect 7870 3440 7910 3455
rect 7870 3420 7880 3440
rect 7900 3420 7910 3440
rect 7870 3390 7910 3420
rect 7870 3370 7880 3390
rect 7900 3370 7910 3390
rect 7870 3340 7910 3370
rect 7870 3320 7880 3340
rect 7900 3320 7910 3340
rect 7870 3290 7910 3320
rect 7870 3270 7880 3290
rect 7900 3270 7910 3290
rect 7870 3255 7910 3270
rect 7980 3440 8020 3455
rect 7980 3420 7990 3440
rect 8010 3420 8020 3440
rect 7980 3390 8020 3420
rect 7980 3370 7990 3390
rect 8010 3370 8020 3390
rect 7980 3340 8020 3370
rect 7980 3320 7990 3340
rect 8010 3320 8020 3340
rect 7980 3290 8020 3320
rect 7980 3270 7990 3290
rect 8010 3270 8020 3290
rect 7980 3255 8020 3270
rect 8035 3440 8075 3455
rect 8035 3420 8045 3440
rect 8065 3420 8075 3440
rect 8035 3390 8075 3420
rect 8035 3370 8045 3390
rect 8065 3370 8075 3390
rect 8035 3340 8075 3370
rect 8035 3320 8045 3340
rect 8065 3320 8075 3340
rect 8035 3290 8075 3320
rect 8035 3270 8045 3290
rect 8065 3270 8075 3290
rect 8035 3255 8075 3270
rect 8190 3440 8240 3455
rect 8190 3420 8205 3440
rect 8225 3420 8240 3440
rect 8190 3390 8240 3420
rect 8190 3370 8205 3390
rect 8225 3370 8240 3390
rect 8190 3340 8240 3370
rect 8190 3320 8205 3340
rect 8225 3320 8240 3340
rect 8190 3290 8240 3320
rect 8190 3270 8205 3290
rect 8225 3270 8240 3290
rect 8190 3255 8240 3270
rect 8255 3440 8305 3455
rect 8255 3420 8270 3440
rect 8290 3420 8305 3440
rect 8255 3390 8305 3420
rect 8255 3370 8270 3390
rect 8290 3370 8305 3390
rect 8255 3340 8305 3370
rect 8255 3320 8270 3340
rect 8290 3320 8305 3340
rect 8255 3290 8305 3320
rect 8255 3270 8270 3290
rect 8290 3270 8305 3290
rect 8255 3255 8305 3270
rect 8385 3440 8435 3455
rect 8385 3420 8400 3440
rect 8420 3420 8435 3440
rect 8385 3390 8435 3420
rect 8385 3370 8400 3390
rect 8420 3370 8435 3390
rect 8385 3340 8435 3370
rect 8385 3320 8400 3340
rect 8420 3320 8435 3340
rect 8385 3290 8435 3320
rect 8385 3270 8400 3290
rect 8420 3270 8435 3290
rect 8385 3255 8435 3270
rect 8450 3440 8500 3455
rect 8450 3420 8465 3440
rect 8485 3420 8500 3440
rect 8450 3390 8500 3420
rect 8450 3370 8465 3390
rect 8485 3370 8500 3390
rect 8450 3340 8500 3370
rect 8450 3320 8465 3340
rect 8485 3320 8500 3340
rect 8450 3290 8500 3320
rect 8450 3270 8465 3290
rect 8485 3270 8500 3290
rect 8450 3255 8500 3270
rect 8580 3440 8630 3455
rect 8580 3420 8595 3440
rect 8615 3420 8630 3440
rect 8580 3390 8630 3420
rect 8580 3370 8595 3390
rect 8615 3370 8630 3390
rect 8580 3340 8630 3370
rect 8580 3320 8595 3340
rect 8615 3320 8630 3340
rect 8580 3290 8630 3320
rect 8580 3270 8595 3290
rect 8615 3270 8630 3290
rect 8580 3255 8630 3270
rect 8645 3440 8695 3455
rect 8645 3420 8660 3440
rect 8680 3420 8695 3440
rect 8645 3390 8695 3420
rect 8645 3370 8660 3390
rect 8680 3370 8695 3390
rect 8645 3340 8695 3370
rect 8645 3320 8660 3340
rect 8680 3320 8695 3340
rect 8645 3290 8695 3320
rect 8645 3270 8660 3290
rect 8680 3270 8695 3290
rect 8645 3255 8695 3270
rect 8725 3440 8775 3455
rect 8725 3420 8740 3440
rect 8760 3420 8775 3440
rect 8725 3390 8775 3420
rect 8725 3370 8740 3390
rect 8760 3370 8775 3390
rect 8725 3340 8775 3370
rect 8725 3320 8740 3340
rect 8760 3320 8775 3340
rect 8725 3290 8775 3320
rect 8725 3270 8740 3290
rect 8760 3270 8775 3290
rect 8725 3255 8775 3270
rect 8790 3440 8840 3455
rect 8790 3420 8805 3440
rect 8825 3420 8840 3440
rect 8790 3390 8840 3420
rect 8790 3370 8805 3390
rect 8825 3370 8840 3390
rect 8790 3340 8840 3370
rect 8790 3320 8805 3340
rect 8825 3320 8840 3340
rect 8790 3290 8840 3320
rect 8790 3270 8805 3290
rect 8825 3270 8840 3290
rect 8790 3255 8840 3270
rect 8920 3440 8970 3455
rect 8920 3420 8935 3440
rect 8955 3420 8970 3440
rect 8920 3390 8970 3420
rect 8920 3370 8935 3390
rect 8955 3370 8970 3390
rect 8920 3340 8970 3370
rect 8920 3320 8935 3340
rect 8955 3320 8970 3340
rect 8920 3290 8970 3320
rect 8920 3270 8935 3290
rect 8955 3270 8970 3290
rect 8920 3255 8970 3270
rect 8985 3440 9035 3455
rect 8985 3420 9000 3440
rect 9020 3420 9035 3440
rect 8985 3390 9035 3420
rect 8985 3370 9000 3390
rect 9020 3370 9035 3390
rect 8985 3340 9035 3370
rect 8985 3320 9000 3340
rect 9020 3320 9035 3340
rect 8985 3290 9035 3320
rect 8985 3270 9000 3290
rect 9020 3270 9035 3290
rect 9765 3435 9780 3455
rect 9800 3435 9815 3455
rect 9765 3405 9815 3435
rect 9765 3385 9780 3405
rect 9800 3385 9815 3405
rect 9765 3355 9815 3385
rect 9765 3335 9780 3355
rect 9800 3335 9815 3355
rect 9765 3305 9815 3335
rect 9765 3285 9780 3305
rect 9800 3285 9815 3305
rect 9765 3270 9815 3285
rect 9875 3455 9925 3470
rect 9875 3435 9890 3455
rect 9910 3435 9925 3455
rect 9875 3405 9925 3435
rect 9875 3385 9890 3405
rect 9910 3385 9925 3405
rect 9875 3355 9925 3385
rect 9875 3335 9890 3355
rect 9910 3335 9925 3355
rect 9875 3305 9925 3335
rect 9875 3285 9890 3305
rect 9910 3285 9925 3305
rect 9875 3270 9925 3285
rect 9985 3455 10035 3470
rect 9985 3435 10000 3455
rect 10020 3435 10035 3455
rect 9985 3405 10035 3435
rect 9985 3385 10000 3405
rect 10020 3385 10035 3405
rect 9985 3355 10035 3385
rect 9985 3335 10000 3355
rect 10020 3335 10035 3355
rect 9985 3305 10035 3335
rect 9985 3285 10000 3305
rect 10020 3285 10035 3305
rect 9985 3270 10035 3285
rect 10095 3455 10145 3470
rect 10095 3435 10110 3455
rect 10130 3435 10145 3455
rect 10095 3405 10145 3435
rect 10095 3385 10110 3405
rect 10130 3385 10145 3405
rect 10095 3355 10145 3385
rect 10095 3335 10110 3355
rect 10130 3335 10145 3355
rect 10095 3305 10145 3335
rect 10095 3285 10110 3305
rect 10130 3285 10145 3305
rect 10095 3270 10145 3285
rect 10205 3455 10255 3470
rect 10205 3435 10220 3455
rect 10240 3435 10255 3455
rect 10205 3405 10255 3435
rect 10205 3385 10220 3405
rect 10240 3385 10255 3405
rect 10205 3355 10255 3385
rect 10205 3335 10220 3355
rect 10240 3335 10255 3355
rect 10205 3305 10255 3335
rect 10205 3285 10220 3305
rect 10240 3285 10255 3305
rect 10205 3270 10255 3285
rect 10315 3455 10365 3470
rect 10315 3435 10330 3455
rect 10350 3435 10365 3455
rect 10315 3405 10365 3435
rect 10315 3385 10330 3405
rect 10350 3385 10365 3405
rect 10315 3355 10365 3385
rect 10315 3335 10330 3355
rect 10350 3335 10365 3355
rect 10315 3305 10365 3335
rect 10315 3285 10330 3305
rect 10350 3285 10365 3305
rect 10315 3270 10365 3285
rect 10425 3455 10475 3470
rect 10525 3455 10575 3470
rect 10425 3435 10440 3455
rect 10460 3435 10475 3455
rect 10525 3435 10540 3455
rect 10560 3435 10575 3455
rect 10425 3405 10475 3435
rect 10525 3405 10575 3435
rect 10425 3385 10440 3405
rect 10460 3385 10475 3405
rect 10525 3385 10540 3405
rect 10560 3385 10575 3405
rect 10425 3355 10475 3385
rect 10525 3355 10575 3385
rect 10425 3335 10440 3355
rect 10460 3335 10475 3355
rect 10525 3335 10540 3355
rect 10560 3335 10575 3355
rect 10425 3305 10475 3335
rect 10525 3305 10575 3335
rect 10425 3285 10440 3305
rect 10460 3285 10475 3305
rect 10525 3285 10540 3305
rect 10560 3285 10575 3305
rect 10425 3270 10475 3285
rect 10525 3270 10575 3285
rect 10635 3455 10685 3470
rect 10635 3435 10650 3455
rect 10670 3435 10685 3455
rect 10635 3405 10685 3435
rect 10635 3385 10650 3405
rect 10670 3385 10685 3405
rect 10635 3355 10685 3385
rect 10635 3335 10650 3355
rect 10670 3335 10685 3355
rect 10635 3305 10685 3335
rect 10635 3285 10650 3305
rect 10670 3285 10685 3305
rect 10635 3270 10685 3285
rect 10745 3455 10795 3470
rect 10745 3435 10760 3455
rect 10780 3435 10795 3455
rect 10745 3405 10795 3435
rect 10745 3385 10760 3405
rect 10780 3385 10795 3405
rect 10745 3355 10795 3385
rect 10745 3335 10760 3355
rect 10780 3335 10795 3355
rect 10745 3305 10795 3335
rect 10745 3285 10760 3305
rect 10780 3285 10795 3305
rect 10745 3270 10795 3285
rect 10855 3455 10905 3470
rect 10855 3435 10870 3455
rect 10890 3435 10905 3455
rect 10855 3405 10905 3435
rect 10855 3385 10870 3405
rect 10890 3385 10905 3405
rect 10855 3355 10905 3385
rect 10855 3335 10870 3355
rect 10890 3335 10905 3355
rect 10855 3305 10905 3335
rect 10855 3285 10870 3305
rect 10890 3285 10905 3305
rect 10855 3270 10905 3285
rect 10965 3455 11015 3470
rect 10965 3435 10980 3455
rect 11000 3435 11015 3455
rect 10965 3405 11015 3435
rect 10965 3385 10980 3405
rect 11000 3385 11015 3405
rect 10965 3355 11015 3385
rect 10965 3335 10980 3355
rect 11000 3335 11015 3355
rect 10965 3305 11015 3335
rect 10965 3285 10980 3305
rect 11000 3285 11015 3305
rect 10965 3270 11015 3285
rect 11075 3455 11125 3470
rect 11075 3435 11090 3455
rect 11110 3435 11125 3455
rect 11075 3405 11125 3435
rect 11075 3385 11090 3405
rect 11110 3385 11125 3405
rect 11075 3355 11125 3385
rect 11075 3335 11090 3355
rect 11110 3335 11125 3355
rect 11075 3305 11125 3335
rect 11075 3285 11090 3305
rect 11110 3285 11125 3305
rect 11075 3270 11125 3285
rect 11185 3455 11235 3470
rect 11185 3435 11200 3455
rect 11220 3435 11235 3455
rect 11185 3405 11235 3435
rect 11185 3385 11200 3405
rect 11220 3385 11235 3405
rect 11185 3355 11235 3385
rect 11185 3335 11200 3355
rect 11220 3335 11235 3355
rect 11185 3305 11235 3335
rect 11185 3285 11200 3305
rect 11220 3285 11235 3305
rect 11185 3270 11235 3285
rect 8985 3255 9035 3270
<< ndiffc >>
rect 6635 4010 6655 4030
rect 6635 3960 6655 3980
rect 6690 4010 6710 4030
rect 6690 3960 6710 3980
rect 6745 4010 6765 4030
rect 6745 3960 6765 3980
rect 6895 4010 6915 4030
rect 6895 3960 6915 3980
rect 6950 4010 6970 4030
rect 6950 3960 6970 3980
rect 7005 4010 7025 4030
rect 7085 4010 7105 4030
rect 7005 3960 7025 3980
rect 7085 3960 7105 3980
rect 7140 4010 7160 4030
rect 7140 3960 7160 3980
rect 7195 4010 7215 4030
rect 7195 3960 7215 3980
rect 7345 4010 7365 4030
rect 7345 3960 7365 3980
rect 7400 4010 7420 4030
rect 7400 3960 7420 3980
rect 7455 4010 7475 4030
rect 7455 3960 7475 3980
rect 7600 4010 7620 4030
rect 7600 3960 7620 3980
rect 7655 4010 7675 4030
rect 7655 3960 7675 3980
rect 7765 4010 7785 4030
rect 7765 3960 7785 3980
rect 7820 4010 7840 4030
rect 7820 3960 7840 3980
rect 7930 4010 7950 4030
rect 7930 3960 7950 3980
rect 7985 4010 8005 4030
rect 7985 3960 8005 3980
rect 8205 4010 8225 4030
rect 8205 3960 8225 3980
rect 8270 4010 8290 4030
rect 8270 3960 8290 3980
rect 8400 4010 8420 4030
rect 8400 3960 8420 3980
rect 8465 4010 8485 4030
rect 8465 3960 8485 3980
rect 8595 4010 8615 4030
rect 8595 3960 8615 3980
rect 8660 4010 8680 4030
rect 8660 3960 8680 3980
rect 8740 4010 8760 4030
rect 8740 3960 8760 3980
rect 8805 4010 8825 4030
rect 8805 3960 8825 3980
rect 8935 4010 8955 4030
rect 8935 3960 8955 3980
rect 9000 4010 9020 4030
rect 9000 3960 9020 3980
rect 9680 3985 9700 4005
rect 9680 3935 9700 3955
rect 9680 3885 9700 3905
rect 9680 3835 9700 3855
rect 9790 3985 9810 4005
rect 9790 3935 9810 3955
rect 9790 3885 9810 3905
rect 9790 3835 9810 3855
rect 9900 3985 9920 4005
rect 9900 3935 9920 3955
rect 9900 3885 9920 3905
rect 9900 3835 9920 3855
rect 10010 3985 10030 4005
rect 10010 3935 10030 3955
rect 10010 3885 10030 3905
rect 10010 3835 10030 3855
rect 10120 3985 10140 4005
rect 10220 3985 10240 4005
rect 10120 3935 10140 3955
rect 10220 3935 10240 3955
rect 10120 3885 10140 3905
rect 10220 3885 10240 3905
rect 10120 3835 10140 3855
rect 10220 3835 10240 3855
rect 10330 3985 10350 4005
rect 10330 3935 10350 3955
rect 10330 3885 10350 3905
rect 10330 3835 10350 3855
rect 10440 3985 10460 4005
rect 10440 3935 10460 3955
rect 10440 3885 10460 3905
rect 10440 3835 10460 3855
rect 10550 3985 10570 4005
rect 10550 3935 10570 3955
rect 10550 3885 10570 3905
rect 10550 3835 10570 3855
rect 10660 3985 10680 4005
rect 10760 3985 10780 4005
rect 10660 3935 10680 3955
rect 10760 3935 10780 3955
rect 10660 3885 10680 3905
rect 10760 3885 10780 3905
rect 10660 3835 10680 3855
rect 10760 3835 10780 3855
rect 10870 3985 10890 4005
rect 10870 3935 10890 3955
rect 10870 3885 10890 3905
rect 10870 3835 10890 3855
rect 10980 3985 11000 4005
rect 10980 3935 11000 3955
rect 10980 3885 11000 3905
rect 10980 3835 11000 3855
rect 11090 3985 11110 4005
rect 11090 3935 11110 3955
rect 11090 3885 11110 3905
rect 11090 3835 11110 3855
rect 11200 3985 11220 4005
rect 11200 3935 11220 3955
rect 11200 3885 11220 3905
rect 11200 3835 11220 3855
rect 6635 3110 6655 3130
rect 6635 3060 6655 3080
rect 6690 3110 6710 3130
rect 6690 3060 6710 3080
rect 6745 3110 6765 3130
rect 6745 3060 6765 3080
rect 6895 3110 6915 3130
rect 6895 3060 6915 3080
rect 6950 3110 6970 3130
rect 6950 3060 6970 3080
rect 7005 3110 7025 3130
rect 7085 3110 7105 3130
rect 7005 3060 7025 3080
rect 7085 3060 7105 3080
rect 7140 3110 7160 3130
rect 7140 3060 7160 3080
rect 7195 3110 7215 3130
rect 7195 3060 7215 3080
rect 7345 3110 7365 3130
rect 7345 3060 7365 3080
rect 7400 3110 7420 3130
rect 7400 3060 7420 3080
rect 7455 3110 7475 3130
rect 7455 3060 7475 3080
rect 7605 3110 7625 3130
rect 7605 3060 7625 3080
rect 7660 3110 7680 3130
rect 7660 3060 7680 3080
rect 7715 3110 7735 3130
rect 7715 3060 7735 3080
rect 7825 3110 7845 3130
rect 7825 3060 7845 3080
rect 7880 3110 7900 3130
rect 7880 3060 7900 3080
rect 7990 3110 8010 3130
rect 7990 3060 8010 3080
rect 8045 3110 8065 3130
rect 8045 3060 8065 3080
rect 8205 3110 8225 3130
rect 8205 3060 8225 3080
rect 8270 3110 8290 3130
rect 8270 3060 8290 3080
rect 8400 3110 8420 3130
rect 8400 3060 8420 3080
rect 8465 3110 8485 3130
rect 8465 3060 8485 3080
rect 8595 3110 8615 3130
rect 8595 3060 8615 3080
rect 8660 3110 8680 3130
rect 8660 3060 8680 3080
rect 8740 3110 8760 3130
rect 8740 3060 8760 3080
rect 8805 3110 8825 3130
rect 8805 3060 8825 3080
<< pdiffc >>
rect 6635 3800 6655 3820
rect 6635 3750 6655 3770
rect 6635 3700 6655 3720
rect 6635 3650 6655 3670
rect 6690 3800 6710 3820
rect 6690 3750 6710 3770
rect 6690 3700 6710 3720
rect 6690 3650 6710 3670
rect 6745 3800 6765 3820
rect 6745 3750 6765 3770
rect 6745 3700 6765 3720
rect 6745 3650 6765 3670
rect 6895 3800 6915 3820
rect 6895 3750 6915 3770
rect 6895 3700 6915 3720
rect 6895 3650 6915 3670
rect 6950 3800 6970 3820
rect 6950 3750 6970 3770
rect 6950 3700 6970 3720
rect 6950 3650 6970 3670
rect 7005 3800 7025 3820
rect 7085 3800 7105 3820
rect 7005 3750 7025 3770
rect 7085 3750 7105 3770
rect 7005 3700 7025 3720
rect 7085 3700 7105 3720
rect 7005 3650 7025 3670
rect 7085 3650 7105 3670
rect 7140 3800 7160 3820
rect 7140 3750 7160 3770
rect 7140 3700 7160 3720
rect 7140 3650 7160 3670
rect 7195 3800 7215 3820
rect 7195 3750 7215 3770
rect 7195 3700 7215 3720
rect 7195 3650 7215 3670
rect 7345 3800 7365 3820
rect 7345 3750 7365 3770
rect 7345 3700 7365 3720
rect 7345 3650 7365 3670
rect 7400 3800 7420 3820
rect 7400 3750 7420 3770
rect 7400 3700 7420 3720
rect 7400 3650 7420 3670
rect 7455 3800 7475 3820
rect 7455 3750 7475 3770
rect 7455 3700 7475 3720
rect 7455 3650 7475 3670
rect 7600 3800 7620 3820
rect 7600 3750 7620 3770
rect 7600 3700 7620 3720
rect 7600 3650 7620 3670
rect 7655 3800 7675 3820
rect 7655 3750 7675 3770
rect 7655 3700 7675 3720
rect 7655 3650 7675 3670
rect 7765 3800 7785 3820
rect 7765 3750 7785 3770
rect 7765 3700 7785 3720
rect 7765 3650 7785 3670
rect 7820 3800 7840 3820
rect 7820 3750 7840 3770
rect 7820 3700 7840 3720
rect 7820 3650 7840 3670
rect 7930 3800 7950 3820
rect 7930 3750 7950 3770
rect 7930 3700 7950 3720
rect 7930 3650 7950 3670
rect 7985 3800 8005 3820
rect 7985 3750 8005 3770
rect 7985 3700 8005 3720
rect 7985 3650 8005 3670
rect 8205 3800 8225 3820
rect 8205 3750 8225 3770
rect 8205 3700 8225 3720
rect 8205 3650 8225 3670
rect 8270 3800 8290 3820
rect 8270 3750 8290 3770
rect 8270 3700 8290 3720
rect 8270 3650 8290 3670
rect 8400 3800 8420 3820
rect 8400 3750 8420 3770
rect 8400 3700 8420 3720
rect 8400 3650 8420 3670
rect 8465 3800 8485 3820
rect 8465 3750 8485 3770
rect 8465 3700 8485 3720
rect 8465 3650 8485 3670
rect 8595 3800 8615 3820
rect 8595 3750 8615 3770
rect 8595 3700 8615 3720
rect 8595 3650 8615 3670
rect 8660 3800 8680 3820
rect 8660 3750 8680 3770
rect 8660 3700 8680 3720
rect 8660 3650 8680 3670
rect 8740 3800 8760 3820
rect 8740 3750 8760 3770
rect 8740 3700 8760 3720
rect 8740 3650 8760 3670
rect 8805 3800 8825 3820
rect 8805 3750 8825 3770
rect 8805 3700 8825 3720
rect 8805 3650 8825 3670
rect 6635 3420 6655 3440
rect 6635 3370 6655 3390
rect 6635 3320 6655 3340
rect 6635 3270 6655 3290
rect 6690 3420 6710 3440
rect 6690 3370 6710 3390
rect 6690 3320 6710 3340
rect 6690 3270 6710 3290
rect 6745 3420 6765 3440
rect 6745 3370 6765 3390
rect 6745 3320 6765 3340
rect 6745 3270 6765 3290
rect 6895 3420 6915 3440
rect 6895 3370 6915 3390
rect 6895 3320 6915 3340
rect 6895 3270 6915 3290
rect 6950 3420 6970 3440
rect 6950 3370 6970 3390
rect 6950 3320 6970 3340
rect 6950 3270 6970 3290
rect 7005 3420 7025 3440
rect 7085 3420 7105 3440
rect 7005 3370 7025 3390
rect 7085 3370 7105 3390
rect 7005 3320 7025 3340
rect 7085 3320 7105 3340
rect 7005 3270 7025 3290
rect 7085 3270 7105 3290
rect 7140 3420 7160 3440
rect 7140 3370 7160 3390
rect 7140 3320 7160 3340
rect 7140 3270 7160 3290
rect 7195 3420 7215 3440
rect 7195 3370 7215 3390
rect 7195 3320 7215 3340
rect 7195 3270 7215 3290
rect 7345 3420 7365 3440
rect 7345 3370 7365 3390
rect 7345 3320 7365 3340
rect 7345 3270 7365 3290
rect 7400 3420 7420 3440
rect 7400 3370 7420 3390
rect 7400 3320 7420 3340
rect 7400 3270 7420 3290
rect 7455 3420 7475 3440
rect 7455 3370 7475 3390
rect 7455 3320 7475 3340
rect 7455 3270 7475 3290
rect 7605 3420 7625 3440
rect 7605 3370 7625 3390
rect 7605 3320 7625 3340
rect 7605 3270 7625 3290
rect 7660 3420 7680 3440
rect 7660 3370 7680 3390
rect 7660 3320 7680 3340
rect 7660 3270 7680 3290
rect 7715 3420 7735 3440
rect 7715 3370 7735 3390
rect 7715 3320 7735 3340
rect 7715 3270 7735 3290
rect 7825 3420 7845 3440
rect 7825 3370 7845 3390
rect 7825 3320 7845 3340
rect 7825 3270 7845 3290
rect 7880 3420 7900 3440
rect 7880 3370 7900 3390
rect 7880 3320 7900 3340
rect 7880 3270 7900 3290
rect 7990 3420 8010 3440
rect 7990 3370 8010 3390
rect 7990 3320 8010 3340
rect 7990 3270 8010 3290
rect 8045 3420 8065 3440
rect 8045 3370 8065 3390
rect 8045 3320 8065 3340
rect 8045 3270 8065 3290
rect 8205 3420 8225 3440
rect 8205 3370 8225 3390
rect 8205 3320 8225 3340
rect 8205 3270 8225 3290
rect 8270 3420 8290 3440
rect 8270 3370 8290 3390
rect 8270 3320 8290 3340
rect 8270 3270 8290 3290
rect 8400 3420 8420 3440
rect 8400 3370 8420 3390
rect 8400 3320 8420 3340
rect 8400 3270 8420 3290
rect 8465 3420 8485 3440
rect 8465 3370 8485 3390
rect 8465 3320 8485 3340
rect 8465 3270 8485 3290
rect 8595 3420 8615 3440
rect 8595 3370 8615 3390
rect 8595 3320 8615 3340
rect 8595 3270 8615 3290
rect 8660 3420 8680 3440
rect 8660 3370 8680 3390
rect 8660 3320 8680 3340
rect 8660 3270 8680 3290
rect 8740 3420 8760 3440
rect 8740 3370 8760 3390
rect 8740 3320 8760 3340
rect 8740 3270 8760 3290
rect 8805 3420 8825 3440
rect 8805 3370 8825 3390
rect 8805 3320 8825 3340
rect 8805 3270 8825 3290
rect 8935 3420 8955 3440
rect 8935 3370 8955 3390
rect 8935 3320 8955 3340
rect 8935 3270 8955 3290
rect 9000 3420 9020 3440
rect 9000 3370 9020 3390
rect 9000 3320 9020 3340
rect 9000 3270 9020 3290
rect 9780 3435 9800 3455
rect 9780 3385 9800 3405
rect 9780 3335 9800 3355
rect 9780 3285 9800 3305
rect 9890 3435 9910 3455
rect 9890 3385 9910 3405
rect 9890 3335 9910 3355
rect 9890 3285 9910 3305
rect 10000 3435 10020 3455
rect 10000 3385 10020 3405
rect 10000 3335 10020 3355
rect 10000 3285 10020 3305
rect 10110 3435 10130 3455
rect 10110 3385 10130 3405
rect 10110 3335 10130 3355
rect 10110 3285 10130 3305
rect 10220 3435 10240 3455
rect 10220 3385 10240 3405
rect 10220 3335 10240 3355
rect 10220 3285 10240 3305
rect 10330 3435 10350 3455
rect 10330 3385 10350 3405
rect 10330 3335 10350 3355
rect 10330 3285 10350 3305
rect 10440 3435 10460 3455
rect 10540 3435 10560 3455
rect 10440 3385 10460 3405
rect 10540 3385 10560 3405
rect 10440 3335 10460 3355
rect 10540 3335 10560 3355
rect 10440 3285 10460 3305
rect 10540 3285 10560 3305
rect 10650 3435 10670 3455
rect 10650 3385 10670 3405
rect 10650 3335 10670 3355
rect 10650 3285 10670 3305
rect 10760 3435 10780 3455
rect 10760 3385 10780 3405
rect 10760 3335 10780 3355
rect 10760 3285 10780 3305
rect 10870 3435 10890 3455
rect 10870 3385 10890 3405
rect 10870 3335 10890 3355
rect 10870 3285 10890 3305
rect 10980 3435 11000 3455
rect 10980 3385 11000 3405
rect 10980 3335 11000 3355
rect 10980 3285 11000 3305
rect 11090 3435 11110 3455
rect 11090 3385 11110 3405
rect 11090 3335 11110 3355
rect 11090 3285 11110 3305
rect 11200 3435 11220 3455
rect 11200 3385 11220 3405
rect 11200 3335 11220 3355
rect 11200 3285 11220 3305
<< psubdiff >>
rect 6585 4030 6625 4045
rect 6585 4010 6595 4030
rect 6615 4010 6625 4030
rect 6585 3980 6625 4010
rect 6585 3960 6595 3980
rect 6615 3960 6625 3980
rect 6585 3945 6625 3960
rect 7035 4030 7075 4045
rect 7035 4010 7045 4030
rect 7065 4010 7075 4030
rect 7035 3980 7075 4010
rect 7035 3960 7045 3980
rect 7065 3960 7075 3980
rect 7035 3945 7075 3960
rect 7485 4030 7525 4045
rect 7485 4010 7495 4030
rect 7515 4010 7525 4030
rect 7485 3980 7525 4010
rect 7485 3960 7495 3980
rect 7515 3960 7525 3980
rect 7485 3945 7525 3960
rect 7685 4030 7725 4045
rect 7685 4010 7695 4030
rect 7715 4010 7725 4030
rect 7685 3980 7725 4010
rect 7685 3960 7695 3980
rect 7715 3960 7725 3980
rect 7685 3945 7725 3960
rect 7850 4030 7890 4045
rect 7850 4010 7860 4030
rect 7880 4010 7890 4030
rect 7850 3980 7890 4010
rect 7850 3960 7860 3980
rect 7880 3960 7890 3980
rect 7850 3945 7890 3960
rect 8015 4030 8055 4045
rect 8015 4010 8025 4030
rect 8045 4010 8055 4030
rect 8015 3980 8055 4010
rect 8015 3960 8025 3980
rect 8045 3960 8055 3980
rect 8015 3945 8055 3960
rect 8140 4030 8190 4045
rect 8140 4010 8155 4030
rect 8175 4010 8190 4030
rect 8140 3980 8190 4010
rect 8140 3960 8155 3980
rect 8175 3960 8190 3980
rect 8140 3945 8190 3960
rect 8530 4030 8580 4045
rect 8530 4010 8545 4030
rect 8565 4010 8580 4030
rect 8530 3980 8580 4010
rect 8530 3960 8545 3980
rect 8565 3960 8580 3980
rect 8530 3945 8580 3960
rect 8870 4030 8920 4045
rect 8870 4010 8885 4030
rect 8905 4010 8920 4030
rect 8870 3980 8920 4010
rect 8870 3960 8885 3980
rect 8905 3960 8920 3980
rect 8870 3945 8920 3960
rect 9615 4005 9665 4020
rect 9615 3985 9630 4005
rect 9650 3985 9665 4005
rect 9615 3955 9665 3985
rect 9615 3935 9630 3955
rect 9650 3935 9665 3955
rect 9615 3905 9665 3935
rect 9615 3885 9630 3905
rect 9650 3885 9665 3905
rect 9615 3855 9665 3885
rect 9615 3835 9630 3855
rect 9650 3835 9665 3855
rect 9615 3820 9665 3835
rect 10155 4005 10205 4020
rect 10155 3985 10170 4005
rect 10190 3985 10205 4005
rect 10155 3955 10205 3985
rect 10155 3935 10170 3955
rect 10190 3935 10205 3955
rect 10155 3905 10205 3935
rect 10155 3885 10170 3905
rect 10190 3885 10205 3905
rect 10155 3855 10205 3885
rect 10155 3835 10170 3855
rect 10190 3835 10205 3855
rect 10155 3820 10205 3835
rect 10695 4005 10745 4020
rect 10695 3985 10710 4005
rect 10730 3985 10745 4005
rect 10695 3955 10745 3985
rect 10695 3935 10710 3955
rect 10730 3935 10745 3955
rect 10695 3905 10745 3935
rect 10695 3885 10710 3905
rect 10730 3885 10745 3905
rect 10695 3855 10745 3885
rect 10695 3835 10710 3855
rect 10730 3835 10745 3855
rect 10695 3820 10745 3835
rect 11235 4005 11285 4020
rect 11235 3985 11250 4005
rect 11270 3985 11285 4005
rect 11235 3955 11285 3985
rect 11235 3935 11250 3955
rect 11270 3935 11285 3955
rect 11235 3905 11285 3935
rect 11235 3885 11250 3905
rect 11270 3885 11285 3905
rect 11235 3855 11285 3885
rect 11235 3835 11250 3855
rect 11270 3835 11285 3855
rect 11235 3820 11285 3835
rect 6585 3130 6625 3145
rect 6585 3110 6595 3130
rect 6615 3110 6625 3130
rect 6585 3080 6625 3110
rect 6585 3060 6595 3080
rect 6615 3060 6625 3080
rect 6585 3045 6625 3060
rect 7035 3130 7075 3145
rect 7035 3110 7045 3130
rect 7065 3110 7075 3130
rect 7035 3080 7075 3110
rect 7035 3060 7045 3080
rect 7065 3060 7075 3080
rect 7035 3045 7075 3060
rect 7485 3130 7525 3145
rect 7485 3110 7495 3130
rect 7515 3110 7525 3130
rect 7485 3080 7525 3110
rect 7485 3060 7495 3080
rect 7515 3060 7525 3080
rect 7485 3045 7525 3060
rect 7555 3130 7595 3145
rect 7555 3110 7565 3130
rect 7585 3110 7595 3130
rect 7555 3080 7595 3110
rect 7555 3060 7565 3080
rect 7585 3060 7595 3080
rect 7555 3045 7595 3060
rect 7775 3130 7815 3145
rect 7775 3110 7785 3130
rect 7805 3110 7815 3130
rect 7775 3080 7815 3110
rect 7775 3060 7785 3080
rect 7805 3060 7815 3080
rect 7775 3045 7815 3060
rect 7940 3130 7980 3145
rect 7940 3110 7950 3130
rect 7970 3110 7980 3130
rect 7940 3080 7980 3110
rect 7940 3060 7950 3080
rect 7970 3060 7980 3080
rect 7940 3045 7980 3060
rect 8150 3130 8190 3145
rect 8150 3110 8160 3130
rect 8180 3110 8190 3130
rect 8150 3080 8190 3110
rect 8150 3060 8160 3080
rect 8180 3060 8190 3080
rect 8150 3045 8190 3060
rect 8345 3130 8385 3145
rect 8345 3110 8355 3130
rect 8375 3110 8385 3130
rect 8345 3080 8385 3110
rect 8345 3060 8355 3080
rect 8375 3060 8385 3080
rect 8345 3045 8385 3060
rect 8540 3130 8580 3145
rect 8540 3110 8550 3130
rect 8570 3110 8580 3130
rect 8540 3080 8580 3110
rect 8540 3060 8550 3080
rect 8570 3060 8580 3080
rect 8540 3045 8580 3060
<< nsubdiff >>
rect 6585 3820 6625 3835
rect 6585 3800 6595 3820
rect 6615 3800 6625 3820
rect 6585 3770 6625 3800
rect 6585 3750 6595 3770
rect 6615 3750 6625 3770
rect 6585 3720 6625 3750
rect 6585 3700 6595 3720
rect 6615 3700 6625 3720
rect 6585 3670 6625 3700
rect 6585 3650 6595 3670
rect 6615 3650 6625 3670
rect 6585 3635 6625 3650
rect 7035 3820 7075 3835
rect 7035 3800 7045 3820
rect 7065 3800 7075 3820
rect 7035 3770 7075 3800
rect 7035 3750 7045 3770
rect 7065 3750 7075 3770
rect 7035 3720 7075 3750
rect 7035 3700 7045 3720
rect 7065 3700 7075 3720
rect 7035 3670 7075 3700
rect 7035 3650 7045 3670
rect 7065 3650 7075 3670
rect 7035 3635 7075 3650
rect 7485 3820 7525 3835
rect 7485 3800 7495 3820
rect 7515 3800 7525 3820
rect 7485 3770 7525 3800
rect 7485 3750 7495 3770
rect 7515 3750 7525 3770
rect 7485 3720 7525 3750
rect 7485 3700 7495 3720
rect 7515 3700 7525 3720
rect 7485 3670 7525 3700
rect 7485 3650 7495 3670
rect 7515 3650 7525 3670
rect 7485 3635 7525 3650
rect 7685 3820 7725 3835
rect 7685 3800 7695 3820
rect 7715 3800 7725 3820
rect 7685 3770 7725 3800
rect 7685 3750 7695 3770
rect 7715 3750 7725 3770
rect 7685 3720 7725 3750
rect 7685 3700 7695 3720
rect 7715 3700 7725 3720
rect 7685 3670 7725 3700
rect 7685 3650 7695 3670
rect 7715 3650 7725 3670
rect 7685 3635 7725 3650
rect 7850 3820 7890 3835
rect 7850 3800 7860 3820
rect 7880 3800 7890 3820
rect 7850 3770 7890 3800
rect 7850 3750 7860 3770
rect 7880 3750 7890 3770
rect 7850 3720 7890 3750
rect 7850 3700 7860 3720
rect 7880 3700 7890 3720
rect 7850 3670 7890 3700
rect 7850 3650 7860 3670
rect 7880 3650 7890 3670
rect 7850 3635 7890 3650
rect 8015 3820 8055 3835
rect 8015 3800 8025 3820
rect 8045 3800 8055 3820
rect 8015 3770 8055 3800
rect 8015 3750 8025 3770
rect 8045 3750 8055 3770
rect 8015 3720 8055 3750
rect 8015 3700 8025 3720
rect 8045 3700 8055 3720
rect 8015 3670 8055 3700
rect 8015 3650 8025 3670
rect 8045 3650 8055 3670
rect 8015 3635 8055 3650
rect 8140 3820 8190 3835
rect 8140 3800 8155 3820
rect 8175 3800 8190 3820
rect 8140 3770 8190 3800
rect 8140 3750 8155 3770
rect 8175 3750 8190 3770
rect 8140 3720 8190 3750
rect 8140 3700 8155 3720
rect 8175 3700 8190 3720
rect 8140 3670 8190 3700
rect 8140 3650 8155 3670
rect 8175 3650 8190 3670
rect 8140 3635 8190 3650
rect 8530 3820 8580 3835
rect 8530 3800 8545 3820
rect 8565 3800 8580 3820
rect 8530 3770 8580 3800
rect 8530 3750 8545 3770
rect 8565 3750 8580 3770
rect 8530 3720 8580 3750
rect 8530 3700 8545 3720
rect 8565 3700 8580 3720
rect 8530 3670 8580 3700
rect 8530 3650 8545 3670
rect 8565 3650 8580 3670
rect 8530 3635 8580 3650
rect 9715 3455 9765 3470
rect 6585 3440 6625 3455
rect 6585 3420 6595 3440
rect 6615 3420 6625 3440
rect 6585 3390 6625 3420
rect 6585 3370 6595 3390
rect 6615 3370 6625 3390
rect 6585 3340 6625 3370
rect 6585 3320 6595 3340
rect 6615 3320 6625 3340
rect 6585 3290 6625 3320
rect 6585 3270 6595 3290
rect 6615 3270 6625 3290
rect 6585 3255 6625 3270
rect 7035 3440 7075 3455
rect 7035 3420 7045 3440
rect 7065 3420 7075 3440
rect 7035 3390 7075 3420
rect 7035 3370 7045 3390
rect 7065 3370 7075 3390
rect 7035 3340 7075 3370
rect 7035 3320 7045 3340
rect 7065 3320 7075 3340
rect 7035 3290 7075 3320
rect 7035 3270 7045 3290
rect 7065 3270 7075 3290
rect 7035 3255 7075 3270
rect 7485 3440 7525 3455
rect 7485 3420 7495 3440
rect 7515 3420 7525 3440
rect 7485 3390 7525 3420
rect 7485 3370 7495 3390
rect 7515 3370 7525 3390
rect 7485 3340 7525 3370
rect 7485 3320 7495 3340
rect 7515 3320 7525 3340
rect 7485 3290 7525 3320
rect 7485 3270 7495 3290
rect 7515 3270 7525 3290
rect 7485 3255 7525 3270
rect 7555 3440 7595 3455
rect 7555 3420 7565 3440
rect 7585 3420 7595 3440
rect 7555 3390 7595 3420
rect 7555 3370 7565 3390
rect 7585 3370 7595 3390
rect 7555 3340 7595 3370
rect 7555 3320 7565 3340
rect 7585 3320 7595 3340
rect 7555 3290 7595 3320
rect 7555 3270 7565 3290
rect 7585 3270 7595 3290
rect 7555 3255 7595 3270
rect 7775 3440 7815 3455
rect 7775 3420 7785 3440
rect 7805 3420 7815 3440
rect 7775 3390 7815 3420
rect 7775 3370 7785 3390
rect 7805 3370 7815 3390
rect 7775 3340 7815 3370
rect 7775 3320 7785 3340
rect 7805 3320 7815 3340
rect 7775 3290 7815 3320
rect 7775 3270 7785 3290
rect 7805 3270 7815 3290
rect 7775 3255 7815 3270
rect 7940 3440 7980 3455
rect 7940 3420 7950 3440
rect 7970 3420 7980 3440
rect 7940 3390 7980 3420
rect 7940 3370 7950 3390
rect 7970 3370 7980 3390
rect 7940 3340 7980 3370
rect 7940 3320 7950 3340
rect 7970 3320 7980 3340
rect 7940 3290 7980 3320
rect 7940 3270 7950 3290
rect 7970 3270 7980 3290
rect 7940 3255 7980 3270
rect 8140 3440 8190 3455
rect 8140 3420 8155 3440
rect 8175 3420 8190 3440
rect 8140 3390 8190 3420
rect 8140 3370 8155 3390
rect 8175 3370 8190 3390
rect 8140 3340 8190 3370
rect 8140 3320 8155 3340
rect 8175 3320 8190 3340
rect 8140 3290 8190 3320
rect 8140 3270 8155 3290
rect 8175 3270 8190 3290
rect 8140 3255 8190 3270
rect 8335 3440 8385 3455
rect 8335 3420 8350 3440
rect 8370 3420 8385 3440
rect 8335 3390 8385 3420
rect 8335 3370 8350 3390
rect 8370 3370 8385 3390
rect 8335 3340 8385 3370
rect 8335 3320 8350 3340
rect 8370 3320 8385 3340
rect 8335 3290 8385 3320
rect 8335 3270 8350 3290
rect 8370 3270 8385 3290
rect 8335 3255 8385 3270
rect 8530 3440 8580 3455
rect 8530 3420 8545 3440
rect 8565 3420 8580 3440
rect 8530 3390 8580 3420
rect 8530 3370 8545 3390
rect 8565 3370 8580 3390
rect 8530 3340 8580 3370
rect 8530 3320 8545 3340
rect 8565 3320 8580 3340
rect 8530 3290 8580 3320
rect 8530 3270 8545 3290
rect 8565 3270 8580 3290
rect 8530 3255 8580 3270
rect 8870 3440 8920 3455
rect 8870 3420 8885 3440
rect 8905 3420 8920 3440
rect 8870 3390 8920 3420
rect 8870 3370 8885 3390
rect 8905 3370 8920 3390
rect 8870 3340 8920 3370
rect 8870 3320 8885 3340
rect 8905 3320 8920 3340
rect 8870 3290 8920 3320
rect 8870 3270 8885 3290
rect 8905 3270 8920 3290
rect 8870 3255 8920 3270
rect 9715 3435 9730 3455
rect 9750 3435 9765 3455
rect 9715 3405 9765 3435
rect 9715 3385 9730 3405
rect 9750 3385 9765 3405
rect 9715 3355 9765 3385
rect 9715 3335 9730 3355
rect 9750 3335 9765 3355
rect 9715 3305 9765 3335
rect 9715 3285 9730 3305
rect 9750 3285 9765 3305
rect 9715 3270 9765 3285
rect 10475 3455 10525 3470
rect 10475 3435 10490 3455
rect 10510 3435 10525 3455
rect 10475 3405 10525 3435
rect 10475 3385 10490 3405
rect 10510 3385 10525 3405
rect 10475 3355 10525 3385
rect 10475 3335 10490 3355
rect 10510 3335 10525 3355
rect 10475 3305 10525 3335
rect 10475 3285 10490 3305
rect 10510 3285 10525 3305
rect 10475 3270 10525 3285
rect 11235 3455 11285 3470
rect 11235 3435 11250 3455
rect 11270 3435 11285 3455
rect 11235 3405 11285 3435
rect 11235 3385 11250 3405
rect 11270 3385 11285 3405
rect 11235 3355 11285 3385
rect 11235 3335 11250 3355
rect 11270 3335 11285 3355
rect 11235 3305 11285 3335
rect 11235 3285 11250 3305
rect 11270 3285 11285 3305
rect 11235 3270 11285 3285
<< psubdiffcont >>
rect 6595 4010 6615 4030
rect 6595 3960 6615 3980
rect 7045 4010 7065 4030
rect 7045 3960 7065 3980
rect 7495 4010 7515 4030
rect 7495 3960 7515 3980
rect 7695 4010 7715 4030
rect 7695 3960 7715 3980
rect 7860 4010 7880 4030
rect 7860 3960 7880 3980
rect 8025 4010 8045 4030
rect 8025 3960 8045 3980
rect 8155 4010 8175 4030
rect 8155 3960 8175 3980
rect 8545 4010 8565 4030
rect 8545 3960 8565 3980
rect 8885 4010 8905 4030
rect 8885 3960 8905 3980
rect 9630 3985 9650 4005
rect 9630 3935 9650 3955
rect 9630 3885 9650 3905
rect 9630 3835 9650 3855
rect 10170 3985 10190 4005
rect 10170 3935 10190 3955
rect 10170 3885 10190 3905
rect 10170 3835 10190 3855
rect 10710 3985 10730 4005
rect 10710 3935 10730 3955
rect 10710 3885 10730 3905
rect 10710 3835 10730 3855
rect 11250 3985 11270 4005
rect 11250 3935 11270 3955
rect 11250 3885 11270 3905
rect 11250 3835 11270 3855
rect 6595 3110 6615 3130
rect 6595 3060 6615 3080
rect 7045 3110 7065 3130
rect 7045 3060 7065 3080
rect 7495 3110 7515 3130
rect 7495 3060 7515 3080
rect 7565 3110 7585 3130
rect 7565 3060 7585 3080
rect 7785 3110 7805 3130
rect 7785 3060 7805 3080
rect 7950 3110 7970 3130
rect 7950 3060 7970 3080
rect 8160 3110 8180 3130
rect 8160 3060 8180 3080
rect 8355 3110 8375 3130
rect 8355 3060 8375 3080
rect 8550 3110 8570 3130
rect 8550 3060 8570 3080
<< nsubdiffcont >>
rect 6595 3800 6615 3820
rect 6595 3750 6615 3770
rect 6595 3700 6615 3720
rect 6595 3650 6615 3670
rect 7045 3800 7065 3820
rect 7045 3750 7065 3770
rect 7045 3700 7065 3720
rect 7045 3650 7065 3670
rect 7495 3800 7515 3820
rect 7495 3750 7515 3770
rect 7495 3700 7515 3720
rect 7495 3650 7515 3670
rect 7695 3800 7715 3820
rect 7695 3750 7715 3770
rect 7695 3700 7715 3720
rect 7695 3650 7715 3670
rect 7860 3800 7880 3820
rect 7860 3750 7880 3770
rect 7860 3700 7880 3720
rect 7860 3650 7880 3670
rect 8025 3800 8045 3820
rect 8025 3750 8045 3770
rect 8025 3700 8045 3720
rect 8025 3650 8045 3670
rect 8155 3800 8175 3820
rect 8155 3750 8175 3770
rect 8155 3700 8175 3720
rect 8155 3650 8175 3670
rect 8545 3800 8565 3820
rect 8545 3750 8565 3770
rect 8545 3700 8565 3720
rect 8545 3650 8565 3670
rect 6595 3420 6615 3440
rect 6595 3370 6615 3390
rect 6595 3320 6615 3340
rect 6595 3270 6615 3290
rect 7045 3420 7065 3440
rect 7045 3370 7065 3390
rect 7045 3320 7065 3340
rect 7045 3270 7065 3290
rect 7495 3420 7515 3440
rect 7495 3370 7515 3390
rect 7495 3320 7515 3340
rect 7495 3270 7515 3290
rect 7565 3420 7585 3440
rect 7565 3370 7585 3390
rect 7565 3320 7585 3340
rect 7565 3270 7585 3290
rect 7785 3420 7805 3440
rect 7785 3370 7805 3390
rect 7785 3320 7805 3340
rect 7785 3270 7805 3290
rect 7950 3420 7970 3440
rect 7950 3370 7970 3390
rect 7950 3320 7970 3340
rect 7950 3270 7970 3290
rect 8155 3420 8175 3440
rect 8155 3370 8175 3390
rect 8155 3320 8175 3340
rect 8155 3270 8175 3290
rect 8350 3420 8370 3440
rect 8350 3370 8370 3390
rect 8350 3320 8370 3340
rect 8350 3270 8370 3290
rect 8545 3420 8565 3440
rect 8545 3370 8565 3390
rect 8545 3320 8565 3340
rect 8545 3270 8565 3290
rect 8885 3420 8905 3440
rect 8885 3370 8905 3390
rect 8885 3320 8905 3340
rect 8885 3270 8905 3290
rect 9730 3435 9750 3455
rect 9730 3385 9750 3405
rect 9730 3335 9750 3355
rect 9730 3285 9750 3305
rect 10490 3435 10510 3455
rect 10490 3385 10510 3405
rect 10490 3335 10510 3355
rect 10490 3285 10510 3305
rect 11250 3435 11270 3455
rect 11250 3385 11270 3405
rect 11250 3335 11270 3355
rect 11250 3285 11270 3305
<< poly >>
rect 6925 4085 7130 4100
rect 6665 4045 6680 4060
rect 6720 4045 6735 4060
rect 6925 4045 6940 4085
rect 6980 4045 6995 4060
rect 7115 4045 7130 4085
rect 8435 4090 8490 4100
rect 8435 4070 8460 4090
rect 8480 4070 8490 4090
rect 8435 4060 8490 4070
rect 8765 4090 8805 4100
rect 8765 4070 8775 4090
rect 8795 4070 8805 4090
rect 8765 4060 8805 4070
rect 9670 4065 9710 4075
rect 7170 4045 7185 4060
rect 7375 4045 7390 4060
rect 7430 4045 7445 4060
rect 7630 4045 7645 4060
rect 7795 4045 7810 4060
rect 7960 4045 7975 4060
rect 8240 4045 8255 4060
rect 8435 4045 8450 4060
rect 8630 4045 8645 4060
rect 8775 4045 8790 4060
rect 8970 4045 8985 4060
rect 9670 4045 9680 4065
rect 9700 4050 9710 4065
rect 9935 4060 10425 4075
rect 9935 4050 9995 4060
rect 9700 4045 9775 4050
rect 9670 4035 9775 4045
rect 9715 4020 9775 4035
rect 9825 4030 9995 4050
rect 10365 4050 10425 4060
rect 11190 4065 11230 4075
rect 11190 4050 11200 4065
rect 9825 4020 9885 4030
rect 9935 4020 9995 4030
rect 10045 4020 10105 4035
rect 10255 4020 10315 4035
rect 10365 4030 10535 4050
rect 10365 4020 10425 4030
rect 10475 4020 10535 4030
rect 10585 4020 10645 4035
rect 10795 4020 10855 4035
rect 10905 4030 11075 4050
rect 10905 4020 10965 4030
rect 11015 4020 11075 4030
rect 11125 4045 11200 4050
rect 11220 4045 11230 4065
rect 11125 4035 11230 4045
rect 11125 4020 11185 4035
rect 6665 3910 6680 3945
rect 6565 3900 6680 3910
rect 6565 3880 6575 3900
rect 6595 3895 6680 3900
rect 6595 3880 6605 3895
rect 6565 3870 6605 3880
rect 6665 3835 6680 3895
rect 6720 3930 6735 3945
rect 6720 3920 6770 3930
rect 6925 3925 6940 3945
rect 6720 3900 6740 3920
rect 6760 3900 6770 3920
rect 6720 3890 6770 3900
rect 6815 3910 6940 3925
rect 6720 3835 6735 3890
rect 6815 3680 6830 3910
rect 6925 3835 6940 3910
rect 6980 3890 6995 3945
rect 6980 3880 7030 3890
rect 6980 3860 7000 3880
rect 7020 3860 7030 3880
rect 6980 3850 7030 3860
rect 6980 3835 6995 3850
rect 7115 3835 7130 3945
rect 7170 3930 7185 3945
rect 7170 3920 7220 3930
rect 7375 3925 7390 3945
rect 7170 3900 7190 3920
rect 7210 3900 7220 3920
rect 7170 3890 7220 3900
rect 7265 3910 7390 3925
rect 7170 3835 7185 3890
rect 6790 3670 6830 3680
rect 6790 3650 6800 3670
rect 6820 3650 6830 3670
rect 6790 3640 6830 3650
rect 7265 3680 7280 3910
rect 7375 3835 7390 3910
rect 7430 3880 7445 3945
rect 7525 3895 7605 3905
rect 7525 3880 7535 3895
rect 7430 3875 7535 3880
rect 7555 3875 7575 3895
rect 7595 3875 7605 3895
rect 7430 3865 7605 3875
rect 7630 3895 7645 3945
rect 7730 3895 7770 3905
rect 7630 3880 7740 3895
rect 7430 3835 7445 3865
rect 7630 3835 7645 3880
rect 7730 3875 7740 3880
rect 7760 3875 7770 3895
rect 7730 3865 7770 3875
rect 7795 3895 7810 3945
rect 7895 3895 7935 3905
rect 7795 3880 7905 3895
rect 7795 3835 7810 3880
rect 7895 3875 7905 3880
rect 7925 3875 7935 3895
rect 7895 3865 7935 3875
rect 7960 3895 7975 3945
rect 8240 3910 8255 3945
rect 8435 3930 8450 3945
rect 8040 3895 8080 3905
rect 7960 3880 8050 3895
rect 7960 3835 7975 3880
rect 8040 3875 8050 3880
rect 8070 3875 8080 3895
rect 8040 3865 8080 3875
rect 8115 3900 8255 3910
rect 8115 3880 8125 3900
rect 8145 3895 8255 3900
rect 8145 3880 8155 3895
rect 8115 3870 8155 3880
rect 8240 3835 8255 3895
rect 8475 3885 8515 3895
rect 8475 3865 8485 3885
rect 8505 3870 8515 3885
rect 8630 3870 8645 3945
rect 8775 3935 8790 3945
rect 8670 3925 8790 3935
rect 8670 3905 8680 3925
rect 8700 3920 8790 3925
rect 8700 3905 8710 3920
rect 8670 3900 8710 3905
rect 8970 3870 8985 3945
rect 8505 3865 8985 3870
rect 8475 3855 8985 3865
rect 8435 3835 8450 3850
rect 8630 3835 8645 3855
rect 8775 3835 8790 3855
rect 7240 3670 7280 3680
rect 7240 3650 7250 3670
rect 7270 3650 7280 3670
rect 7240 3640 7280 3650
rect 9715 3805 9775 3820
rect 9825 3810 9885 3820
rect 9935 3810 9995 3820
rect 9825 3800 9995 3810
rect 9825 3795 9900 3800
rect 9890 3780 9900 3795
rect 9920 3795 9995 3800
rect 10045 3810 10105 3820
rect 10255 3810 10315 3820
rect 10045 3795 10315 3810
rect 10365 3810 10425 3820
rect 10475 3810 10535 3820
rect 10365 3795 10535 3810
rect 10585 3810 10645 3820
rect 10795 3810 10855 3820
rect 10585 3795 10855 3810
rect 10905 3805 10965 3820
rect 11015 3805 11075 3820
rect 11125 3805 11185 3820
rect 9920 3780 9930 3795
rect 9890 3770 9930 3780
rect 10160 3775 10170 3795
rect 10190 3775 10200 3795
rect 10160 3765 10200 3775
rect 10700 3775 10710 3795
rect 10730 3775 10740 3795
rect 10700 3765 10740 3775
rect 10905 3790 11075 3805
rect 10905 3780 10945 3790
rect 10905 3760 10915 3780
rect 10935 3760 10945 3780
rect 10905 3750 10945 3760
rect 11035 3780 11075 3790
rect 11035 3760 11045 3780
rect 11065 3760 11075 3780
rect 11035 3750 11075 3760
rect 6665 3620 6680 3635
rect 6720 3620 6735 3635
rect 6925 3620 6940 3635
rect 6980 3620 6995 3635
rect 7115 3620 7130 3635
rect 7170 3620 7185 3635
rect 7375 3620 7390 3635
rect 7430 3620 7445 3635
rect 7630 3620 7645 3635
rect 7795 3620 7810 3635
rect 7960 3620 7975 3635
rect 8240 3620 8255 3635
rect 8435 3620 8450 3635
rect 8630 3620 8645 3635
rect 8775 3620 8790 3635
rect 6850 3610 6890 3620
rect 6850 3590 6860 3610
rect 6880 3590 6890 3610
rect 6850 3580 6890 3590
rect 8410 3610 8450 3620
rect 8410 3590 8420 3610
rect 8440 3590 8450 3610
rect 8410 3585 8450 3590
rect 10685 3530 10725 3540
rect 10100 3515 10140 3525
rect 7625 3500 7665 3505
rect 10100 3500 10110 3515
rect 7625 3480 7635 3500
rect 7655 3480 7665 3500
rect 9925 3495 10110 3500
rect 10130 3500 10140 3515
rect 10480 3515 10520 3525
rect 10130 3495 10315 3500
rect 10480 3495 10490 3515
rect 10510 3495 10520 3515
rect 10685 3510 10695 3530
rect 10715 3510 10725 3530
rect 10685 3500 10725 3510
rect 11035 3530 11075 3540
rect 11035 3510 11045 3530
rect 11065 3510 11075 3530
rect 11035 3500 11075 3510
rect 7625 3470 7665 3480
rect 9815 3470 9875 3485
rect 9925 3480 10315 3495
rect 9925 3470 9985 3480
rect 10035 3470 10095 3480
rect 10145 3470 10205 3480
rect 10255 3470 10315 3480
rect 10365 3480 10635 3495
rect 10365 3470 10425 3480
rect 10575 3470 10635 3480
rect 10685 3485 11075 3500
rect 10685 3470 10745 3485
rect 10795 3470 10855 3485
rect 10905 3470 10965 3485
rect 11015 3470 11075 3485
rect 11125 3470 11185 3485
rect 6665 3455 6680 3470
rect 6720 3455 6735 3470
rect 6925 3455 6940 3470
rect 6980 3455 6995 3470
rect 7115 3455 7130 3470
rect 7170 3455 7185 3470
rect 7375 3455 7390 3470
rect 7430 3455 7445 3470
rect 7635 3455 7650 3470
rect 7690 3455 7705 3470
rect 7855 3455 7870 3470
rect 8020 3455 8035 3470
rect 8240 3455 8255 3470
rect 8435 3455 8450 3470
rect 8630 3455 8645 3470
rect 8775 3455 8790 3470
rect 8970 3455 8985 3470
rect 6790 3440 6830 3450
rect 6790 3420 6800 3440
rect 6820 3420 6830 3440
rect 6790 3410 6830 3420
rect 6565 3210 6605 3220
rect 6565 3190 6575 3210
rect 6595 3195 6605 3210
rect 6665 3195 6680 3255
rect 6595 3190 6680 3195
rect 6565 3180 6680 3190
rect 6665 3145 6680 3180
rect 6720 3200 6735 3255
rect 6720 3190 6770 3200
rect 6720 3170 6740 3190
rect 6760 3170 6770 3190
rect 6720 3160 6770 3170
rect 6815 3180 6830 3410
rect 7240 3440 7280 3450
rect 7240 3420 7250 3440
rect 7270 3420 7280 3440
rect 7240 3410 7280 3420
rect 6925 3180 6940 3255
rect 6815 3165 6940 3180
rect 6720 3145 6735 3160
rect 6925 3145 6940 3165
rect 6980 3240 6995 3255
rect 6980 3230 7030 3240
rect 6980 3210 7000 3230
rect 7020 3210 7030 3230
rect 6980 3200 7030 3210
rect 6980 3145 6995 3200
rect 7115 3145 7130 3255
rect 7170 3200 7185 3255
rect 7170 3190 7220 3200
rect 7170 3170 7190 3190
rect 7210 3170 7220 3190
rect 7170 3160 7220 3170
rect 7265 3180 7280 3410
rect 9815 3255 9875 3270
rect 7375 3180 7390 3255
rect 7265 3165 7390 3180
rect 7170 3145 7185 3160
rect 7375 3145 7390 3165
rect 7430 3180 7445 3255
rect 7515 3195 7555 3205
rect 7515 3180 7525 3195
rect 7430 3175 7525 3180
rect 7545 3175 7555 3195
rect 7430 3165 7555 3175
rect 7430 3145 7445 3165
rect 7635 3145 7650 3255
rect 7690 3145 7705 3255
rect 7730 3215 7770 3225
rect 7730 3195 7740 3215
rect 7760 3210 7770 3215
rect 7855 3210 7870 3255
rect 7760 3195 7870 3210
rect 7730 3185 7770 3195
rect 7855 3145 7870 3195
rect 7895 3215 7935 3225
rect 7895 3195 7905 3215
rect 7925 3210 7935 3215
rect 8020 3210 8035 3255
rect 7925 3195 8035 3210
rect 7895 3185 7935 3195
rect 8020 3145 8035 3195
rect 8060 3215 8100 3225
rect 8060 3195 8070 3215
rect 8090 3195 8100 3215
rect 8240 3210 8255 3255
rect 8435 3225 8450 3255
rect 8060 3185 8100 3195
rect 8125 3200 8255 3210
rect 8125 3180 8135 3200
rect 8155 3195 8255 3200
rect 8155 3180 8165 3195
rect 8125 3170 8165 3180
rect 8240 3145 8255 3195
rect 8410 3215 8450 3225
rect 8410 3195 8420 3215
rect 8440 3195 8450 3215
rect 8630 3200 8645 3255
rect 8775 3240 8790 3255
rect 8670 3230 8885 3240
rect 8670 3210 8680 3230
rect 8700 3225 8855 3230
rect 8700 3210 8710 3225
rect 8670 3200 8710 3210
rect 8845 3210 8855 3225
rect 8875 3210 8885 3230
rect 8845 3200 8885 3210
rect 8410 3185 8450 3195
rect 8435 3145 8450 3185
rect 8605 3190 8645 3200
rect 8605 3170 8615 3190
rect 8635 3175 8645 3190
rect 8970 3175 8985 3255
rect 9770 3245 9875 3255
rect 9770 3225 9780 3245
rect 9800 3240 9875 3245
rect 9925 3260 9985 3270
rect 10035 3260 10095 3270
rect 10145 3260 10205 3270
rect 10255 3260 10315 3270
rect 9925 3240 10315 3260
rect 10365 3255 10425 3270
rect 10575 3255 10635 3270
rect 10685 3260 10745 3270
rect 10795 3260 10855 3270
rect 10905 3260 10965 3270
rect 11015 3260 11075 3270
rect 10685 3240 11075 3260
rect 11125 3255 11185 3270
rect 11125 3245 11230 3255
rect 11125 3240 11200 3245
rect 9800 3225 9810 3240
rect 9770 3215 9810 3225
rect 11190 3225 11200 3240
rect 11220 3225 11230 3245
rect 11190 3215 11230 3225
rect 8635 3170 8985 3175
rect 8605 3160 8985 3170
rect 8630 3145 8645 3160
rect 8775 3145 8790 3160
rect 6665 3030 6680 3045
rect 6720 3030 6735 3045
rect 6925 3005 6940 3045
rect 6980 3030 6995 3045
rect 7115 3005 7130 3045
rect 7170 3030 7185 3045
rect 7375 3030 7390 3045
rect 7430 3030 7445 3045
rect 7635 3030 7650 3045
rect 7690 3030 7705 3045
rect 7855 3030 7870 3045
rect 8020 3030 8035 3045
rect 8240 3030 8255 3045
rect 8435 3030 8450 3045
rect 8630 3030 8645 3045
rect 8775 3030 8790 3045
rect 6925 2990 7130 3005
rect 7690 3020 7730 3030
rect 7690 3000 7700 3020
rect 7720 3000 7730 3020
rect 7690 2990 7730 3000
<< polycont >>
rect 8460 4070 8480 4090
rect 8775 4070 8795 4090
rect 9680 4045 9700 4065
rect 11200 4045 11220 4065
rect 6575 3880 6595 3900
rect 6740 3900 6760 3920
rect 7000 3860 7020 3880
rect 7190 3900 7210 3920
rect 6800 3650 6820 3670
rect 7535 3875 7555 3895
rect 7575 3875 7595 3895
rect 7740 3875 7760 3895
rect 7905 3875 7925 3895
rect 8050 3875 8070 3895
rect 8125 3880 8145 3900
rect 8485 3865 8505 3885
rect 8680 3905 8700 3925
rect 7250 3650 7270 3670
rect 9900 3780 9920 3800
rect 10170 3775 10190 3795
rect 10710 3775 10730 3795
rect 10915 3760 10935 3780
rect 11045 3760 11065 3780
rect 6860 3590 6880 3610
rect 8420 3590 8440 3610
rect 7635 3480 7655 3500
rect 10110 3495 10130 3515
rect 10490 3495 10510 3515
rect 10695 3510 10715 3530
rect 11045 3510 11065 3530
rect 6800 3420 6820 3440
rect 6575 3190 6595 3210
rect 6740 3170 6760 3190
rect 7250 3420 7270 3440
rect 7000 3210 7020 3230
rect 7190 3170 7210 3190
rect 7525 3175 7545 3195
rect 7740 3195 7760 3215
rect 7905 3195 7925 3215
rect 8070 3195 8090 3215
rect 8135 3180 8155 3200
rect 8420 3195 8440 3215
rect 8680 3210 8700 3230
rect 8855 3210 8875 3230
rect 8615 3170 8635 3190
rect 9780 3225 9800 3245
rect 11200 3225 11220 3245
rect 7700 3000 7720 3020
<< locali >>
rect 11545 4190 11600 4200
rect 11545 4155 11555 4190
rect 11590 4155 11600 4190
rect 6625 4145 6665 4155
rect 6625 4125 6635 4145
rect 6655 4125 6665 4145
rect 6625 4115 6665 4125
rect 6735 4145 6775 4155
rect 6735 4125 6745 4145
rect 6765 4125 6775 4145
rect 6735 4115 6775 4125
rect 6885 4145 6925 4155
rect 6885 4125 6895 4145
rect 6915 4125 6925 4145
rect 6885 4115 6925 4125
rect 7000 4145 7040 4155
rect 7000 4125 7010 4145
rect 7030 4125 7040 4145
rect 7000 4115 7040 4125
rect 7075 4145 7115 4155
rect 7075 4125 7085 4145
rect 7105 4125 7115 4145
rect 7075 4115 7115 4125
rect 7185 4145 7225 4155
rect 7185 4125 7195 4145
rect 7215 4125 7225 4145
rect 7185 4115 7225 4125
rect 7335 4145 7375 4155
rect 7335 4125 7345 4145
rect 7365 4125 7375 4145
rect 7335 4115 7375 4125
rect 7445 4145 7485 4155
rect 7445 4125 7455 4145
rect 7475 4125 7485 4145
rect 7445 4115 7485 4125
rect 7645 4145 7685 4155
rect 7645 4125 7655 4145
rect 7675 4125 7685 4145
rect 7645 4115 7685 4125
rect 7810 4145 7850 4155
rect 7810 4125 7820 4145
rect 7840 4125 7850 4145
rect 7810 4115 7850 4125
rect 7975 4145 8015 4155
rect 7975 4125 7985 4145
rect 8005 4125 8015 4145
rect 7975 4115 8015 4125
rect 8195 4145 8235 4155
rect 8195 4125 8205 4145
rect 8225 4125 8235 4145
rect 8195 4115 8235 4125
rect 8585 4145 8625 4155
rect 8585 4125 8595 4145
rect 8615 4125 8625 4145
rect 8585 4115 8625 4125
rect 8925 4145 8965 4155
rect 11545 4145 11600 4155
rect 8925 4125 8935 4145
rect 8955 4125 8965 4145
rect 8925 4115 8965 4125
rect 6635 4040 6655 4115
rect 6745 4040 6765 4115
rect 6895 4040 6915 4115
rect 7010 4040 7030 4115
rect 7085 4040 7105 4115
rect 7195 4040 7215 4115
rect 7345 4040 7365 4115
rect 7455 4040 7475 4115
rect 7655 4040 7675 4115
rect 7820 4040 7840 4115
rect 7985 4040 8005 4115
rect 8205 4040 8225 4115
rect 8450 4090 8490 4100
rect 8450 4070 8460 4090
rect 8480 4070 8490 4090
rect 8450 4060 8490 4070
rect 8595 4040 8615 4115
rect 8765 4090 8805 4100
rect 8765 4070 8775 4090
rect 8795 4070 8805 4090
rect 8765 4060 8805 4070
rect 8935 4040 8955 4115
rect 9670 4065 9710 4075
rect 9670 4045 9680 4065
rect 9700 4045 9710 4065
rect 6590 4030 6660 4040
rect 6590 4010 6595 4030
rect 6615 4010 6635 4030
rect 6655 4010 6660 4030
rect 6590 3980 6660 4010
rect 6590 3960 6595 3980
rect 6615 3960 6635 3980
rect 6655 3960 6660 3980
rect 6590 3950 6660 3960
rect 6685 4030 6715 4040
rect 6685 4010 6690 4030
rect 6710 4010 6715 4030
rect 6685 3980 6715 4010
rect 6685 3960 6690 3980
rect 6710 3960 6715 3980
rect 6685 3950 6715 3960
rect 6740 4030 6770 4040
rect 6740 4010 6745 4030
rect 6765 4010 6770 4030
rect 6740 3980 6770 4010
rect 6740 3960 6745 3980
rect 6765 3960 6770 3980
rect 6740 3950 6770 3960
rect 6890 4030 6920 4040
rect 6890 4010 6895 4030
rect 6915 4010 6920 4030
rect 6890 3980 6920 4010
rect 6890 3960 6895 3980
rect 6915 3960 6920 3980
rect 6890 3950 6920 3960
rect 6945 4030 6975 4040
rect 6945 4010 6950 4030
rect 6970 4010 6975 4030
rect 6945 3980 6975 4010
rect 6945 3960 6950 3980
rect 6970 3960 6975 3980
rect 6945 3950 6975 3960
rect 7000 4030 7110 4040
rect 7000 4010 7005 4030
rect 7025 4010 7045 4030
rect 7065 4010 7085 4030
rect 7105 4010 7110 4030
rect 7000 3980 7110 4010
rect 7000 3960 7005 3980
rect 7025 3960 7045 3980
rect 7065 3960 7085 3980
rect 7105 3960 7110 3980
rect 7000 3950 7110 3960
rect 7135 4030 7165 4040
rect 7135 4010 7140 4030
rect 7160 4010 7165 4030
rect 7135 3980 7165 4010
rect 7135 3960 7140 3980
rect 7160 3960 7165 3980
rect 7135 3950 7165 3960
rect 7190 4030 7220 4040
rect 7190 4010 7195 4030
rect 7215 4010 7220 4030
rect 7190 3980 7220 4010
rect 7190 3960 7195 3980
rect 7215 3960 7220 3980
rect 7190 3950 7220 3960
rect 7340 4030 7370 4040
rect 7340 4010 7345 4030
rect 7365 4010 7370 4030
rect 7340 3980 7370 4010
rect 7340 3960 7345 3980
rect 7365 3960 7370 3980
rect 7340 3950 7370 3960
rect 7395 4030 7425 4040
rect 7395 4010 7400 4030
rect 7420 4010 7425 4030
rect 7395 3980 7425 4010
rect 7395 3960 7400 3980
rect 7420 3960 7425 3980
rect 7395 3950 7425 3960
rect 7450 4030 7520 4040
rect 7450 4010 7455 4030
rect 7475 4010 7495 4030
rect 7515 4010 7520 4030
rect 7450 3980 7520 4010
rect 7450 3960 7455 3980
rect 7475 3960 7495 3980
rect 7515 3960 7520 3980
rect 7450 3950 7520 3960
rect 7595 4030 7625 4040
rect 7595 4010 7600 4030
rect 7620 4010 7625 4030
rect 7595 3980 7625 4010
rect 7595 3960 7600 3980
rect 7620 3960 7625 3980
rect 7595 3950 7625 3960
rect 7650 4030 7720 4040
rect 7650 4010 7655 4030
rect 7675 4010 7695 4030
rect 7715 4010 7720 4030
rect 7650 3980 7720 4010
rect 7650 3960 7655 3980
rect 7675 3960 7695 3980
rect 7715 3960 7720 3980
rect 7650 3950 7720 3960
rect 7760 4030 7790 4040
rect 7760 4010 7765 4030
rect 7785 4010 7790 4030
rect 7760 3980 7790 4010
rect 7760 3960 7765 3980
rect 7785 3960 7790 3980
rect 7760 3950 7790 3960
rect 7815 4030 7885 4040
rect 7815 4010 7820 4030
rect 7840 4010 7860 4030
rect 7880 4010 7885 4030
rect 7815 3980 7885 4010
rect 7815 3960 7820 3980
rect 7840 3960 7860 3980
rect 7880 3960 7885 3980
rect 7815 3950 7885 3960
rect 7925 4030 7955 4040
rect 7925 4010 7930 4030
rect 7950 4010 7955 4030
rect 7925 3980 7955 4010
rect 7925 3960 7930 3980
rect 7950 3960 7955 3980
rect 7925 3950 7955 3960
rect 7980 4030 8050 4040
rect 7980 4010 7985 4030
rect 8005 4010 8025 4030
rect 8045 4010 8050 4030
rect 7980 3980 8050 4010
rect 7980 3960 7985 3980
rect 8005 3960 8025 3980
rect 8045 3960 8050 3980
rect 7980 3950 8050 3960
rect 8145 4030 8235 4040
rect 8145 4010 8155 4030
rect 8175 4010 8205 4030
rect 8225 4010 8235 4030
rect 8145 3980 8235 4010
rect 8145 3960 8155 3980
rect 8175 3960 8205 3980
rect 8225 3960 8235 3980
rect 8145 3950 8235 3960
rect 8260 4030 8300 4040
rect 8260 4010 8270 4030
rect 8290 4010 8300 4030
rect 8260 3980 8300 4010
rect 8260 3960 8270 3980
rect 8290 3960 8300 3980
rect 8260 3950 8300 3960
rect 8390 4030 8430 4040
rect 8390 4010 8400 4030
rect 8420 4010 8430 4030
rect 8390 3980 8430 4010
rect 8390 3960 8400 3980
rect 8420 3960 8430 3980
rect 8390 3950 8430 3960
rect 8455 4030 8495 4040
rect 8455 4010 8465 4030
rect 8485 4010 8495 4030
rect 8455 3980 8495 4010
rect 8455 3960 8465 3980
rect 8485 3960 8495 3980
rect 8455 3950 8495 3960
rect 8535 4030 8625 4040
rect 8535 4010 8545 4030
rect 8565 4010 8595 4030
rect 8615 4010 8625 4030
rect 8535 3980 8625 4010
rect 8535 3960 8545 3980
rect 8565 3960 8595 3980
rect 8615 3960 8625 3980
rect 8535 3950 8625 3960
rect 8650 4030 8690 4040
rect 8650 4010 8660 4030
rect 8680 4010 8690 4030
rect 8650 3980 8690 4010
rect 8650 3960 8660 3980
rect 8680 3960 8690 3980
rect 8650 3950 8690 3960
rect 8730 4030 8770 4040
rect 8730 4010 8740 4030
rect 8760 4010 8770 4030
rect 8730 3980 8770 4010
rect 8730 3960 8740 3980
rect 8760 3960 8770 3980
rect 8730 3950 8770 3960
rect 8795 4030 8835 4040
rect 8795 4010 8805 4030
rect 8825 4010 8835 4030
rect 8795 3980 8835 4010
rect 8795 3960 8805 3980
rect 8825 3960 8835 3980
rect 8795 3950 8835 3960
rect 8875 4030 8965 4040
rect 8875 4010 8885 4030
rect 8905 4010 8935 4030
rect 8955 4010 8965 4030
rect 8875 3980 8965 4010
rect 8875 3960 8885 3980
rect 8905 3960 8935 3980
rect 8955 3960 8965 3980
rect 8875 3950 8965 3960
rect 8990 4030 9030 4040
rect 9670 4035 9710 4045
rect 11190 4065 11230 4075
rect 11190 4045 11200 4065
rect 11220 4045 11230 4065
rect 11190 4035 11230 4045
rect 8990 4010 9000 4030
rect 9020 4010 9030 4030
rect 8990 3980 9030 4010
rect 8990 3960 9000 3980
rect 9020 3960 9030 3980
rect 8990 3950 9030 3960
rect 9620 4005 9710 4015
rect 9620 3985 9630 4005
rect 9650 3985 9680 4005
rect 9700 3985 9710 4005
rect 9620 3955 9710 3985
rect 6565 3900 6605 3910
rect 6565 3880 6575 3900
rect 6595 3880 6605 3900
rect 6565 3870 6605 3880
rect 6685 3870 6705 3950
rect 6730 3920 6770 3930
rect 6730 3900 6740 3920
rect 6760 3910 6770 3920
rect 6760 3900 6870 3910
rect 6730 3890 6870 3900
rect 6685 3850 6765 3870
rect 6745 3830 6765 3850
rect 6590 3820 6660 3830
rect 6590 3800 6595 3820
rect 6615 3800 6635 3820
rect 6655 3800 6660 3820
rect 6590 3770 6660 3800
rect 6590 3750 6595 3770
rect 6615 3750 6635 3770
rect 6655 3750 6660 3770
rect 6590 3720 6660 3750
rect 6590 3700 6595 3720
rect 6615 3700 6635 3720
rect 6655 3700 6660 3720
rect 6590 3670 6660 3700
rect 6590 3650 6595 3670
rect 6615 3650 6635 3670
rect 6655 3650 6660 3670
rect 6590 3640 6660 3650
rect 6685 3820 6715 3830
rect 6685 3800 6690 3820
rect 6710 3800 6715 3820
rect 6685 3770 6715 3800
rect 6685 3750 6690 3770
rect 6710 3750 6715 3770
rect 6685 3720 6715 3750
rect 6685 3700 6690 3720
rect 6710 3700 6715 3720
rect 6685 3670 6715 3700
rect 6685 3650 6690 3670
rect 6710 3650 6715 3670
rect 6685 3640 6715 3650
rect 6740 3820 6770 3830
rect 6740 3800 6745 3820
rect 6765 3800 6770 3820
rect 6740 3770 6770 3800
rect 6740 3750 6745 3770
rect 6765 3750 6770 3770
rect 6740 3720 6770 3750
rect 6740 3700 6745 3720
rect 6765 3700 6770 3720
rect 6740 3670 6770 3700
rect 6740 3650 6745 3670
rect 6765 3665 6770 3670
rect 6790 3670 6830 3680
rect 6790 3665 6800 3670
rect 6765 3650 6800 3665
rect 6820 3650 6830 3670
rect 6740 3640 6830 3650
rect 6850 3660 6870 3890
rect 6950 3870 6970 3950
rect 6895 3850 6970 3870
rect 6990 3880 7030 3890
rect 6990 3860 7000 3880
rect 7020 3870 7030 3880
rect 7135 3870 7155 3950
rect 7180 3920 7220 3930
rect 7180 3900 7190 3920
rect 7210 3910 7220 3920
rect 7210 3900 7320 3910
rect 7180 3890 7320 3900
rect 7020 3860 7215 3870
rect 6990 3850 7215 3860
rect 6895 3830 6915 3850
rect 7195 3830 7215 3850
rect 6890 3820 6920 3830
rect 6890 3800 6895 3820
rect 6915 3800 6920 3820
rect 6890 3770 6920 3800
rect 6890 3750 6895 3770
rect 6915 3750 6920 3770
rect 6890 3720 6920 3750
rect 6890 3700 6895 3720
rect 6915 3700 6920 3720
rect 6890 3670 6920 3700
rect 6890 3660 6895 3670
rect 6850 3650 6895 3660
rect 6915 3650 6920 3670
rect 6850 3640 6920 3650
rect 6945 3820 6975 3830
rect 6945 3800 6950 3820
rect 6970 3800 6975 3820
rect 6945 3770 6975 3800
rect 6945 3750 6950 3770
rect 6970 3750 6975 3770
rect 6945 3720 6975 3750
rect 6945 3700 6950 3720
rect 6970 3700 6975 3720
rect 6945 3670 6975 3700
rect 6945 3650 6950 3670
rect 6970 3650 6975 3670
rect 6945 3640 6975 3650
rect 7000 3820 7110 3830
rect 7000 3800 7005 3820
rect 7025 3800 7045 3820
rect 7065 3800 7085 3820
rect 7105 3800 7110 3820
rect 7000 3770 7110 3800
rect 7000 3750 7005 3770
rect 7025 3750 7045 3770
rect 7065 3750 7085 3770
rect 7105 3750 7110 3770
rect 7000 3720 7110 3750
rect 7000 3700 7005 3720
rect 7025 3700 7045 3720
rect 7065 3700 7085 3720
rect 7105 3700 7110 3720
rect 7000 3670 7110 3700
rect 7000 3650 7005 3670
rect 7025 3650 7045 3670
rect 7065 3650 7085 3670
rect 7105 3650 7110 3670
rect 7000 3640 7110 3650
rect 7135 3820 7165 3830
rect 7135 3800 7140 3820
rect 7160 3800 7165 3820
rect 7135 3770 7165 3800
rect 7135 3750 7140 3770
rect 7160 3750 7165 3770
rect 7135 3720 7165 3750
rect 7135 3700 7140 3720
rect 7160 3700 7165 3720
rect 7135 3670 7165 3700
rect 7135 3650 7140 3670
rect 7160 3650 7165 3670
rect 7135 3640 7165 3650
rect 7190 3820 7220 3830
rect 7190 3800 7195 3820
rect 7215 3800 7220 3820
rect 7190 3770 7220 3800
rect 7190 3750 7195 3770
rect 7215 3750 7220 3770
rect 7190 3720 7220 3750
rect 7190 3700 7195 3720
rect 7215 3700 7220 3720
rect 7190 3670 7220 3700
rect 7190 3650 7195 3670
rect 7215 3665 7220 3670
rect 7240 3670 7280 3680
rect 7240 3665 7250 3670
rect 7215 3650 7250 3665
rect 7270 3650 7280 3670
rect 7190 3640 7280 3650
rect 7300 3660 7320 3890
rect 7400 3870 7420 3950
rect 7595 3905 7615 3950
rect 7760 3905 7780 3950
rect 7925 3905 7945 3950
rect 7345 3850 7420 3870
rect 7525 3895 7615 3905
rect 7525 3875 7535 3895
rect 7555 3875 7575 3895
rect 7595 3875 7615 3895
rect 7525 3865 7615 3875
rect 7730 3895 7780 3905
rect 7730 3875 7740 3895
rect 7760 3875 7780 3895
rect 7730 3865 7780 3875
rect 7895 3895 7945 3905
rect 7895 3875 7905 3895
rect 7925 3875 7945 3895
rect 7895 3865 7945 3875
rect 8040 3895 8080 3905
rect 8040 3875 8050 3895
rect 8070 3875 8080 3895
rect 8040 3865 8080 3875
rect 8115 3900 8155 3910
rect 8115 3880 8125 3900
rect 8145 3880 8155 3900
rect 8115 3870 8155 3880
rect 8270 3870 8290 3950
rect 8400 3870 8420 3950
rect 7345 3830 7365 3850
rect 7595 3830 7615 3865
rect 7760 3830 7780 3865
rect 7925 3830 7945 3865
rect 8270 3850 8420 3870
rect 8270 3830 8290 3850
rect 8400 3830 8420 3850
rect 8465 3895 8485 3950
rect 8670 3935 8690 3950
rect 8670 3925 8710 3935
rect 8670 3905 8680 3925
rect 8700 3905 8710 3925
rect 8670 3900 8710 3905
rect 8465 3885 8515 3895
rect 8465 3865 8485 3885
rect 8505 3865 8515 3885
rect 8465 3855 8515 3865
rect 8465 3830 8485 3855
rect 8670 3830 8690 3900
rect 8740 3830 8760 3950
rect 8805 3910 8825 3950
rect 9000 3930 9020 3950
rect 9620 3935 9630 3955
rect 9650 3935 9680 3955
rect 9700 3935 9710 3955
rect 9000 3920 9040 3930
rect 9000 3910 9010 3920
rect 8805 3900 9010 3910
rect 9030 3900 9040 3920
rect 8805 3890 9040 3900
rect 9620 3905 9710 3935
rect 8805 3830 8825 3890
rect 9620 3885 9630 3905
rect 9650 3885 9680 3905
rect 9700 3885 9710 3905
rect 9620 3855 9710 3885
rect 9620 3835 9630 3855
rect 9650 3835 9680 3855
rect 9700 3835 9710 3855
rect 7340 3820 7370 3830
rect 7340 3800 7345 3820
rect 7365 3800 7370 3820
rect 7340 3770 7370 3800
rect 7340 3750 7345 3770
rect 7365 3750 7370 3770
rect 7340 3720 7370 3750
rect 7340 3700 7345 3720
rect 7365 3700 7370 3720
rect 7340 3670 7370 3700
rect 7340 3660 7345 3670
rect 7300 3650 7345 3660
rect 7365 3650 7370 3670
rect 7300 3640 7370 3650
rect 7395 3820 7425 3830
rect 7395 3800 7400 3820
rect 7420 3800 7425 3820
rect 7395 3770 7425 3800
rect 7395 3750 7400 3770
rect 7420 3750 7425 3770
rect 7395 3720 7425 3750
rect 7395 3700 7400 3720
rect 7420 3700 7425 3720
rect 7395 3670 7425 3700
rect 7395 3650 7400 3670
rect 7420 3650 7425 3670
rect 7395 3640 7425 3650
rect 7450 3820 7520 3830
rect 7450 3800 7455 3820
rect 7475 3800 7495 3820
rect 7515 3800 7520 3820
rect 7450 3770 7520 3800
rect 7450 3750 7455 3770
rect 7475 3750 7495 3770
rect 7515 3750 7520 3770
rect 7450 3720 7520 3750
rect 7450 3700 7455 3720
rect 7475 3700 7495 3720
rect 7515 3700 7520 3720
rect 7450 3670 7520 3700
rect 7450 3650 7455 3670
rect 7475 3650 7495 3670
rect 7515 3650 7520 3670
rect 7450 3640 7520 3650
rect 7595 3820 7625 3830
rect 7595 3800 7600 3820
rect 7620 3800 7625 3820
rect 7595 3770 7625 3800
rect 7595 3750 7600 3770
rect 7620 3750 7625 3770
rect 7595 3720 7625 3750
rect 7595 3700 7600 3720
rect 7620 3700 7625 3720
rect 7595 3670 7625 3700
rect 7595 3650 7600 3670
rect 7620 3650 7625 3670
rect 7595 3640 7625 3650
rect 7650 3820 7720 3830
rect 7650 3800 7655 3820
rect 7675 3800 7695 3820
rect 7715 3800 7720 3820
rect 7650 3770 7720 3800
rect 7650 3750 7655 3770
rect 7675 3750 7695 3770
rect 7715 3750 7720 3770
rect 7650 3720 7720 3750
rect 7650 3700 7655 3720
rect 7675 3700 7695 3720
rect 7715 3700 7720 3720
rect 7650 3670 7720 3700
rect 7650 3650 7655 3670
rect 7675 3650 7695 3670
rect 7715 3650 7720 3670
rect 7650 3640 7720 3650
rect 7760 3820 7790 3830
rect 7760 3800 7765 3820
rect 7785 3800 7790 3820
rect 7760 3770 7790 3800
rect 7760 3750 7765 3770
rect 7785 3750 7790 3770
rect 7760 3720 7790 3750
rect 7760 3700 7765 3720
rect 7785 3700 7790 3720
rect 7760 3670 7790 3700
rect 7760 3650 7765 3670
rect 7785 3650 7790 3670
rect 7760 3640 7790 3650
rect 7815 3820 7885 3830
rect 7815 3800 7820 3820
rect 7840 3800 7860 3820
rect 7880 3800 7885 3820
rect 7815 3770 7885 3800
rect 7815 3750 7820 3770
rect 7840 3750 7860 3770
rect 7880 3750 7885 3770
rect 7815 3720 7885 3750
rect 7815 3700 7820 3720
rect 7840 3700 7860 3720
rect 7880 3700 7885 3720
rect 7815 3670 7885 3700
rect 7815 3650 7820 3670
rect 7840 3650 7860 3670
rect 7880 3650 7885 3670
rect 7815 3640 7885 3650
rect 7925 3820 7955 3830
rect 7925 3800 7930 3820
rect 7950 3800 7955 3820
rect 7925 3770 7955 3800
rect 7925 3750 7930 3770
rect 7950 3750 7955 3770
rect 7925 3720 7955 3750
rect 7925 3700 7930 3720
rect 7950 3700 7955 3720
rect 7925 3670 7955 3700
rect 7925 3650 7930 3670
rect 7950 3650 7955 3670
rect 7925 3640 7955 3650
rect 7980 3820 8050 3830
rect 7980 3800 7985 3820
rect 8005 3800 8025 3820
rect 8045 3800 8050 3820
rect 7980 3770 8050 3800
rect 7980 3750 7985 3770
rect 8005 3750 8025 3770
rect 8045 3750 8050 3770
rect 7980 3720 8050 3750
rect 7980 3700 7985 3720
rect 8005 3700 8025 3720
rect 8045 3700 8050 3720
rect 7980 3670 8050 3700
rect 7980 3650 7985 3670
rect 8005 3650 8025 3670
rect 8045 3650 8050 3670
rect 7980 3640 8050 3650
rect 8145 3820 8235 3830
rect 8145 3800 8155 3820
rect 8175 3800 8205 3820
rect 8225 3800 8235 3820
rect 8145 3770 8235 3800
rect 8145 3750 8155 3770
rect 8175 3750 8205 3770
rect 8225 3750 8235 3770
rect 8145 3720 8235 3750
rect 8145 3700 8155 3720
rect 8175 3700 8205 3720
rect 8225 3700 8235 3720
rect 8145 3670 8235 3700
rect 8145 3650 8155 3670
rect 8175 3650 8205 3670
rect 8225 3650 8235 3670
rect 8145 3640 8235 3650
rect 8260 3820 8300 3830
rect 8260 3800 8270 3820
rect 8290 3800 8300 3820
rect 8260 3770 8300 3800
rect 8260 3750 8270 3770
rect 8290 3750 8300 3770
rect 8260 3720 8300 3750
rect 8260 3700 8270 3720
rect 8290 3700 8300 3720
rect 8260 3670 8300 3700
rect 8260 3650 8270 3670
rect 8290 3650 8300 3670
rect 8260 3640 8300 3650
rect 8390 3820 8430 3830
rect 8390 3800 8400 3820
rect 8420 3800 8430 3820
rect 8390 3770 8430 3800
rect 8390 3750 8400 3770
rect 8420 3750 8430 3770
rect 8390 3720 8430 3750
rect 8390 3700 8400 3720
rect 8420 3700 8430 3720
rect 8390 3670 8430 3700
rect 8390 3650 8400 3670
rect 8420 3650 8430 3670
rect 8390 3640 8430 3650
rect 8455 3820 8495 3830
rect 8455 3800 8465 3820
rect 8485 3800 8495 3820
rect 8455 3770 8495 3800
rect 8455 3750 8465 3770
rect 8485 3750 8495 3770
rect 8455 3720 8495 3750
rect 8455 3700 8465 3720
rect 8485 3700 8495 3720
rect 8455 3670 8495 3700
rect 8455 3650 8465 3670
rect 8485 3650 8495 3670
rect 8455 3640 8495 3650
rect 8535 3820 8625 3830
rect 8535 3800 8545 3820
rect 8565 3800 8595 3820
rect 8615 3800 8625 3820
rect 8535 3770 8625 3800
rect 8535 3750 8545 3770
rect 8565 3750 8595 3770
rect 8615 3750 8625 3770
rect 8535 3720 8625 3750
rect 8535 3700 8545 3720
rect 8565 3700 8595 3720
rect 8615 3700 8625 3720
rect 8535 3670 8625 3700
rect 8535 3650 8545 3670
rect 8565 3650 8595 3670
rect 8615 3650 8625 3670
rect 8535 3640 8625 3650
rect 8650 3820 8690 3830
rect 8650 3800 8660 3820
rect 8680 3800 8690 3820
rect 8650 3770 8690 3800
rect 8650 3750 8660 3770
rect 8680 3750 8690 3770
rect 8650 3720 8690 3750
rect 8650 3700 8660 3720
rect 8680 3700 8690 3720
rect 8650 3670 8690 3700
rect 8650 3650 8660 3670
rect 8680 3650 8690 3670
rect 8650 3640 8690 3650
rect 8730 3820 8770 3830
rect 8730 3800 8740 3820
rect 8760 3800 8770 3820
rect 8730 3770 8770 3800
rect 8730 3750 8740 3770
rect 8760 3750 8770 3770
rect 8730 3720 8770 3750
rect 8730 3700 8740 3720
rect 8760 3700 8770 3720
rect 8730 3670 8770 3700
rect 8730 3650 8740 3670
rect 8760 3650 8770 3670
rect 8730 3640 8770 3650
rect 8795 3820 8835 3830
rect 9620 3825 9710 3835
rect 9780 4005 9820 4015
rect 9780 3985 9790 4005
rect 9810 3985 9820 4005
rect 9780 3955 9820 3985
rect 9780 3935 9790 3955
rect 9810 3935 9820 3955
rect 9780 3905 9820 3935
rect 9780 3885 9790 3905
rect 9810 3885 9820 3905
rect 9780 3855 9820 3885
rect 9780 3835 9790 3855
rect 9810 3835 9820 3855
rect 9780 3825 9820 3835
rect 9890 4005 9930 4015
rect 9890 3985 9900 4005
rect 9920 3985 9930 4005
rect 9890 3955 9930 3985
rect 9890 3935 9900 3955
rect 9920 3935 9930 3955
rect 9890 3905 9930 3935
rect 9890 3885 9900 3905
rect 9920 3885 9930 3905
rect 9890 3855 9930 3885
rect 9890 3835 9900 3855
rect 9920 3835 9930 3855
rect 8795 3800 8805 3820
rect 8825 3800 8835 3820
rect 8795 3770 8835 3800
rect 9890 3800 9930 3835
rect 10000 4005 10040 4015
rect 10000 3985 10010 4005
rect 10030 3985 10040 4005
rect 10000 3955 10040 3985
rect 10000 3935 10010 3955
rect 10030 3935 10040 3955
rect 10000 3905 10040 3935
rect 10000 3885 10010 3905
rect 10030 3885 10040 3905
rect 10000 3855 10040 3885
rect 10000 3835 10010 3855
rect 10030 3835 10040 3855
rect 10000 3825 10040 3835
rect 10110 4005 10250 4015
rect 10110 3985 10120 4005
rect 10140 3985 10170 4005
rect 10190 3985 10220 4005
rect 10240 3985 10250 4005
rect 10110 3955 10250 3985
rect 10110 3935 10120 3955
rect 10140 3935 10170 3955
rect 10190 3935 10220 3955
rect 10240 3935 10250 3955
rect 10110 3905 10250 3935
rect 10110 3885 10120 3905
rect 10140 3885 10170 3905
rect 10190 3885 10220 3905
rect 10240 3885 10250 3905
rect 10110 3855 10250 3885
rect 10110 3835 10120 3855
rect 10140 3835 10170 3855
rect 10190 3835 10220 3855
rect 10240 3835 10250 3855
rect 10110 3825 10250 3835
rect 10320 4005 10360 4015
rect 10320 3985 10330 4005
rect 10350 3985 10360 4005
rect 10320 3955 10360 3985
rect 10320 3935 10330 3955
rect 10350 3935 10360 3955
rect 10320 3905 10360 3935
rect 10320 3885 10330 3905
rect 10350 3885 10360 3905
rect 10320 3855 10360 3885
rect 10320 3835 10330 3855
rect 10350 3835 10360 3855
rect 10320 3825 10360 3835
rect 10430 4005 10470 4015
rect 10430 3985 10440 4005
rect 10460 3985 10470 4005
rect 10430 3955 10470 3985
rect 10430 3935 10440 3955
rect 10460 3935 10470 3955
rect 10430 3905 10470 3935
rect 10430 3885 10440 3905
rect 10460 3885 10470 3905
rect 10430 3855 10470 3885
rect 10430 3835 10440 3855
rect 10460 3835 10470 3855
rect 10430 3825 10470 3835
rect 10540 4005 10580 4015
rect 10540 3985 10550 4005
rect 10570 3985 10580 4005
rect 10540 3955 10580 3985
rect 10540 3935 10550 3955
rect 10570 3935 10580 3955
rect 10540 3905 10580 3935
rect 10540 3885 10550 3905
rect 10570 3885 10580 3905
rect 10540 3855 10580 3885
rect 10540 3835 10550 3855
rect 10570 3835 10580 3855
rect 10540 3825 10580 3835
rect 10650 4005 10790 4015
rect 10650 3985 10660 4005
rect 10680 3985 10710 4005
rect 10730 3985 10760 4005
rect 10780 3985 10790 4005
rect 10650 3955 10790 3985
rect 10650 3935 10660 3955
rect 10680 3935 10710 3955
rect 10730 3935 10760 3955
rect 10780 3935 10790 3955
rect 10650 3905 10790 3935
rect 10650 3885 10660 3905
rect 10680 3885 10710 3905
rect 10730 3885 10760 3905
rect 10780 3885 10790 3905
rect 10650 3855 10790 3885
rect 10650 3835 10660 3855
rect 10680 3835 10710 3855
rect 10730 3835 10760 3855
rect 10780 3835 10790 3855
rect 10650 3825 10790 3835
rect 10860 4005 10900 4015
rect 10860 3985 10870 4005
rect 10890 3985 10900 4005
rect 10860 3955 10900 3985
rect 10860 3935 10870 3955
rect 10890 3935 10900 3955
rect 10860 3905 10900 3935
rect 10860 3885 10870 3905
rect 10890 3885 10900 3905
rect 10860 3855 10900 3885
rect 10860 3835 10870 3855
rect 10890 3835 10900 3855
rect 10860 3825 10900 3835
rect 10970 4005 11010 4015
rect 10970 3985 10980 4005
rect 11000 3985 11010 4005
rect 10970 3955 11010 3985
rect 10970 3935 10980 3955
rect 11000 3935 11010 3955
rect 10970 3905 11010 3935
rect 10970 3885 10980 3905
rect 11000 3885 11010 3905
rect 10970 3855 11010 3885
rect 10970 3835 10980 3855
rect 11000 3835 11010 3855
rect 10970 3825 11010 3835
rect 11080 4005 11120 4015
rect 11080 3985 11090 4005
rect 11110 3985 11120 4005
rect 11080 3955 11120 3985
rect 11080 3935 11090 3955
rect 11110 3935 11120 3955
rect 11080 3905 11120 3935
rect 11080 3885 11090 3905
rect 11110 3885 11120 3905
rect 11080 3855 11120 3885
rect 11080 3835 11090 3855
rect 11110 3835 11120 3855
rect 11080 3825 11120 3835
rect 11190 4005 11280 4015
rect 11190 3985 11200 4005
rect 11220 3985 11250 4005
rect 11270 3985 11280 4005
rect 11190 3955 11280 3985
rect 11190 3935 11200 3955
rect 11220 3935 11250 3955
rect 11270 3935 11280 3955
rect 11190 3905 11280 3935
rect 11190 3885 11200 3905
rect 11220 3885 11250 3905
rect 11270 3885 11280 3905
rect 11190 3855 11280 3885
rect 11190 3835 11200 3855
rect 11220 3835 11250 3855
rect 11270 3835 11280 3855
rect 11190 3825 11280 3835
rect 9890 3780 9900 3800
rect 9920 3780 9930 3800
rect 9890 3770 9930 3780
rect 10160 3795 10200 3825
rect 10160 3775 10170 3795
rect 10190 3775 10200 3795
rect 8795 3750 8805 3770
rect 8825 3750 8835 3770
rect 10160 3765 10200 3775
rect 10700 3795 10740 3825
rect 10700 3775 10710 3795
rect 10730 3775 10740 3795
rect 11370 3795 11425 3805
rect 10700 3765 10740 3775
rect 10905 3780 10945 3790
rect 10905 3760 10915 3780
rect 10935 3760 10945 3780
rect 10905 3750 10945 3760
rect 11035 3780 11075 3790
rect 11035 3760 11045 3780
rect 11065 3760 11075 3780
rect 11035 3750 11075 3760
rect 11370 3760 11380 3795
rect 11415 3760 11425 3795
rect 11370 3750 11425 3760
rect 8795 3720 8835 3750
rect 8795 3700 8805 3720
rect 8825 3700 8835 3720
rect 8795 3670 8835 3700
rect 8795 3650 8805 3670
rect 8825 3650 8835 3670
rect 8795 3640 8835 3650
rect 6635 3565 6655 3640
rect 6850 3620 6870 3640
rect 6850 3610 6890 3620
rect 6850 3590 6860 3610
rect 6880 3590 6890 3610
rect 6850 3580 6890 3590
rect 7005 3565 7025 3640
rect 7085 3565 7105 3640
rect 7455 3565 7475 3640
rect 7665 3565 7685 3640
rect 7820 3565 7840 3640
rect 7985 3565 8005 3640
rect 8205 3565 8225 3640
rect 8410 3610 8450 3620
rect 8410 3590 8420 3610
rect 8440 3590 8450 3610
rect 8410 3585 8450 3590
rect 8595 3565 8615 3640
rect 8740 3620 8760 3640
rect 8730 3610 8770 3620
rect 8730 3590 8740 3610
rect 8760 3590 8770 3610
rect 8730 3580 8770 3590
rect 6625 3555 6665 3565
rect 6625 3535 6635 3555
rect 6655 3535 6665 3555
rect 6625 3525 6665 3535
rect 6995 3555 7035 3565
rect 6995 3535 7005 3555
rect 7025 3535 7035 3555
rect 6995 3525 7035 3535
rect 7075 3555 7115 3565
rect 7075 3535 7085 3555
rect 7105 3535 7115 3555
rect 7075 3525 7115 3535
rect 7445 3555 7485 3565
rect 7445 3535 7455 3555
rect 7475 3535 7485 3555
rect 7445 3525 7485 3535
rect 7570 3555 7610 3565
rect 7570 3535 7580 3555
rect 7600 3535 7610 3555
rect 7570 3525 7610 3535
rect 7665 3555 7745 3565
rect 7665 3535 7675 3555
rect 7695 3535 7715 3555
rect 7735 3535 7745 3555
rect 7665 3525 7745 3535
rect 7810 3555 7850 3565
rect 7810 3535 7820 3555
rect 7840 3535 7850 3555
rect 7810 3525 7850 3535
rect 7975 3555 8015 3565
rect 7975 3535 7985 3555
rect 8005 3535 8015 3555
rect 7975 3525 8015 3535
rect 8195 3555 8235 3565
rect 8195 3535 8205 3555
rect 8225 3535 8235 3555
rect 8195 3525 8235 3535
rect 8390 3555 8430 3565
rect 8390 3535 8400 3555
rect 8420 3535 8430 3555
rect 8390 3525 8430 3535
rect 8585 3555 8625 3565
rect 8585 3535 8595 3555
rect 8615 3535 8625 3555
rect 8585 3525 8625 3535
rect 8925 3555 8965 3565
rect 8925 3535 8935 3555
rect 8955 3535 8965 3555
rect 8925 3525 8965 3535
rect 10685 3530 10725 3540
rect 6635 3450 6655 3525
rect 7005 3450 7025 3525
rect 7085 3450 7105 3525
rect 7455 3450 7475 3525
rect 7580 3450 7600 3525
rect 7625 3500 7665 3505
rect 7625 3480 7635 3500
rect 7655 3480 7665 3500
rect 7625 3470 7665 3480
rect 7715 3450 7735 3525
rect 7825 3450 7845 3525
rect 7990 3450 8010 3525
rect 8205 3450 8225 3525
rect 8400 3450 8420 3525
rect 8595 3450 8615 3525
rect 8935 3450 8955 3525
rect 10100 3515 10140 3525
rect 10100 3495 10110 3515
rect 10130 3495 10140 3515
rect 10100 3485 10140 3495
rect 10480 3515 10520 3525
rect 10480 3495 10490 3515
rect 10510 3495 10520 3515
rect 10685 3510 10695 3530
rect 10715 3510 10725 3530
rect 10685 3500 10725 3510
rect 11035 3530 11075 3540
rect 11035 3510 11045 3530
rect 11065 3510 11075 3530
rect 11035 3500 11075 3510
rect 11370 3530 11425 3540
rect 10480 3465 10520 3495
rect 11370 3495 11380 3530
rect 11415 3495 11425 3530
rect 11370 3485 11425 3495
rect 9720 3455 9810 3465
rect 6590 3440 6660 3450
rect 6590 3420 6595 3440
rect 6615 3420 6635 3440
rect 6655 3420 6660 3440
rect 6590 3390 6660 3420
rect 6590 3370 6595 3390
rect 6615 3370 6635 3390
rect 6655 3370 6660 3390
rect 6590 3340 6660 3370
rect 6590 3320 6595 3340
rect 6615 3320 6635 3340
rect 6655 3320 6660 3340
rect 6590 3290 6660 3320
rect 6590 3270 6595 3290
rect 6615 3270 6635 3290
rect 6655 3270 6660 3290
rect 6590 3260 6660 3270
rect 6685 3440 6715 3450
rect 6685 3420 6690 3440
rect 6710 3420 6715 3440
rect 6685 3390 6715 3420
rect 6685 3370 6690 3390
rect 6710 3370 6715 3390
rect 6685 3340 6715 3370
rect 6685 3320 6690 3340
rect 6710 3320 6715 3340
rect 6685 3290 6715 3320
rect 6685 3270 6690 3290
rect 6710 3270 6715 3290
rect 6685 3260 6715 3270
rect 6740 3440 6830 3450
rect 6740 3420 6745 3440
rect 6765 3425 6800 3440
rect 6765 3420 6770 3425
rect 6740 3390 6770 3420
rect 6790 3420 6800 3425
rect 6820 3420 6830 3440
rect 6790 3410 6830 3420
rect 6850 3440 6920 3450
rect 6850 3430 6895 3440
rect 6740 3370 6745 3390
rect 6765 3370 6770 3390
rect 6740 3340 6770 3370
rect 6740 3320 6745 3340
rect 6765 3320 6770 3340
rect 6740 3290 6770 3320
rect 6740 3270 6745 3290
rect 6765 3270 6770 3290
rect 6740 3260 6770 3270
rect 6745 3240 6765 3260
rect 6685 3220 6765 3240
rect 6565 3210 6605 3220
rect 6565 3190 6575 3210
rect 6595 3190 6605 3210
rect 6565 3180 6605 3190
rect 6685 3140 6705 3220
rect 6850 3200 6870 3430
rect 6890 3420 6895 3430
rect 6915 3420 6920 3440
rect 6890 3390 6920 3420
rect 6890 3370 6895 3390
rect 6915 3370 6920 3390
rect 6890 3340 6920 3370
rect 6890 3320 6895 3340
rect 6915 3320 6920 3340
rect 6890 3290 6920 3320
rect 6890 3270 6895 3290
rect 6915 3270 6920 3290
rect 6890 3260 6920 3270
rect 6945 3440 6975 3450
rect 6945 3420 6950 3440
rect 6970 3420 6975 3440
rect 6945 3390 6975 3420
rect 6945 3370 6950 3390
rect 6970 3370 6975 3390
rect 6945 3340 6975 3370
rect 6945 3320 6950 3340
rect 6970 3320 6975 3340
rect 6945 3290 6975 3320
rect 6945 3270 6950 3290
rect 6970 3270 6975 3290
rect 6945 3260 6975 3270
rect 7000 3440 7110 3450
rect 7000 3420 7005 3440
rect 7025 3420 7045 3440
rect 7065 3420 7085 3440
rect 7105 3420 7110 3440
rect 7000 3390 7110 3420
rect 7000 3370 7005 3390
rect 7025 3370 7045 3390
rect 7065 3370 7085 3390
rect 7105 3370 7110 3390
rect 7000 3340 7110 3370
rect 7000 3320 7005 3340
rect 7025 3320 7045 3340
rect 7065 3320 7085 3340
rect 7105 3320 7110 3340
rect 7000 3290 7110 3320
rect 7000 3270 7005 3290
rect 7025 3270 7045 3290
rect 7065 3270 7085 3290
rect 7105 3270 7110 3290
rect 7000 3260 7110 3270
rect 7135 3440 7165 3450
rect 7135 3420 7140 3440
rect 7160 3420 7165 3440
rect 7135 3390 7165 3420
rect 7135 3370 7140 3390
rect 7160 3370 7165 3390
rect 7135 3340 7165 3370
rect 7135 3320 7140 3340
rect 7160 3320 7165 3340
rect 7135 3290 7165 3320
rect 7135 3270 7140 3290
rect 7160 3270 7165 3290
rect 7135 3260 7165 3270
rect 7190 3440 7280 3450
rect 7190 3420 7195 3440
rect 7215 3425 7250 3440
rect 7215 3420 7220 3425
rect 7190 3390 7220 3420
rect 7240 3420 7250 3425
rect 7270 3420 7280 3440
rect 7240 3410 7280 3420
rect 7300 3440 7370 3450
rect 7300 3430 7345 3440
rect 7190 3370 7195 3390
rect 7215 3370 7220 3390
rect 7190 3340 7220 3370
rect 7190 3320 7195 3340
rect 7215 3320 7220 3340
rect 7190 3290 7220 3320
rect 7190 3270 7195 3290
rect 7215 3270 7220 3290
rect 7190 3260 7220 3270
rect 6895 3240 6915 3260
rect 7195 3240 7215 3260
rect 6895 3220 6970 3240
rect 6730 3190 6870 3200
rect 6730 3170 6740 3190
rect 6760 3180 6870 3190
rect 6760 3170 6770 3180
rect 6730 3160 6770 3170
rect 6590 3130 6660 3140
rect 6590 3110 6595 3130
rect 6615 3110 6635 3130
rect 6655 3110 6660 3130
rect 6590 3080 6660 3110
rect 6590 3060 6595 3080
rect 6615 3060 6635 3080
rect 6655 3060 6660 3080
rect 6590 3050 6660 3060
rect 6685 3130 6715 3140
rect 6685 3110 6690 3130
rect 6710 3110 6715 3130
rect 6685 3080 6715 3110
rect 6685 3060 6690 3080
rect 6710 3060 6715 3080
rect 6685 3050 6715 3060
rect 6740 3130 6770 3140
rect 6740 3110 6745 3130
rect 6765 3110 6770 3130
rect 6740 3080 6770 3110
rect 6740 3060 6745 3080
rect 6765 3060 6770 3080
rect 6740 3050 6770 3060
rect 6635 2975 6655 3050
rect 6745 2975 6765 3050
rect 6850 3030 6870 3180
rect 6950 3140 6970 3220
rect 6990 3230 7215 3240
rect 6990 3210 7000 3230
rect 7020 3220 7215 3230
rect 7020 3210 7030 3220
rect 6990 3200 7030 3210
rect 7135 3140 7155 3220
rect 7300 3200 7320 3430
rect 7340 3420 7345 3430
rect 7365 3420 7370 3440
rect 7340 3390 7370 3420
rect 7340 3370 7345 3390
rect 7365 3370 7370 3390
rect 7340 3340 7370 3370
rect 7340 3320 7345 3340
rect 7365 3320 7370 3340
rect 7340 3290 7370 3320
rect 7340 3270 7345 3290
rect 7365 3270 7370 3290
rect 7340 3260 7370 3270
rect 7395 3440 7425 3450
rect 7395 3420 7400 3440
rect 7420 3420 7425 3440
rect 7395 3390 7425 3420
rect 7395 3370 7400 3390
rect 7420 3370 7425 3390
rect 7395 3340 7425 3370
rect 7395 3320 7400 3340
rect 7420 3320 7425 3340
rect 7395 3290 7425 3320
rect 7395 3270 7400 3290
rect 7420 3270 7425 3290
rect 7395 3260 7425 3270
rect 7450 3440 7520 3450
rect 7450 3420 7455 3440
rect 7475 3420 7495 3440
rect 7515 3420 7520 3440
rect 7450 3390 7520 3420
rect 7450 3370 7455 3390
rect 7475 3370 7495 3390
rect 7515 3370 7520 3390
rect 7450 3340 7520 3370
rect 7450 3320 7455 3340
rect 7475 3320 7495 3340
rect 7515 3320 7520 3340
rect 7450 3290 7520 3320
rect 7450 3270 7455 3290
rect 7475 3270 7495 3290
rect 7515 3270 7520 3290
rect 7450 3260 7520 3270
rect 7560 3440 7630 3450
rect 7560 3420 7565 3440
rect 7585 3420 7605 3440
rect 7625 3420 7630 3440
rect 7560 3390 7630 3420
rect 7560 3370 7565 3390
rect 7585 3370 7605 3390
rect 7625 3370 7630 3390
rect 7560 3340 7630 3370
rect 7560 3320 7565 3340
rect 7585 3320 7605 3340
rect 7625 3320 7630 3340
rect 7560 3290 7630 3320
rect 7560 3270 7565 3290
rect 7585 3270 7605 3290
rect 7625 3270 7630 3290
rect 7560 3260 7630 3270
rect 7655 3440 7685 3450
rect 7655 3420 7660 3440
rect 7680 3420 7685 3440
rect 7655 3390 7685 3420
rect 7655 3370 7660 3390
rect 7680 3370 7685 3390
rect 7655 3340 7685 3370
rect 7655 3320 7660 3340
rect 7680 3320 7685 3340
rect 7655 3290 7685 3320
rect 7655 3270 7660 3290
rect 7680 3270 7685 3290
rect 7655 3260 7685 3270
rect 7710 3440 7740 3450
rect 7710 3420 7715 3440
rect 7735 3420 7740 3440
rect 7710 3390 7740 3420
rect 7710 3370 7715 3390
rect 7735 3370 7740 3390
rect 7710 3340 7740 3370
rect 7710 3320 7715 3340
rect 7735 3320 7740 3340
rect 7710 3290 7740 3320
rect 7710 3270 7715 3290
rect 7735 3270 7740 3290
rect 7710 3260 7740 3270
rect 7780 3440 7850 3450
rect 7780 3420 7785 3440
rect 7805 3420 7825 3440
rect 7845 3420 7850 3440
rect 7780 3390 7850 3420
rect 7780 3370 7785 3390
rect 7805 3370 7825 3390
rect 7845 3370 7850 3390
rect 7780 3340 7850 3370
rect 7780 3320 7785 3340
rect 7805 3320 7825 3340
rect 7845 3320 7850 3340
rect 7780 3290 7850 3320
rect 7780 3270 7785 3290
rect 7805 3270 7825 3290
rect 7845 3270 7850 3290
rect 7780 3260 7850 3270
rect 7875 3440 7905 3450
rect 7875 3420 7880 3440
rect 7900 3420 7905 3440
rect 7875 3390 7905 3420
rect 7875 3370 7880 3390
rect 7900 3370 7905 3390
rect 7875 3340 7905 3370
rect 7875 3320 7880 3340
rect 7900 3320 7905 3340
rect 7875 3290 7905 3320
rect 7875 3270 7880 3290
rect 7900 3270 7905 3290
rect 7875 3260 7905 3270
rect 7945 3440 8015 3450
rect 7945 3420 7950 3440
rect 7970 3420 7990 3440
rect 8010 3420 8015 3440
rect 7945 3390 8015 3420
rect 7945 3370 7950 3390
rect 7970 3370 7990 3390
rect 8010 3370 8015 3390
rect 7945 3340 8015 3370
rect 7945 3320 7950 3340
rect 7970 3320 7990 3340
rect 8010 3320 8015 3340
rect 7945 3290 8015 3320
rect 7945 3270 7950 3290
rect 7970 3270 7990 3290
rect 8010 3270 8015 3290
rect 7945 3260 8015 3270
rect 8040 3440 8070 3450
rect 8040 3420 8045 3440
rect 8065 3420 8070 3440
rect 8040 3390 8070 3420
rect 8040 3370 8045 3390
rect 8065 3370 8070 3390
rect 8040 3340 8070 3370
rect 8040 3320 8045 3340
rect 8065 3320 8070 3340
rect 8040 3290 8070 3320
rect 8040 3270 8045 3290
rect 8065 3270 8070 3290
rect 8040 3260 8070 3270
rect 8145 3440 8235 3450
rect 8145 3420 8155 3440
rect 8175 3420 8205 3440
rect 8225 3420 8235 3440
rect 8145 3390 8235 3420
rect 8145 3370 8155 3390
rect 8175 3370 8205 3390
rect 8225 3370 8235 3390
rect 8145 3340 8235 3370
rect 8145 3320 8155 3340
rect 8175 3320 8205 3340
rect 8225 3320 8235 3340
rect 8145 3290 8235 3320
rect 8145 3270 8155 3290
rect 8175 3270 8205 3290
rect 8225 3270 8235 3290
rect 8145 3260 8235 3270
rect 8260 3440 8300 3450
rect 8260 3420 8270 3440
rect 8290 3420 8300 3440
rect 8260 3390 8300 3420
rect 8260 3370 8270 3390
rect 8290 3370 8300 3390
rect 8260 3340 8300 3370
rect 8260 3320 8270 3340
rect 8290 3320 8300 3340
rect 8260 3290 8300 3320
rect 8260 3270 8270 3290
rect 8290 3270 8300 3290
rect 8260 3260 8300 3270
rect 8340 3440 8430 3450
rect 8340 3420 8350 3440
rect 8370 3420 8400 3440
rect 8420 3420 8430 3440
rect 8340 3390 8430 3420
rect 8340 3370 8350 3390
rect 8370 3370 8400 3390
rect 8420 3370 8430 3390
rect 8340 3340 8430 3370
rect 8340 3320 8350 3340
rect 8370 3320 8400 3340
rect 8420 3320 8430 3340
rect 8340 3290 8430 3320
rect 8340 3270 8350 3290
rect 8370 3270 8400 3290
rect 8420 3270 8430 3290
rect 8340 3260 8430 3270
rect 8455 3440 8495 3450
rect 8455 3420 8465 3440
rect 8485 3420 8495 3440
rect 8455 3390 8495 3420
rect 8455 3370 8465 3390
rect 8485 3370 8495 3390
rect 8455 3340 8495 3370
rect 8455 3320 8465 3340
rect 8485 3320 8495 3340
rect 8455 3290 8495 3320
rect 8455 3270 8465 3290
rect 8485 3270 8495 3290
rect 8455 3260 8495 3270
rect 8535 3440 8625 3450
rect 8535 3420 8545 3440
rect 8565 3420 8595 3440
rect 8615 3420 8625 3440
rect 8535 3390 8625 3420
rect 8535 3370 8545 3390
rect 8565 3370 8595 3390
rect 8615 3370 8625 3390
rect 8535 3340 8625 3370
rect 8535 3320 8545 3340
rect 8565 3320 8595 3340
rect 8615 3320 8625 3340
rect 8535 3290 8625 3320
rect 8535 3270 8545 3290
rect 8565 3270 8595 3290
rect 8615 3270 8625 3290
rect 8535 3260 8625 3270
rect 8650 3440 8690 3450
rect 8650 3420 8660 3440
rect 8680 3420 8690 3440
rect 8650 3390 8690 3420
rect 8650 3370 8660 3390
rect 8680 3370 8690 3390
rect 8650 3340 8690 3370
rect 8650 3320 8660 3340
rect 8680 3320 8690 3340
rect 8650 3290 8690 3320
rect 8650 3270 8660 3290
rect 8680 3270 8690 3290
rect 8650 3260 8690 3270
rect 8730 3440 8770 3450
rect 8730 3420 8740 3440
rect 8760 3420 8770 3440
rect 8730 3390 8770 3420
rect 8730 3370 8740 3390
rect 8760 3370 8770 3390
rect 8730 3340 8770 3370
rect 8730 3320 8740 3340
rect 8760 3320 8770 3340
rect 8730 3290 8770 3320
rect 8730 3270 8740 3290
rect 8760 3270 8770 3290
rect 8730 3260 8770 3270
rect 8795 3440 8835 3450
rect 8795 3420 8805 3440
rect 8825 3420 8835 3440
rect 8795 3390 8835 3420
rect 8795 3370 8805 3390
rect 8825 3370 8835 3390
rect 8795 3340 8835 3370
rect 8795 3320 8805 3340
rect 8825 3320 8835 3340
rect 8795 3290 8835 3320
rect 8795 3270 8805 3290
rect 8825 3270 8835 3290
rect 8795 3260 8835 3270
rect 8875 3440 8965 3450
rect 8875 3420 8885 3440
rect 8905 3420 8935 3440
rect 8955 3420 8965 3440
rect 8875 3390 8965 3420
rect 8875 3370 8885 3390
rect 8905 3370 8935 3390
rect 8955 3370 8965 3390
rect 8875 3340 8965 3370
rect 8875 3320 8885 3340
rect 8905 3320 8935 3340
rect 8955 3320 8965 3340
rect 8875 3290 8965 3320
rect 8875 3270 8885 3290
rect 8905 3270 8935 3290
rect 8955 3270 8965 3290
rect 8875 3260 8965 3270
rect 8990 3440 9030 3450
rect 8990 3420 9000 3440
rect 9020 3420 9030 3440
rect 8990 3390 9030 3420
rect 8990 3370 9000 3390
rect 9020 3370 9030 3390
rect 8990 3340 9030 3370
rect 8990 3320 9000 3340
rect 9020 3320 9030 3340
rect 8990 3290 9030 3320
rect 8990 3270 9000 3290
rect 9020 3270 9030 3290
rect 9720 3435 9730 3455
rect 9750 3435 9780 3455
rect 9800 3435 9810 3455
rect 9720 3405 9810 3435
rect 9720 3385 9730 3405
rect 9750 3385 9780 3405
rect 9800 3385 9810 3405
rect 9720 3355 9810 3385
rect 9720 3335 9730 3355
rect 9750 3335 9780 3355
rect 9800 3335 9810 3355
rect 9720 3305 9810 3335
rect 9720 3285 9730 3305
rect 9750 3285 9780 3305
rect 9800 3285 9810 3305
rect 9720 3275 9810 3285
rect 9880 3455 9920 3465
rect 9880 3435 9890 3455
rect 9910 3435 9920 3455
rect 9880 3405 9920 3435
rect 9880 3385 9890 3405
rect 9910 3385 9920 3405
rect 9880 3355 9920 3385
rect 9880 3335 9890 3355
rect 9910 3335 9920 3355
rect 9880 3305 9920 3335
rect 9880 3285 9890 3305
rect 9910 3285 9920 3305
rect 9880 3275 9920 3285
rect 9990 3455 10030 3465
rect 9990 3435 10000 3455
rect 10020 3435 10030 3455
rect 9990 3405 10030 3435
rect 9990 3385 10000 3405
rect 10020 3385 10030 3405
rect 9990 3355 10030 3385
rect 9990 3335 10000 3355
rect 10020 3335 10030 3355
rect 9990 3305 10030 3335
rect 9990 3285 10000 3305
rect 10020 3285 10030 3305
rect 9990 3275 10030 3285
rect 10100 3455 10140 3465
rect 10100 3435 10110 3455
rect 10130 3435 10140 3455
rect 10100 3405 10140 3435
rect 10100 3385 10110 3405
rect 10130 3385 10140 3405
rect 10100 3355 10140 3385
rect 10100 3335 10110 3355
rect 10130 3335 10140 3355
rect 10100 3305 10140 3335
rect 10100 3285 10110 3305
rect 10130 3285 10140 3305
rect 10100 3275 10140 3285
rect 10210 3455 10250 3465
rect 10210 3435 10220 3455
rect 10240 3435 10250 3455
rect 10210 3405 10250 3435
rect 10210 3385 10220 3405
rect 10240 3385 10250 3405
rect 10210 3355 10250 3385
rect 10210 3335 10220 3355
rect 10240 3335 10250 3355
rect 10210 3305 10250 3335
rect 10210 3285 10220 3305
rect 10240 3285 10250 3305
rect 10210 3275 10250 3285
rect 10320 3455 10360 3465
rect 10320 3435 10330 3455
rect 10350 3435 10360 3455
rect 10320 3405 10360 3435
rect 10320 3385 10330 3405
rect 10350 3385 10360 3405
rect 10320 3355 10360 3385
rect 10320 3335 10330 3355
rect 10350 3335 10360 3355
rect 10320 3305 10360 3335
rect 10320 3285 10330 3305
rect 10350 3285 10360 3305
rect 10320 3275 10360 3285
rect 10430 3455 10570 3465
rect 10430 3435 10440 3455
rect 10460 3435 10490 3455
rect 10510 3435 10540 3455
rect 10560 3435 10570 3455
rect 10430 3405 10570 3435
rect 10430 3385 10440 3405
rect 10460 3385 10490 3405
rect 10510 3385 10540 3405
rect 10560 3385 10570 3405
rect 10430 3355 10570 3385
rect 10430 3335 10440 3355
rect 10460 3335 10490 3355
rect 10510 3335 10540 3355
rect 10560 3335 10570 3355
rect 10430 3305 10570 3335
rect 10430 3285 10440 3305
rect 10460 3285 10490 3305
rect 10510 3285 10540 3305
rect 10560 3285 10570 3305
rect 10430 3275 10570 3285
rect 10640 3455 10680 3465
rect 10640 3435 10650 3455
rect 10670 3435 10680 3455
rect 10640 3405 10680 3435
rect 10640 3385 10650 3405
rect 10670 3385 10680 3405
rect 10640 3355 10680 3385
rect 10640 3335 10650 3355
rect 10670 3335 10680 3355
rect 10640 3305 10680 3335
rect 10640 3285 10650 3305
rect 10670 3285 10680 3305
rect 10640 3275 10680 3285
rect 10750 3455 10790 3465
rect 10750 3435 10760 3455
rect 10780 3435 10790 3455
rect 10750 3405 10790 3435
rect 10750 3385 10760 3405
rect 10780 3385 10790 3405
rect 10750 3355 10790 3385
rect 10750 3335 10760 3355
rect 10780 3335 10790 3355
rect 10750 3305 10790 3335
rect 10750 3285 10760 3305
rect 10780 3285 10790 3305
rect 10750 3275 10790 3285
rect 10860 3455 10900 3465
rect 10860 3435 10870 3455
rect 10890 3435 10900 3455
rect 10860 3405 10900 3435
rect 10860 3385 10870 3405
rect 10890 3385 10900 3405
rect 10860 3355 10900 3385
rect 10860 3335 10870 3355
rect 10890 3335 10900 3355
rect 10860 3305 10900 3335
rect 10860 3285 10870 3305
rect 10890 3285 10900 3305
rect 10860 3275 10900 3285
rect 10970 3455 11010 3465
rect 10970 3435 10980 3455
rect 11000 3435 11010 3455
rect 10970 3405 11010 3435
rect 10970 3385 10980 3405
rect 11000 3385 11010 3405
rect 10970 3355 11010 3385
rect 10970 3335 10980 3355
rect 11000 3335 11010 3355
rect 10970 3305 11010 3335
rect 10970 3285 10980 3305
rect 11000 3285 11010 3305
rect 10970 3275 11010 3285
rect 11080 3455 11120 3465
rect 11080 3435 11090 3455
rect 11110 3435 11120 3455
rect 11080 3405 11120 3435
rect 11080 3385 11090 3405
rect 11110 3385 11120 3405
rect 11080 3355 11120 3385
rect 11080 3335 11090 3355
rect 11110 3335 11120 3355
rect 11080 3305 11120 3335
rect 11080 3285 11090 3305
rect 11110 3285 11120 3305
rect 11080 3275 11120 3285
rect 11190 3455 11280 3465
rect 11190 3435 11200 3455
rect 11220 3435 11250 3455
rect 11270 3435 11280 3455
rect 11190 3405 11280 3435
rect 11190 3385 11200 3405
rect 11220 3385 11250 3405
rect 11270 3385 11280 3405
rect 11190 3355 11280 3385
rect 11190 3335 11200 3355
rect 11220 3335 11250 3355
rect 11270 3335 11280 3355
rect 11190 3305 11280 3335
rect 11190 3285 11200 3305
rect 11220 3285 11250 3305
rect 11270 3285 11280 3305
rect 11190 3275 11280 3285
rect 8990 3260 9030 3270
rect 7345 3240 7365 3260
rect 7345 3220 7420 3240
rect 7180 3190 7320 3200
rect 7180 3170 7190 3190
rect 7210 3180 7320 3190
rect 7210 3170 7220 3180
rect 7180 3160 7220 3170
rect 7400 3140 7420 3220
rect 7660 3225 7680 3260
rect 7885 3225 7905 3260
rect 8050 3225 8070 3260
rect 7660 3215 7770 3225
rect 7660 3205 7740 3215
rect 7515 3195 7555 3205
rect 7515 3175 7525 3195
rect 7545 3175 7555 3195
rect 7515 3165 7555 3175
rect 7715 3195 7740 3205
rect 7760 3195 7770 3215
rect 7715 3185 7770 3195
rect 7885 3215 7935 3225
rect 7885 3195 7905 3215
rect 7925 3195 7935 3215
rect 7885 3185 7935 3195
rect 8050 3215 8100 3225
rect 8050 3195 8070 3215
rect 8090 3195 8100 3215
rect 8280 3215 8300 3260
rect 8410 3215 8450 3225
rect 8050 3185 8100 3195
rect 8125 3200 8165 3210
rect 7715 3140 7735 3185
rect 7885 3140 7905 3185
rect 8050 3140 8070 3185
rect 8125 3180 8135 3200
rect 8155 3180 8165 3200
rect 8125 3170 8165 3180
rect 8280 3195 8420 3215
rect 8440 3195 8450 3215
rect 8280 3140 8300 3195
rect 8410 3185 8450 3195
rect 8475 3200 8495 3260
rect 8670 3240 8690 3260
rect 8670 3230 8710 3240
rect 8670 3210 8680 3230
rect 8700 3210 8710 3230
rect 8670 3200 8710 3210
rect 8475 3190 8645 3200
rect 8475 3180 8615 3190
rect 8475 3140 8495 3180
rect 8605 3170 8615 3180
rect 8635 3170 8645 3190
rect 8605 3160 8645 3170
rect 8670 3140 8690 3200
rect 8740 3140 8760 3260
rect 8805 3180 8825 3260
rect 8845 3230 8885 3240
rect 8845 3210 8855 3230
rect 8875 3210 8885 3230
rect 8845 3200 8885 3210
rect 9000 3200 9020 3260
rect 9770 3245 9810 3255
rect 9770 3225 9780 3245
rect 9800 3225 9810 3245
rect 9770 3215 9810 3225
rect 11190 3245 11230 3255
rect 11190 3225 11200 3245
rect 11220 3225 11230 3245
rect 11190 3215 11230 3225
rect 9000 3190 9040 3200
rect 9000 3180 9010 3190
rect 8805 3170 9010 3180
rect 9030 3170 9040 3190
rect 8805 3160 9040 3170
rect 8805 3140 8825 3160
rect 6890 3130 6920 3140
rect 6890 3110 6895 3130
rect 6915 3110 6920 3130
rect 6890 3080 6920 3110
rect 6890 3060 6895 3080
rect 6915 3060 6920 3080
rect 6890 3050 6920 3060
rect 6945 3130 6975 3140
rect 6945 3110 6950 3130
rect 6970 3110 6975 3130
rect 6945 3080 6975 3110
rect 6945 3060 6950 3080
rect 6970 3060 6975 3080
rect 6945 3050 6975 3060
rect 7000 3130 7110 3140
rect 7000 3110 7005 3130
rect 7025 3110 7045 3130
rect 7065 3110 7085 3130
rect 7105 3110 7110 3130
rect 7000 3080 7110 3110
rect 7000 3060 7005 3080
rect 7025 3060 7045 3080
rect 7065 3060 7085 3080
rect 7105 3060 7110 3080
rect 7000 3050 7110 3060
rect 7135 3130 7165 3140
rect 7135 3110 7140 3130
rect 7160 3110 7165 3130
rect 7135 3080 7165 3110
rect 7135 3060 7140 3080
rect 7160 3060 7165 3080
rect 7135 3050 7165 3060
rect 7190 3130 7220 3140
rect 7190 3110 7195 3130
rect 7215 3110 7220 3130
rect 7190 3080 7220 3110
rect 7190 3060 7195 3080
rect 7215 3060 7220 3080
rect 7190 3050 7220 3060
rect 7340 3130 7370 3140
rect 7340 3110 7345 3130
rect 7365 3110 7370 3130
rect 7340 3080 7370 3110
rect 7340 3060 7345 3080
rect 7365 3060 7370 3080
rect 7340 3050 7370 3060
rect 7395 3130 7425 3140
rect 7395 3110 7400 3130
rect 7420 3110 7425 3130
rect 7395 3080 7425 3110
rect 7395 3060 7400 3080
rect 7420 3060 7425 3080
rect 7395 3050 7425 3060
rect 7450 3130 7520 3140
rect 7450 3110 7455 3130
rect 7475 3110 7495 3130
rect 7515 3110 7520 3130
rect 7450 3080 7520 3110
rect 7450 3060 7455 3080
rect 7475 3060 7495 3080
rect 7515 3060 7520 3080
rect 7450 3050 7520 3060
rect 7560 3130 7630 3140
rect 7560 3110 7565 3130
rect 7585 3110 7605 3130
rect 7625 3110 7630 3130
rect 7560 3080 7630 3110
rect 7560 3060 7565 3080
rect 7585 3060 7605 3080
rect 7625 3060 7630 3080
rect 7560 3050 7630 3060
rect 7655 3130 7685 3140
rect 7655 3110 7660 3130
rect 7680 3110 7685 3130
rect 7655 3080 7685 3110
rect 7655 3060 7660 3080
rect 7680 3060 7685 3080
rect 7655 3050 7685 3060
rect 7710 3130 7740 3140
rect 7710 3110 7715 3130
rect 7735 3110 7740 3130
rect 7710 3080 7740 3110
rect 7710 3060 7715 3080
rect 7735 3060 7740 3080
rect 7710 3050 7740 3060
rect 7780 3130 7850 3140
rect 7780 3110 7785 3130
rect 7805 3110 7825 3130
rect 7845 3110 7850 3130
rect 7780 3080 7850 3110
rect 7780 3060 7785 3080
rect 7805 3060 7825 3080
rect 7845 3060 7850 3080
rect 7780 3050 7850 3060
rect 7875 3130 7905 3140
rect 7875 3110 7880 3130
rect 7900 3110 7905 3130
rect 7875 3080 7905 3110
rect 7875 3060 7880 3080
rect 7900 3060 7905 3080
rect 7875 3050 7905 3060
rect 7945 3130 8015 3140
rect 7945 3110 7950 3130
rect 7970 3110 7990 3130
rect 8010 3110 8015 3130
rect 7945 3080 8015 3110
rect 7945 3060 7950 3080
rect 7970 3060 7990 3080
rect 8010 3060 8015 3080
rect 7945 3050 8015 3060
rect 8040 3130 8070 3140
rect 8040 3110 8045 3130
rect 8065 3110 8070 3130
rect 8040 3080 8070 3110
rect 8040 3060 8045 3080
rect 8065 3060 8070 3080
rect 8040 3050 8070 3060
rect 8155 3130 8235 3140
rect 8155 3110 8160 3130
rect 8180 3110 8205 3130
rect 8225 3110 8235 3130
rect 8155 3080 8235 3110
rect 8155 3060 8160 3080
rect 8180 3060 8205 3080
rect 8225 3060 8235 3080
rect 8155 3050 8235 3060
rect 8260 3130 8300 3140
rect 8260 3110 8270 3130
rect 8290 3110 8300 3130
rect 8260 3080 8300 3110
rect 8260 3060 8270 3080
rect 8290 3060 8300 3080
rect 8260 3050 8300 3060
rect 8350 3130 8430 3140
rect 8350 3110 8355 3130
rect 8375 3110 8400 3130
rect 8420 3110 8430 3130
rect 8350 3080 8430 3110
rect 8350 3060 8355 3080
rect 8375 3060 8400 3080
rect 8420 3060 8430 3080
rect 8350 3050 8430 3060
rect 8455 3130 8495 3140
rect 8455 3110 8465 3130
rect 8485 3110 8495 3130
rect 8455 3080 8495 3110
rect 8455 3060 8465 3080
rect 8485 3060 8495 3080
rect 8455 3050 8495 3060
rect 8545 3130 8625 3140
rect 8545 3110 8550 3130
rect 8570 3110 8595 3130
rect 8615 3110 8625 3130
rect 8545 3080 8625 3110
rect 8545 3060 8550 3080
rect 8570 3060 8595 3080
rect 8615 3060 8625 3080
rect 8545 3050 8625 3060
rect 8650 3130 8690 3140
rect 8650 3110 8660 3130
rect 8680 3110 8690 3130
rect 8650 3080 8690 3110
rect 8650 3060 8660 3080
rect 8680 3060 8690 3080
rect 8650 3050 8690 3060
rect 8730 3130 8770 3140
rect 8730 3110 8740 3130
rect 8760 3110 8770 3130
rect 8730 3080 8770 3110
rect 8730 3060 8740 3080
rect 8760 3060 8770 3080
rect 8730 3050 8770 3060
rect 8795 3130 8835 3140
rect 8795 3110 8805 3130
rect 8825 3110 8835 3130
rect 8795 3080 8835 3110
rect 8795 3060 8805 3080
rect 8825 3060 8835 3080
rect 8795 3050 8835 3060
rect 6830 3020 6870 3030
rect 6830 3000 6840 3020
rect 6860 3000 6870 3020
rect 6830 2990 6870 3000
rect 6895 2975 6915 3050
rect 7005 2975 7025 3050
rect 7085 2975 7105 3050
rect 7195 2975 7215 3050
rect 7345 2975 7365 3050
rect 7455 2975 7475 3050
rect 7605 2975 7625 3050
rect 7690 3020 7730 3030
rect 7690 3000 7700 3020
rect 7720 3000 7730 3020
rect 7690 2990 7730 3000
rect 7825 2975 7845 3050
rect 7990 2975 8010 3050
rect 8205 2975 8225 3050
rect 8400 2975 8420 3050
rect 8595 2975 8615 3050
rect 8740 3030 8760 3050
rect 8730 3020 8770 3030
rect 8730 3000 8740 3020
rect 8760 3000 8770 3020
rect 8730 2990 8770 3000
rect 6625 2965 6665 2975
rect 6625 2945 6635 2965
rect 6655 2945 6665 2965
rect 6625 2935 6665 2945
rect 6735 2965 6775 2975
rect 6735 2945 6745 2965
rect 6765 2945 6775 2965
rect 6735 2935 6775 2945
rect 6885 2965 6925 2975
rect 6885 2945 6895 2965
rect 6915 2945 6925 2965
rect 6885 2935 6925 2945
rect 6995 2965 7035 2975
rect 6995 2945 7005 2965
rect 7025 2945 7035 2965
rect 6995 2935 7035 2945
rect 7075 2965 7115 2975
rect 7075 2945 7085 2965
rect 7105 2945 7115 2965
rect 7075 2935 7115 2945
rect 7185 2965 7225 2975
rect 7185 2945 7195 2965
rect 7215 2945 7225 2965
rect 7185 2935 7225 2945
rect 7335 2965 7375 2975
rect 7335 2945 7345 2965
rect 7365 2945 7375 2965
rect 7335 2935 7375 2945
rect 7445 2965 7485 2975
rect 7445 2945 7455 2965
rect 7475 2945 7485 2965
rect 7445 2935 7485 2945
rect 7595 2965 7635 2975
rect 7595 2945 7605 2965
rect 7625 2945 7635 2965
rect 7595 2935 7635 2945
rect 7815 2965 7855 2975
rect 7815 2945 7825 2965
rect 7845 2945 7855 2965
rect 7815 2935 7855 2945
rect 7980 2965 8020 2975
rect 7980 2945 7990 2965
rect 8010 2945 8020 2965
rect 7980 2935 8020 2945
rect 8195 2965 8235 2975
rect 8195 2945 8205 2965
rect 8225 2945 8235 2965
rect 8195 2935 8235 2945
rect 8390 2965 8430 2975
rect 8390 2945 8400 2965
rect 8420 2945 8430 2965
rect 8390 2935 8430 2945
rect 8585 2965 8625 2975
rect 8585 2945 8595 2965
rect 8615 2945 8625 2965
rect 8585 2935 8625 2945
rect 11490 2940 11545 2950
rect 11490 2905 11500 2940
rect 11535 2905 11545 2940
rect 11490 2895 11545 2905
<< viali >>
rect 11555 4155 11590 4190
rect 6635 4125 6655 4145
rect 6745 4125 6765 4145
rect 6895 4125 6915 4145
rect 7010 4125 7030 4145
rect 7085 4125 7105 4145
rect 7195 4125 7215 4145
rect 7345 4125 7365 4145
rect 7455 4125 7475 4145
rect 7655 4125 7675 4145
rect 7820 4125 7840 4145
rect 7985 4125 8005 4145
rect 8205 4125 8225 4145
rect 8595 4125 8615 4145
rect 8935 4125 8955 4145
rect 8460 4070 8480 4090
rect 8775 4070 8795 4090
rect 9680 4045 9700 4065
rect 11200 4045 11220 4065
rect 9680 3985 9700 4005
rect 6575 3880 6595 3900
rect 7535 3875 7555 3895
rect 8050 3875 8070 3895
rect 8125 3880 8145 3900
rect 9680 3935 9700 3955
rect 9010 3900 9030 3920
rect 9680 3885 9700 3905
rect 9680 3835 9700 3855
rect 9790 3985 9810 4005
rect 9790 3935 9810 3955
rect 9790 3885 9810 3905
rect 9790 3835 9810 3855
rect 9900 3985 9920 4005
rect 9900 3935 9920 3955
rect 9900 3885 9920 3905
rect 9900 3835 9920 3855
rect 10010 3985 10030 4005
rect 10010 3935 10030 3955
rect 10010 3885 10030 3905
rect 10010 3835 10030 3855
rect 10120 3985 10140 4005
rect 10170 3985 10190 4005
rect 10220 3985 10240 4005
rect 10120 3935 10140 3955
rect 10170 3935 10190 3955
rect 10220 3935 10240 3955
rect 10120 3885 10140 3905
rect 10170 3885 10190 3905
rect 10220 3885 10240 3905
rect 10120 3835 10140 3855
rect 10170 3835 10190 3855
rect 10220 3835 10240 3855
rect 10330 3985 10350 4005
rect 10330 3935 10350 3955
rect 10330 3885 10350 3905
rect 10330 3835 10350 3855
rect 10440 3985 10460 4005
rect 10440 3935 10460 3955
rect 10440 3885 10460 3905
rect 10440 3835 10460 3855
rect 10550 3985 10570 4005
rect 10550 3935 10570 3955
rect 10550 3885 10570 3905
rect 10550 3835 10570 3855
rect 10660 3985 10680 4005
rect 10710 3985 10730 4005
rect 10760 3985 10780 4005
rect 10660 3935 10680 3955
rect 10710 3935 10730 3955
rect 10760 3935 10780 3955
rect 10660 3885 10680 3905
rect 10710 3885 10730 3905
rect 10760 3885 10780 3905
rect 10660 3835 10680 3855
rect 10710 3835 10730 3855
rect 10760 3835 10780 3855
rect 10870 3985 10890 4005
rect 10870 3935 10890 3955
rect 10870 3885 10890 3905
rect 10870 3835 10890 3855
rect 10980 3985 11000 4005
rect 10980 3935 11000 3955
rect 10980 3885 11000 3905
rect 10980 3835 11000 3855
rect 11090 3985 11110 4005
rect 11090 3935 11110 3955
rect 11090 3885 11110 3905
rect 11090 3835 11110 3855
rect 11200 3985 11220 4005
rect 11200 3935 11220 3955
rect 11200 3885 11220 3905
rect 11200 3835 11220 3855
rect 9900 3780 9920 3800
rect 10915 3760 10935 3780
rect 11045 3760 11065 3780
rect 11380 3760 11415 3795
rect 6860 3590 6880 3610
rect 8420 3590 8440 3610
rect 8740 3590 8760 3610
rect 6635 3535 6655 3555
rect 7005 3535 7025 3555
rect 7085 3535 7105 3555
rect 7455 3535 7475 3555
rect 7580 3535 7600 3555
rect 7675 3535 7695 3555
rect 7715 3535 7735 3555
rect 7820 3535 7840 3555
rect 7985 3535 8005 3555
rect 8205 3535 8225 3555
rect 8400 3535 8420 3555
rect 8595 3535 8615 3555
rect 8935 3535 8955 3555
rect 7635 3480 7655 3500
rect 10110 3495 10130 3515
rect 10695 3510 10715 3530
rect 11045 3510 11065 3530
rect 11380 3495 11415 3530
rect 6575 3190 6595 3210
rect 9780 3435 9800 3455
rect 9780 3385 9800 3405
rect 9780 3335 9800 3355
rect 9780 3285 9800 3305
rect 9890 3435 9910 3455
rect 9890 3385 9910 3405
rect 9890 3335 9910 3355
rect 9890 3285 9910 3305
rect 10000 3435 10020 3455
rect 10000 3385 10020 3405
rect 10000 3335 10020 3355
rect 10000 3285 10020 3305
rect 10110 3435 10130 3455
rect 10110 3385 10130 3405
rect 10110 3335 10130 3355
rect 10110 3285 10130 3305
rect 10220 3435 10240 3455
rect 10220 3385 10240 3405
rect 10220 3335 10240 3355
rect 10220 3285 10240 3305
rect 10330 3435 10350 3455
rect 10330 3385 10350 3405
rect 10330 3335 10350 3355
rect 10330 3285 10350 3305
rect 10440 3435 10460 3455
rect 10490 3435 10510 3455
rect 10540 3435 10560 3455
rect 10440 3385 10460 3405
rect 10490 3385 10510 3405
rect 10540 3385 10560 3405
rect 10440 3335 10460 3355
rect 10490 3335 10510 3355
rect 10540 3335 10560 3355
rect 10440 3285 10460 3305
rect 10490 3285 10510 3305
rect 10540 3285 10560 3305
rect 10650 3435 10670 3455
rect 10650 3385 10670 3405
rect 10650 3335 10670 3355
rect 10650 3285 10670 3305
rect 10760 3435 10780 3455
rect 10760 3385 10780 3405
rect 10760 3335 10780 3355
rect 10760 3285 10780 3305
rect 10870 3435 10890 3455
rect 10870 3385 10890 3405
rect 10870 3335 10890 3355
rect 10870 3285 10890 3305
rect 10980 3435 11000 3455
rect 10980 3385 11000 3405
rect 10980 3335 11000 3355
rect 10980 3285 11000 3305
rect 11090 3435 11110 3455
rect 11090 3385 11110 3405
rect 11090 3335 11110 3355
rect 11090 3285 11110 3305
rect 11200 3435 11220 3455
rect 11200 3385 11220 3405
rect 11200 3335 11220 3355
rect 11200 3285 11220 3305
rect 7525 3175 7545 3195
rect 8070 3195 8090 3215
rect 8135 3180 8155 3200
rect 8855 3210 8875 3230
rect 9780 3225 9800 3245
rect 11200 3225 11220 3245
rect 9010 3170 9030 3190
rect 6840 3000 6860 3020
rect 7700 3000 7720 3020
rect 8740 3000 8760 3020
rect 6635 2945 6655 2965
rect 6745 2945 6765 2965
rect 6895 2945 6915 2965
rect 7005 2945 7025 2965
rect 7085 2945 7105 2965
rect 7195 2945 7215 2965
rect 7345 2945 7365 2965
rect 7455 2945 7475 2965
rect 7605 2945 7625 2965
rect 7825 2945 7845 2965
rect 7990 2945 8010 2965
rect 8205 2945 8225 2965
rect 8400 2945 8420 2965
rect 8595 2945 8615 2965
rect 11500 2905 11535 2940
<< metal1 >>
rect 11545 4190 11600 4200
rect 9050 4185 9090 4190
rect 9050 4155 9055 4185
rect 9085 4155 9090 4185
rect 6625 4150 6665 4155
rect 6625 4120 6630 4150
rect 6660 4120 6665 4150
rect 6625 4115 6665 4120
rect 6735 4150 6775 4155
rect 6735 4120 6740 4150
rect 6770 4120 6775 4150
rect 6735 4115 6775 4120
rect 6885 4150 6925 4155
rect 6885 4120 6890 4150
rect 6920 4120 6925 4150
rect 6885 4115 6925 4120
rect 7000 4150 7040 4155
rect 7000 4120 7005 4150
rect 7035 4120 7040 4150
rect 7000 4115 7040 4120
rect 7075 4150 7115 4155
rect 7075 4120 7080 4150
rect 7110 4120 7115 4150
rect 7075 4115 7115 4120
rect 7185 4150 7225 4155
rect 7185 4120 7190 4150
rect 7220 4120 7225 4150
rect 7185 4115 7225 4120
rect 7335 4150 7375 4155
rect 7335 4120 7340 4150
rect 7370 4120 7375 4150
rect 7335 4115 7375 4120
rect 7445 4150 7485 4155
rect 7445 4120 7450 4150
rect 7480 4120 7485 4150
rect 7445 4115 7485 4120
rect 7645 4150 7685 4155
rect 7645 4120 7650 4150
rect 7680 4120 7685 4150
rect 7645 4115 7685 4120
rect 7810 4150 7850 4155
rect 7810 4120 7815 4150
rect 7845 4120 7850 4150
rect 7810 4115 7850 4120
rect 7975 4150 8015 4155
rect 7975 4120 7980 4150
rect 8010 4120 8015 4150
rect 7975 4115 8015 4120
rect 8195 4150 8235 4155
rect 8195 4120 8200 4150
rect 8230 4120 8235 4150
rect 8195 4115 8235 4120
rect 8325 4150 8365 4155
rect 8325 4120 8330 4150
rect 8360 4120 8365 4150
rect 8325 4115 8365 4120
rect 8585 4150 8625 4155
rect 8585 4120 8590 4150
rect 8620 4120 8625 4150
rect 8585 4115 8625 4120
rect 8925 4150 8965 4155
rect 8925 4120 8930 4150
rect 8960 4120 8965 4150
rect 8925 4115 8965 4120
rect 6565 3905 6605 3910
rect 6565 3875 6570 3905
rect 6600 3875 6605 3905
rect 6565 3870 6605 3875
rect 7525 3900 7565 3905
rect 7525 3870 7530 3900
rect 7560 3870 7565 3900
rect 7525 3865 7565 3870
rect 8040 3900 8100 3905
rect 8040 3870 8045 3900
rect 8075 3870 8100 3900
rect 8040 3865 8100 3870
rect 6850 3615 6890 3620
rect 6850 3585 6855 3615
rect 6885 3585 6890 3615
rect 6850 3580 6890 3585
rect 6625 3560 6665 3565
rect 6625 3530 6630 3560
rect 6660 3530 6665 3560
rect 6625 3525 6665 3530
rect 6995 3560 7035 3565
rect 6995 3530 7000 3560
rect 7030 3530 7035 3560
rect 6995 3525 7035 3530
rect 7075 3560 7115 3565
rect 7075 3530 7080 3560
rect 7110 3530 7115 3560
rect 7075 3525 7115 3530
rect 7445 3560 7485 3565
rect 7445 3530 7450 3560
rect 7480 3530 7485 3560
rect 7445 3525 7485 3530
rect 6565 3215 6605 3220
rect 6565 3185 6570 3215
rect 6600 3185 6605 3215
rect 7535 3205 7555 3865
rect 7615 3615 7655 3620
rect 7615 3585 7620 3615
rect 7650 3585 7655 3615
rect 7615 3580 7655 3585
rect 7570 3560 7610 3565
rect 7570 3530 7575 3560
rect 7605 3530 7610 3560
rect 7570 3525 7610 3530
rect 7625 3505 7645 3580
rect 7665 3560 7745 3565
rect 7665 3530 7670 3560
rect 7700 3530 7710 3560
rect 7740 3530 7745 3560
rect 7665 3525 7745 3530
rect 7810 3560 7850 3565
rect 7810 3530 7815 3560
rect 7845 3530 7850 3560
rect 7810 3525 7850 3530
rect 7975 3560 8015 3565
rect 7975 3530 7980 3560
rect 8010 3530 8015 3560
rect 7975 3525 8015 3530
rect 7625 3475 7630 3505
rect 7660 3475 7665 3505
rect 7625 3470 7665 3475
rect 8080 3225 8100 3865
rect 8115 3900 8155 3910
rect 8115 3880 8125 3900
rect 8145 3880 8155 3900
rect 8115 3870 8155 3880
rect 8115 3625 8135 3870
rect 8115 3620 8155 3625
rect 8115 3590 8120 3620
rect 8150 3590 8155 3620
rect 8335 3615 8355 4115
rect 8450 4095 8525 4100
rect 8450 4065 8455 4095
rect 8485 4065 8525 4095
rect 8450 4060 8525 4065
rect 8765 4095 8805 4100
rect 8765 4065 8770 4095
rect 8800 4065 8805 4095
rect 8765 4060 8805 4065
rect 9050 4095 9090 4155
rect 11545 4155 11555 4190
rect 11590 4155 11600 4190
rect 11545 4145 11600 4155
rect 9050 4065 9055 4095
rect 9085 4065 9090 4095
rect 9050 4060 9090 4065
rect 9670 4115 9710 4120
rect 9670 4085 9675 4115
rect 9705 4085 9710 4115
rect 9670 4065 9710 4085
rect 8410 3615 8450 3620
rect 8115 3585 8155 3590
rect 8325 3585 8330 3615
rect 8360 3585 8365 3615
rect 8410 3585 8415 3615
rect 8445 3585 8450 3615
rect 8505 3565 8525 4060
rect 9670 4045 9680 4065
rect 9700 4045 9710 4065
rect 9670 4005 9710 4045
rect 9670 3985 9680 4005
rect 9700 3985 9710 4005
rect 9670 3955 9710 3985
rect 9670 3935 9680 3955
rect 9700 3935 9710 3955
rect 9000 3925 9040 3930
rect 9000 3895 9005 3925
rect 9035 3895 9040 3925
rect 9000 3890 9040 3895
rect 9090 3925 9130 3930
rect 9090 3895 9095 3925
rect 9125 3895 9130 3925
rect 9090 3745 9130 3895
rect 9670 3905 9710 3935
rect 9670 3885 9680 3905
rect 9700 3885 9710 3905
rect 9670 3855 9710 3885
rect 9670 3835 9680 3855
rect 9700 3835 9710 3855
rect 9670 3825 9710 3835
rect 9780 4115 9820 4120
rect 9780 4085 9785 4115
rect 9815 4085 9820 4115
rect 9780 4005 9820 4085
rect 10000 4115 10040 4120
rect 10000 4085 10005 4115
rect 10035 4085 10040 4115
rect 9780 3985 9790 4005
rect 9810 3985 9820 4005
rect 9780 3955 9820 3985
rect 9780 3935 9790 3955
rect 9810 3935 9820 3955
rect 9780 3905 9820 3935
rect 9780 3885 9790 3905
rect 9810 3885 9820 3905
rect 9780 3855 9820 3885
rect 9780 3835 9790 3855
rect 9810 3835 9820 3855
rect 9780 3825 9820 3835
rect 9890 4005 9930 4015
rect 9890 3985 9900 4005
rect 9920 3985 9930 4005
rect 9890 3955 9930 3985
rect 9890 3935 9900 3955
rect 9920 3935 9930 3955
rect 9890 3905 9930 3935
rect 9890 3885 9900 3905
rect 9920 3885 9930 3905
rect 9890 3855 9930 3885
rect 9890 3835 9900 3855
rect 9920 3835 9930 3855
rect 9890 3825 9930 3835
rect 10000 4005 10040 4085
rect 10160 4115 10200 4120
rect 10160 4085 10165 4115
rect 10195 4085 10200 4115
rect 10160 4015 10200 4085
rect 10320 4115 10360 4120
rect 10320 4085 10325 4115
rect 10355 4085 10360 4115
rect 10000 3985 10010 4005
rect 10030 3985 10040 4005
rect 10000 3955 10040 3985
rect 10000 3935 10010 3955
rect 10030 3935 10040 3955
rect 10000 3905 10040 3935
rect 10000 3885 10010 3905
rect 10030 3885 10040 3905
rect 10000 3855 10040 3885
rect 10000 3835 10010 3855
rect 10030 3835 10040 3855
rect 10000 3825 10040 3835
rect 10110 4005 10250 4015
rect 10110 3985 10120 4005
rect 10140 3985 10170 4005
rect 10190 3985 10220 4005
rect 10240 3985 10250 4005
rect 10110 3955 10250 3985
rect 10110 3935 10120 3955
rect 10140 3935 10170 3955
rect 10190 3935 10220 3955
rect 10240 3935 10250 3955
rect 10110 3905 10250 3935
rect 10110 3885 10120 3905
rect 10140 3885 10170 3905
rect 10190 3885 10220 3905
rect 10240 3885 10250 3905
rect 10110 3855 10250 3885
rect 10110 3835 10120 3855
rect 10140 3835 10170 3855
rect 10190 3835 10220 3855
rect 10240 3835 10250 3855
rect 10110 3825 10250 3835
rect 10320 4005 10360 4085
rect 10540 4115 10580 4120
rect 10540 4085 10545 4115
rect 10575 4085 10580 4115
rect 10320 3985 10330 4005
rect 10350 3985 10360 4005
rect 10320 3955 10360 3985
rect 10320 3935 10330 3955
rect 10350 3935 10360 3955
rect 10320 3905 10360 3935
rect 10320 3885 10330 3905
rect 10350 3885 10360 3905
rect 10320 3855 10360 3885
rect 10320 3835 10330 3855
rect 10350 3835 10360 3855
rect 10320 3825 10360 3835
rect 10430 4005 10470 4015
rect 10430 3985 10440 4005
rect 10460 3985 10470 4005
rect 10430 3955 10470 3985
rect 10430 3935 10440 3955
rect 10460 3935 10470 3955
rect 10430 3905 10470 3935
rect 10430 3885 10440 3905
rect 10460 3885 10470 3905
rect 10430 3855 10470 3885
rect 10430 3835 10440 3855
rect 10460 3835 10470 3855
rect 9090 3715 9095 3745
rect 9125 3715 9130 3745
rect 9090 3710 9130 3715
rect 9890 3800 9930 3810
rect 9890 3780 9900 3800
rect 9920 3780 9930 3800
rect 9090 3690 9130 3695
rect 9090 3660 9095 3690
rect 9125 3660 9130 3690
rect 8730 3615 8770 3620
rect 8730 3585 8735 3615
rect 8765 3585 8770 3615
rect 8730 3580 8770 3585
rect 9090 3615 9130 3660
rect 9890 3690 9930 3780
rect 9890 3660 9895 3690
rect 9925 3660 9930 3690
rect 9890 3655 9930 3660
rect 9090 3585 9095 3615
rect 9125 3585 9130 3615
rect 9090 3580 9130 3585
rect 9145 3635 9185 3640
rect 9145 3605 9150 3635
rect 9180 3605 9185 3635
rect 8195 3560 8235 3565
rect 8195 3530 8200 3560
rect 8230 3530 8235 3560
rect 8195 3525 8235 3530
rect 8390 3560 8430 3565
rect 8390 3530 8395 3560
rect 8425 3530 8430 3560
rect 8390 3525 8430 3530
rect 8495 3560 8535 3565
rect 8495 3530 8500 3560
rect 8530 3530 8535 3560
rect 8495 3525 8535 3530
rect 8585 3560 8625 3565
rect 8585 3530 8590 3560
rect 8620 3530 8625 3560
rect 8585 3525 8625 3530
rect 8925 3560 8965 3565
rect 8925 3530 8930 3560
rect 8960 3530 8965 3560
rect 8925 3525 8965 3530
rect 6565 3180 6605 3185
rect 7515 3200 7555 3205
rect 7515 3170 7520 3200
rect 7550 3170 7555 3200
rect 8060 3220 8100 3225
rect 8060 3190 8065 3220
rect 8095 3190 8100 3220
rect 8845 3235 8885 3240
rect 8060 3185 8100 3190
rect 8125 3200 8165 3210
rect 7515 3165 7555 3170
rect 8125 3180 8135 3200
rect 8155 3180 8165 3200
rect 8125 3170 8165 3180
rect 8845 3205 8850 3235
rect 8880 3205 8885 3235
rect 8125 3040 8145 3170
rect 8115 3035 8155 3040
rect 6830 3025 6870 3030
rect 6830 2995 6835 3025
rect 6865 2995 6870 3025
rect 6830 2990 6870 2995
rect 7690 3025 7730 3030
rect 7690 2995 7695 3025
rect 7725 2995 7730 3025
rect 8115 3005 8120 3035
rect 8150 3005 8155 3035
rect 8115 3000 8155 3005
rect 8730 3025 8770 3030
rect 7690 2990 7730 2995
rect 8730 2995 8735 3025
rect 8765 2995 8770 3025
rect 8730 2990 8770 2995
rect 6625 2970 6665 2975
rect 6625 2940 6630 2970
rect 6660 2940 6665 2970
rect 6625 2935 6665 2940
rect 6735 2970 6775 2975
rect 6735 2940 6740 2970
rect 6770 2940 6775 2970
rect 6735 2935 6775 2940
rect 6885 2970 6925 2975
rect 6885 2940 6890 2970
rect 6920 2940 6925 2970
rect 6885 2935 6925 2940
rect 6995 2970 7035 2975
rect 6995 2940 7000 2970
rect 7030 2940 7035 2970
rect 6995 2935 7035 2940
rect 7075 2970 7115 2975
rect 7075 2940 7080 2970
rect 7110 2940 7115 2970
rect 7075 2935 7115 2940
rect 7185 2970 7225 2975
rect 7185 2940 7190 2970
rect 7220 2940 7225 2970
rect 7185 2935 7225 2940
rect 7335 2970 7375 2975
rect 7335 2940 7340 2970
rect 7370 2940 7375 2970
rect 7335 2935 7375 2940
rect 7445 2970 7485 2975
rect 7445 2940 7450 2970
rect 7480 2940 7485 2970
rect 7445 2935 7485 2940
rect 7595 2970 7635 2975
rect 7595 2940 7600 2970
rect 7630 2940 7635 2970
rect 7595 2935 7635 2940
rect 7815 2970 7855 2975
rect 7815 2940 7820 2970
rect 7850 2940 7855 2970
rect 7815 2935 7855 2940
rect 7980 2970 8020 2975
rect 7980 2940 7985 2970
rect 8015 2940 8020 2970
rect 7980 2935 8020 2940
rect 8195 2970 8235 2975
rect 8195 2940 8200 2970
rect 8230 2940 8235 2970
rect 8195 2935 8235 2940
rect 8390 2970 8430 2975
rect 8390 2940 8395 2970
rect 8425 2940 8430 2970
rect 8390 2935 8430 2940
rect 8585 2970 8625 2975
rect 8585 2940 8590 2970
rect 8620 2940 8625 2970
rect 8585 2935 8625 2940
rect 8845 2940 8885 3205
rect 9000 3195 9040 3200
rect 9000 3165 9005 3195
rect 9035 3165 9040 3195
rect 9000 3160 9040 3165
rect 9145 3195 9185 3605
rect 9145 3165 9150 3195
rect 9180 3165 9185 3195
rect 9145 3160 9185 3165
rect 9200 3580 9240 3585
rect 9200 3550 9205 3580
rect 9235 3550 9240 3580
rect 9200 3025 9240 3550
rect 10100 3580 10140 3585
rect 10100 3550 10105 3580
rect 10135 3550 10140 3580
rect 9990 3520 10030 3525
rect 9990 3490 9995 3520
rect 10025 3490 10030 3520
rect 9770 3455 9810 3465
rect 9770 3435 9780 3455
rect 9800 3435 9810 3455
rect 9770 3405 9810 3435
rect 9770 3385 9780 3405
rect 9800 3385 9810 3405
rect 9770 3355 9810 3385
rect 9770 3335 9780 3355
rect 9800 3335 9810 3355
rect 9770 3305 9810 3335
rect 9770 3285 9780 3305
rect 9800 3285 9810 3305
rect 9770 3245 9810 3285
rect 9770 3225 9780 3245
rect 9800 3225 9810 3245
rect 9770 3195 9810 3225
rect 9770 3165 9775 3195
rect 9805 3165 9810 3195
rect 9770 3160 9810 3165
rect 9880 3455 9920 3465
rect 9880 3435 9890 3455
rect 9910 3435 9920 3455
rect 9880 3405 9920 3435
rect 9880 3385 9890 3405
rect 9910 3385 9920 3405
rect 9880 3355 9920 3385
rect 9880 3335 9890 3355
rect 9910 3335 9920 3355
rect 9880 3305 9920 3335
rect 9880 3285 9890 3305
rect 9910 3285 9920 3305
rect 9880 3195 9920 3285
rect 9990 3455 10030 3490
rect 10100 3515 10140 3550
rect 10100 3495 10110 3515
rect 10130 3495 10140 3515
rect 10100 3485 10140 3495
rect 10210 3520 10250 3525
rect 10210 3490 10215 3520
rect 10245 3490 10250 3520
rect 9990 3435 10000 3455
rect 10020 3435 10030 3455
rect 9990 3405 10030 3435
rect 9990 3385 10000 3405
rect 10020 3385 10030 3405
rect 9990 3355 10030 3385
rect 9990 3335 10000 3355
rect 10020 3335 10030 3355
rect 9990 3305 10030 3335
rect 9990 3285 10000 3305
rect 10020 3285 10030 3305
rect 9990 3275 10030 3285
rect 10100 3455 10140 3465
rect 10100 3435 10110 3455
rect 10130 3435 10140 3455
rect 10100 3405 10140 3435
rect 10100 3385 10110 3405
rect 10130 3385 10140 3405
rect 10100 3355 10140 3385
rect 10100 3335 10110 3355
rect 10130 3335 10140 3355
rect 10100 3305 10140 3335
rect 10100 3285 10110 3305
rect 10130 3285 10140 3305
rect 9880 3165 9885 3195
rect 9915 3165 9920 3195
rect 9880 3160 9920 3165
rect 10100 3195 10140 3285
rect 10210 3455 10250 3490
rect 10430 3520 10470 3835
rect 10540 4005 10580 4085
rect 10700 4115 10740 4120
rect 10700 4085 10705 4115
rect 10735 4085 10740 4115
rect 10700 4015 10740 4085
rect 10860 4115 10900 4120
rect 10860 4085 10865 4115
rect 10895 4085 10900 4115
rect 10540 3985 10550 4005
rect 10570 3985 10580 4005
rect 10540 3955 10580 3985
rect 10540 3935 10550 3955
rect 10570 3935 10580 3955
rect 10540 3905 10580 3935
rect 10540 3885 10550 3905
rect 10570 3885 10580 3905
rect 10540 3855 10580 3885
rect 10540 3835 10550 3855
rect 10570 3835 10580 3855
rect 10540 3825 10580 3835
rect 10650 4005 10790 4015
rect 10650 3985 10660 4005
rect 10680 3985 10710 4005
rect 10730 3985 10760 4005
rect 10780 3985 10790 4005
rect 10650 3955 10790 3985
rect 10650 3935 10660 3955
rect 10680 3935 10710 3955
rect 10730 3935 10760 3955
rect 10780 3935 10790 3955
rect 10650 3905 10790 3935
rect 10650 3885 10660 3905
rect 10680 3885 10710 3905
rect 10730 3885 10760 3905
rect 10780 3885 10790 3905
rect 10650 3855 10790 3885
rect 10650 3835 10660 3855
rect 10680 3835 10710 3855
rect 10730 3835 10760 3855
rect 10780 3835 10790 3855
rect 10650 3825 10790 3835
rect 10860 4005 10900 4085
rect 11080 4115 11120 4120
rect 11080 4085 11085 4115
rect 11115 4085 11120 4115
rect 10860 3985 10870 4005
rect 10890 3985 10900 4005
rect 10860 3955 10900 3985
rect 10860 3935 10870 3955
rect 10890 3935 10900 3955
rect 10860 3905 10900 3935
rect 10860 3885 10870 3905
rect 10890 3885 10900 3905
rect 10860 3855 10900 3885
rect 10860 3835 10870 3855
rect 10890 3835 10900 3855
rect 10860 3825 10900 3835
rect 10970 4005 11010 4015
rect 10970 3985 10980 4005
rect 11000 3985 11010 4005
rect 10970 3955 11010 3985
rect 10970 3935 10980 3955
rect 11000 3935 11010 3955
rect 10970 3905 11010 3935
rect 10970 3885 10980 3905
rect 11000 3885 11010 3905
rect 10970 3855 11010 3885
rect 10970 3835 10980 3855
rect 11000 3835 11010 3855
rect 10905 3785 10945 3790
rect 10905 3755 10910 3785
rect 10940 3755 10945 3785
rect 10905 3750 10945 3755
rect 10970 3660 11010 3835
rect 11080 4005 11120 4085
rect 11080 3985 11090 4005
rect 11110 3985 11120 4005
rect 11080 3955 11120 3985
rect 11080 3935 11090 3955
rect 11110 3935 11120 3955
rect 11080 3905 11120 3935
rect 11080 3885 11090 3905
rect 11110 3885 11120 3905
rect 11080 3855 11120 3885
rect 11080 3835 11090 3855
rect 11110 3835 11120 3855
rect 11080 3825 11120 3835
rect 11190 4115 11230 4120
rect 11190 4085 11195 4115
rect 11225 4085 11230 4115
rect 11190 4065 11230 4085
rect 11190 4045 11200 4065
rect 11220 4045 11230 4065
rect 11190 4005 11230 4045
rect 11190 3985 11200 4005
rect 11220 3985 11230 4005
rect 11190 3955 11230 3985
rect 11190 3935 11200 3955
rect 11220 3935 11230 3955
rect 11190 3905 11230 3935
rect 11190 3885 11200 3905
rect 11220 3885 11230 3905
rect 11190 3855 11230 3885
rect 11190 3835 11200 3855
rect 11220 3835 11230 3855
rect 11190 3825 11230 3835
rect 11370 3795 11425 3805
rect 11035 3785 11075 3790
rect 11035 3755 11040 3785
rect 11070 3755 11075 3785
rect 11035 3750 11075 3755
rect 11370 3760 11380 3795
rect 11415 3760 11425 3795
rect 11370 3750 11425 3760
rect 10430 3490 10435 3520
rect 10465 3490 10470 3520
rect 10685 3635 10725 3640
rect 10685 3605 10690 3635
rect 10720 3605 10725 3635
rect 10685 3535 10725 3605
rect 10685 3505 10690 3535
rect 10720 3505 10725 3535
rect 10970 3630 10975 3660
rect 11005 3630 11010 3660
rect 10685 3500 10725 3505
rect 10750 3520 10790 3525
rect 10430 3485 10470 3490
rect 10750 3490 10755 3520
rect 10785 3490 10790 3520
rect 10210 3435 10220 3455
rect 10240 3435 10250 3455
rect 10210 3405 10250 3435
rect 10210 3385 10220 3405
rect 10240 3385 10250 3405
rect 10210 3355 10250 3385
rect 10210 3335 10220 3355
rect 10240 3335 10250 3355
rect 10210 3305 10250 3335
rect 10210 3285 10220 3305
rect 10240 3285 10250 3305
rect 10210 3275 10250 3285
rect 10320 3455 10360 3465
rect 10320 3435 10330 3455
rect 10350 3435 10360 3455
rect 10320 3405 10360 3435
rect 10320 3385 10330 3405
rect 10350 3385 10360 3405
rect 10320 3355 10360 3385
rect 10320 3335 10330 3355
rect 10350 3335 10360 3355
rect 10320 3305 10360 3335
rect 10320 3285 10330 3305
rect 10350 3285 10360 3305
rect 10100 3165 10105 3195
rect 10135 3165 10140 3195
rect 10100 3160 10140 3165
rect 10320 3195 10360 3285
rect 10430 3455 10570 3465
rect 10430 3435 10440 3455
rect 10460 3435 10490 3455
rect 10510 3435 10540 3455
rect 10560 3435 10570 3455
rect 10430 3405 10570 3435
rect 10430 3385 10440 3405
rect 10460 3385 10490 3405
rect 10510 3385 10540 3405
rect 10560 3385 10570 3405
rect 10430 3355 10570 3385
rect 10430 3335 10440 3355
rect 10460 3335 10490 3355
rect 10510 3335 10540 3355
rect 10560 3335 10570 3355
rect 10430 3305 10570 3335
rect 10430 3285 10440 3305
rect 10460 3285 10490 3305
rect 10510 3285 10540 3305
rect 10560 3285 10570 3305
rect 10430 3275 10570 3285
rect 10640 3455 10680 3465
rect 10640 3435 10650 3455
rect 10670 3435 10680 3455
rect 10640 3405 10680 3435
rect 10640 3385 10650 3405
rect 10670 3385 10680 3405
rect 10640 3355 10680 3385
rect 10640 3335 10650 3355
rect 10670 3335 10680 3355
rect 10640 3305 10680 3335
rect 10640 3285 10650 3305
rect 10670 3285 10680 3305
rect 10320 3165 10325 3195
rect 10355 3165 10360 3195
rect 10320 3160 10360 3165
rect 10480 3195 10520 3275
rect 10480 3165 10485 3195
rect 10515 3165 10520 3195
rect 10480 3160 10520 3165
rect 10640 3195 10680 3285
rect 10750 3455 10790 3490
rect 10970 3520 11010 3630
rect 10970 3490 10975 3520
rect 11005 3490 11010 3520
rect 11035 3535 11075 3540
rect 11035 3505 11040 3535
rect 11070 3505 11075 3535
rect 11035 3500 11075 3505
rect 11370 3530 11425 3540
rect 10750 3435 10760 3455
rect 10780 3435 10790 3455
rect 10750 3405 10790 3435
rect 10750 3385 10760 3405
rect 10780 3385 10790 3405
rect 10750 3355 10790 3385
rect 10750 3335 10760 3355
rect 10780 3335 10790 3355
rect 10750 3305 10790 3335
rect 10750 3285 10760 3305
rect 10780 3285 10790 3305
rect 10750 3275 10790 3285
rect 10860 3455 10900 3465
rect 10860 3435 10870 3455
rect 10890 3435 10900 3455
rect 10860 3405 10900 3435
rect 10860 3385 10870 3405
rect 10890 3385 10900 3405
rect 10860 3355 10900 3385
rect 10860 3335 10870 3355
rect 10890 3335 10900 3355
rect 10860 3305 10900 3335
rect 10860 3285 10870 3305
rect 10890 3285 10900 3305
rect 10640 3165 10645 3195
rect 10675 3165 10680 3195
rect 10640 3160 10680 3165
rect 10860 3195 10900 3285
rect 10970 3455 11010 3490
rect 11370 3495 11380 3530
rect 11415 3495 11425 3530
rect 11370 3485 11425 3495
rect 10970 3435 10980 3455
rect 11000 3435 11010 3455
rect 10970 3405 11010 3435
rect 10970 3385 10980 3405
rect 11000 3385 11010 3405
rect 10970 3355 11010 3385
rect 10970 3335 10980 3355
rect 11000 3335 11010 3355
rect 10970 3305 11010 3335
rect 10970 3285 10980 3305
rect 11000 3285 11010 3305
rect 10970 3275 11010 3285
rect 11080 3455 11120 3465
rect 11080 3435 11090 3455
rect 11110 3435 11120 3455
rect 11080 3405 11120 3435
rect 11080 3385 11090 3405
rect 11110 3385 11120 3405
rect 11080 3355 11120 3385
rect 11080 3335 11090 3355
rect 11110 3335 11120 3355
rect 11080 3305 11120 3335
rect 11080 3285 11090 3305
rect 11110 3285 11120 3305
rect 10860 3165 10865 3195
rect 10895 3165 10900 3195
rect 10860 3160 10900 3165
rect 11080 3195 11120 3285
rect 11080 3165 11085 3195
rect 11115 3165 11120 3195
rect 11080 3160 11120 3165
rect 11190 3455 11230 3465
rect 11190 3435 11200 3455
rect 11220 3435 11230 3455
rect 11190 3405 11230 3435
rect 11190 3385 11200 3405
rect 11220 3385 11230 3405
rect 11190 3355 11230 3385
rect 11190 3335 11200 3355
rect 11220 3335 11230 3355
rect 11190 3305 11230 3335
rect 11190 3285 11200 3305
rect 11220 3285 11230 3305
rect 11190 3245 11230 3285
rect 11190 3225 11200 3245
rect 11220 3225 11230 3245
rect 11190 3195 11230 3225
rect 11190 3165 11195 3195
rect 11225 3165 11230 3195
rect 11190 3160 11230 3165
rect 9200 2995 9205 3025
rect 9235 2995 9240 3025
rect 9200 2990 9240 2995
rect 8845 2910 8850 2940
rect 8880 2910 8885 2940
rect 8845 2905 8885 2910
rect 11490 2940 11545 2950
rect 11490 2905 11500 2940
rect 11535 2905 11545 2940
rect 11490 2895 11545 2905
<< via1 >>
rect 9055 4155 9085 4185
rect 6630 4145 6660 4150
rect 6630 4125 6635 4145
rect 6635 4125 6655 4145
rect 6655 4125 6660 4145
rect 6630 4120 6660 4125
rect 6740 4145 6770 4150
rect 6740 4125 6745 4145
rect 6745 4125 6765 4145
rect 6765 4125 6770 4145
rect 6740 4120 6770 4125
rect 6890 4145 6920 4150
rect 6890 4125 6895 4145
rect 6895 4125 6915 4145
rect 6915 4125 6920 4145
rect 6890 4120 6920 4125
rect 7005 4145 7035 4150
rect 7005 4125 7010 4145
rect 7010 4125 7030 4145
rect 7030 4125 7035 4145
rect 7005 4120 7035 4125
rect 7080 4145 7110 4150
rect 7080 4125 7085 4145
rect 7085 4125 7105 4145
rect 7105 4125 7110 4145
rect 7080 4120 7110 4125
rect 7190 4145 7220 4150
rect 7190 4125 7195 4145
rect 7195 4125 7215 4145
rect 7215 4125 7220 4145
rect 7190 4120 7220 4125
rect 7340 4145 7370 4150
rect 7340 4125 7345 4145
rect 7345 4125 7365 4145
rect 7365 4125 7370 4145
rect 7340 4120 7370 4125
rect 7450 4145 7480 4150
rect 7450 4125 7455 4145
rect 7455 4125 7475 4145
rect 7475 4125 7480 4145
rect 7450 4120 7480 4125
rect 7650 4145 7680 4150
rect 7650 4125 7655 4145
rect 7655 4125 7675 4145
rect 7675 4125 7680 4145
rect 7650 4120 7680 4125
rect 7815 4145 7845 4150
rect 7815 4125 7820 4145
rect 7820 4125 7840 4145
rect 7840 4125 7845 4145
rect 7815 4120 7845 4125
rect 7980 4145 8010 4150
rect 7980 4125 7985 4145
rect 7985 4125 8005 4145
rect 8005 4125 8010 4145
rect 7980 4120 8010 4125
rect 8200 4145 8230 4150
rect 8200 4125 8205 4145
rect 8205 4125 8225 4145
rect 8225 4125 8230 4145
rect 8200 4120 8230 4125
rect 8330 4120 8360 4150
rect 8590 4145 8620 4150
rect 8590 4125 8595 4145
rect 8595 4125 8615 4145
rect 8615 4125 8620 4145
rect 8590 4120 8620 4125
rect 8930 4145 8960 4150
rect 8930 4125 8935 4145
rect 8935 4125 8955 4145
rect 8955 4125 8960 4145
rect 8930 4120 8960 4125
rect 6570 3900 6600 3905
rect 6570 3880 6575 3900
rect 6575 3880 6595 3900
rect 6595 3880 6600 3900
rect 6570 3875 6600 3880
rect 7530 3895 7560 3900
rect 7530 3875 7535 3895
rect 7535 3875 7555 3895
rect 7555 3875 7560 3895
rect 7530 3870 7560 3875
rect 8045 3895 8075 3900
rect 8045 3875 8050 3895
rect 8050 3875 8070 3895
rect 8070 3875 8075 3895
rect 8045 3870 8075 3875
rect 6855 3610 6885 3615
rect 6855 3590 6860 3610
rect 6860 3590 6880 3610
rect 6880 3590 6885 3610
rect 6855 3585 6885 3590
rect 6630 3555 6660 3560
rect 6630 3535 6635 3555
rect 6635 3535 6655 3555
rect 6655 3535 6660 3555
rect 6630 3530 6660 3535
rect 7000 3555 7030 3560
rect 7000 3535 7005 3555
rect 7005 3535 7025 3555
rect 7025 3535 7030 3555
rect 7000 3530 7030 3535
rect 7080 3555 7110 3560
rect 7080 3535 7085 3555
rect 7085 3535 7105 3555
rect 7105 3535 7110 3555
rect 7080 3530 7110 3535
rect 7450 3555 7480 3560
rect 7450 3535 7455 3555
rect 7455 3535 7475 3555
rect 7475 3535 7480 3555
rect 7450 3530 7480 3535
rect 6570 3210 6600 3215
rect 6570 3190 6575 3210
rect 6575 3190 6595 3210
rect 6595 3190 6600 3210
rect 6570 3185 6600 3190
rect 7620 3585 7650 3615
rect 7575 3555 7605 3560
rect 7575 3535 7580 3555
rect 7580 3535 7600 3555
rect 7600 3535 7605 3555
rect 7575 3530 7605 3535
rect 7670 3555 7700 3560
rect 7670 3535 7675 3555
rect 7675 3535 7695 3555
rect 7695 3535 7700 3555
rect 7670 3530 7700 3535
rect 7710 3555 7740 3560
rect 7710 3535 7715 3555
rect 7715 3535 7735 3555
rect 7735 3535 7740 3555
rect 7710 3530 7740 3535
rect 7815 3555 7845 3560
rect 7815 3535 7820 3555
rect 7820 3535 7840 3555
rect 7840 3535 7845 3555
rect 7815 3530 7845 3535
rect 7980 3555 8010 3560
rect 7980 3535 7985 3555
rect 7985 3535 8005 3555
rect 8005 3535 8010 3555
rect 7980 3530 8010 3535
rect 7630 3500 7660 3505
rect 7630 3480 7635 3500
rect 7635 3480 7655 3500
rect 7655 3480 7660 3500
rect 7630 3475 7660 3480
rect 8120 3590 8150 3620
rect 8455 4090 8485 4095
rect 8455 4070 8460 4090
rect 8460 4070 8480 4090
rect 8480 4070 8485 4090
rect 8455 4065 8485 4070
rect 8770 4090 8800 4095
rect 8770 4070 8775 4090
rect 8775 4070 8795 4090
rect 8795 4070 8800 4090
rect 8770 4065 8800 4070
rect 11555 4155 11590 4190
rect 9055 4065 9085 4095
rect 9675 4085 9705 4115
rect 8330 3585 8360 3615
rect 8415 3610 8445 3615
rect 8415 3590 8420 3610
rect 8420 3590 8440 3610
rect 8440 3590 8445 3610
rect 8415 3585 8445 3590
rect 9005 3920 9035 3925
rect 9005 3900 9010 3920
rect 9010 3900 9030 3920
rect 9030 3900 9035 3920
rect 9005 3895 9035 3900
rect 9095 3895 9125 3925
rect 9785 4085 9815 4115
rect 10005 4085 10035 4115
rect 10165 4085 10195 4115
rect 10325 4085 10355 4115
rect 10545 4085 10575 4115
rect 9095 3715 9125 3745
rect 9095 3660 9125 3690
rect 8735 3610 8765 3615
rect 8735 3590 8740 3610
rect 8740 3590 8760 3610
rect 8760 3590 8765 3610
rect 8735 3585 8765 3590
rect 9895 3660 9925 3690
rect 9095 3585 9125 3615
rect 9150 3605 9180 3635
rect 8200 3555 8230 3560
rect 8200 3535 8205 3555
rect 8205 3535 8225 3555
rect 8225 3535 8230 3555
rect 8200 3530 8230 3535
rect 8395 3555 8425 3560
rect 8395 3535 8400 3555
rect 8400 3535 8420 3555
rect 8420 3535 8425 3555
rect 8395 3530 8425 3535
rect 8500 3530 8530 3560
rect 8590 3555 8620 3560
rect 8590 3535 8595 3555
rect 8595 3535 8615 3555
rect 8615 3535 8620 3555
rect 8590 3530 8620 3535
rect 8930 3555 8960 3560
rect 8930 3535 8935 3555
rect 8935 3535 8955 3555
rect 8955 3535 8960 3555
rect 8930 3530 8960 3535
rect 7520 3195 7550 3200
rect 7520 3175 7525 3195
rect 7525 3175 7545 3195
rect 7545 3175 7550 3195
rect 7520 3170 7550 3175
rect 8065 3215 8095 3220
rect 8065 3195 8070 3215
rect 8070 3195 8090 3215
rect 8090 3195 8095 3215
rect 8065 3190 8095 3195
rect 8850 3230 8880 3235
rect 8850 3210 8855 3230
rect 8855 3210 8875 3230
rect 8875 3210 8880 3230
rect 8850 3205 8880 3210
rect 6835 3020 6865 3025
rect 6835 3000 6840 3020
rect 6840 3000 6860 3020
rect 6860 3000 6865 3020
rect 6835 2995 6865 3000
rect 7695 3020 7725 3025
rect 7695 3000 7700 3020
rect 7700 3000 7720 3020
rect 7720 3000 7725 3020
rect 7695 2995 7725 3000
rect 8120 3005 8150 3035
rect 8735 3020 8765 3025
rect 8735 3000 8740 3020
rect 8740 3000 8760 3020
rect 8760 3000 8765 3020
rect 8735 2995 8765 3000
rect 6630 2965 6660 2970
rect 6630 2945 6635 2965
rect 6635 2945 6655 2965
rect 6655 2945 6660 2965
rect 6630 2940 6660 2945
rect 6740 2965 6770 2970
rect 6740 2945 6745 2965
rect 6745 2945 6765 2965
rect 6765 2945 6770 2965
rect 6740 2940 6770 2945
rect 6890 2965 6920 2970
rect 6890 2945 6895 2965
rect 6895 2945 6915 2965
rect 6915 2945 6920 2965
rect 6890 2940 6920 2945
rect 7000 2965 7030 2970
rect 7000 2945 7005 2965
rect 7005 2945 7025 2965
rect 7025 2945 7030 2965
rect 7000 2940 7030 2945
rect 7080 2965 7110 2970
rect 7080 2945 7085 2965
rect 7085 2945 7105 2965
rect 7105 2945 7110 2965
rect 7080 2940 7110 2945
rect 7190 2965 7220 2970
rect 7190 2945 7195 2965
rect 7195 2945 7215 2965
rect 7215 2945 7220 2965
rect 7190 2940 7220 2945
rect 7340 2965 7370 2970
rect 7340 2945 7345 2965
rect 7345 2945 7365 2965
rect 7365 2945 7370 2965
rect 7340 2940 7370 2945
rect 7450 2965 7480 2970
rect 7450 2945 7455 2965
rect 7455 2945 7475 2965
rect 7475 2945 7480 2965
rect 7450 2940 7480 2945
rect 7600 2965 7630 2970
rect 7600 2945 7605 2965
rect 7605 2945 7625 2965
rect 7625 2945 7630 2965
rect 7600 2940 7630 2945
rect 7820 2965 7850 2970
rect 7820 2945 7825 2965
rect 7825 2945 7845 2965
rect 7845 2945 7850 2965
rect 7820 2940 7850 2945
rect 7985 2965 8015 2970
rect 7985 2945 7990 2965
rect 7990 2945 8010 2965
rect 8010 2945 8015 2965
rect 7985 2940 8015 2945
rect 8200 2965 8230 2970
rect 8200 2945 8205 2965
rect 8205 2945 8225 2965
rect 8225 2945 8230 2965
rect 8200 2940 8230 2945
rect 8395 2965 8425 2970
rect 8395 2945 8400 2965
rect 8400 2945 8420 2965
rect 8420 2945 8425 2965
rect 8395 2940 8425 2945
rect 8590 2965 8620 2970
rect 8590 2945 8595 2965
rect 8595 2945 8615 2965
rect 8615 2945 8620 2965
rect 8590 2940 8620 2945
rect 9005 3190 9035 3195
rect 9005 3170 9010 3190
rect 9010 3170 9030 3190
rect 9030 3170 9035 3190
rect 9005 3165 9035 3170
rect 9150 3165 9180 3195
rect 9205 3550 9235 3580
rect 10105 3550 10135 3580
rect 9995 3490 10025 3520
rect 9775 3165 9805 3195
rect 10215 3490 10245 3520
rect 9885 3165 9915 3195
rect 10705 4085 10735 4115
rect 10865 4085 10895 4115
rect 11085 4085 11115 4115
rect 10910 3780 10940 3785
rect 10910 3760 10915 3780
rect 10915 3760 10935 3780
rect 10935 3760 10940 3780
rect 10910 3755 10940 3760
rect 11195 4085 11225 4115
rect 11040 3780 11070 3785
rect 11040 3760 11045 3780
rect 11045 3760 11065 3780
rect 11065 3760 11070 3780
rect 11040 3755 11070 3760
rect 11380 3760 11415 3795
rect 10435 3490 10465 3520
rect 10690 3605 10720 3635
rect 10690 3530 10720 3535
rect 10690 3510 10695 3530
rect 10695 3510 10715 3530
rect 10715 3510 10720 3530
rect 10690 3505 10720 3510
rect 10975 3630 11005 3660
rect 10755 3490 10785 3520
rect 10105 3165 10135 3195
rect 10325 3165 10355 3195
rect 10485 3165 10515 3195
rect 10975 3490 11005 3520
rect 11040 3530 11070 3535
rect 11040 3510 11045 3530
rect 11045 3510 11065 3530
rect 11065 3510 11070 3530
rect 11040 3505 11070 3510
rect 10645 3165 10675 3195
rect 11380 3495 11415 3530
rect 10865 3165 10895 3195
rect 11085 3165 11115 3195
rect 11195 3165 11225 3195
rect 9205 2995 9235 3025
rect 8850 2910 8880 2940
rect 11500 2905 11535 2940
<< metal2 >>
rect 11545 4190 11600 4200
rect 9050 4185 11555 4190
rect 9050 4155 9055 4185
rect 9085 4155 11555 4185
rect 11590 4155 11600 4190
rect 6505 4150 8965 4155
rect 9050 4150 11600 4155
rect 6505 4120 6630 4150
rect 6660 4120 6740 4150
rect 6770 4120 6890 4150
rect 6920 4120 7005 4150
rect 7035 4120 7080 4150
rect 7110 4120 7190 4150
rect 7220 4120 7340 4150
rect 7370 4120 7450 4150
rect 7480 4120 7650 4150
rect 7680 4120 7815 4150
rect 7845 4120 7980 4150
rect 8010 4120 8200 4150
rect 8230 4120 8330 4150
rect 8360 4120 8590 4150
rect 8620 4120 8930 4150
rect 8960 4120 8965 4150
rect 11545 4145 11600 4150
rect 6505 4115 8965 4120
rect 9670 4115 11230 4120
rect 8450 4095 8490 4100
rect 8450 4065 8455 4095
rect 8485 4065 8490 4095
rect 8450 4060 8490 4065
rect 8765 4095 9090 4100
rect 8765 4065 8770 4095
rect 8800 4065 9055 4095
rect 9085 4065 9090 4095
rect 9670 4085 9675 4115
rect 9705 4085 9785 4115
rect 9815 4085 10005 4115
rect 10035 4085 10165 4115
rect 10195 4085 10325 4115
rect 10355 4085 10545 4115
rect 10575 4085 10705 4115
rect 10735 4085 10865 4115
rect 10895 4085 11085 4115
rect 11115 4085 11195 4115
rect 11225 4085 11230 4115
rect 9670 4080 11230 4085
rect 8765 4060 9090 4065
rect 9000 3925 9130 3930
rect 6505 3905 6605 3910
rect 6505 3875 6570 3905
rect 6600 3875 6605 3905
rect 6505 3870 6605 3875
rect 7525 3900 7565 3905
rect 7525 3870 7530 3900
rect 7560 3870 7565 3900
rect 7525 3865 7565 3870
rect 8040 3900 8080 3905
rect 8040 3870 8045 3900
rect 8075 3870 8080 3900
rect 9000 3895 9005 3925
rect 9035 3895 9095 3925
rect 9125 3895 9130 3925
rect 9000 3890 9130 3895
rect 8040 3865 8080 3870
rect 11370 3795 11425 3805
rect 11370 3790 11380 3795
rect 10905 3785 10945 3790
rect 10905 3755 10910 3785
rect 10940 3755 10945 3785
rect 10905 3750 10945 3755
rect 11035 3785 11380 3790
rect 11035 3755 11040 3785
rect 11070 3760 11380 3785
rect 11415 3760 11425 3795
rect 11070 3755 11425 3760
rect 11035 3750 11425 3755
rect 9090 3745 10945 3750
rect 9090 3715 9095 3745
rect 9125 3715 10945 3745
rect 9090 3710 10945 3715
rect 9090 3690 9930 3695
rect 9090 3660 9095 3690
rect 9125 3660 9895 3690
rect 9925 3660 9930 3690
rect 9090 3655 9930 3660
rect 10970 3660 12095 3665
rect 9145 3635 10725 3640
rect 8115 3620 8155 3625
rect 6850 3615 6890 3620
rect 6850 3585 6855 3615
rect 6885 3610 6890 3615
rect 7615 3615 7655 3620
rect 8115 3615 8120 3620
rect 7615 3610 7620 3615
rect 6885 3590 7620 3610
rect 6885 3585 6890 3590
rect 6850 3580 6890 3585
rect 7615 3585 7620 3590
rect 7650 3595 8120 3615
rect 7650 3585 7655 3595
rect 8115 3590 8120 3595
rect 8150 3590 8155 3620
rect 8410 3615 8450 3620
rect 8115 3585 8155 3590
rect 8325 3585 8330 3615
rect 8360 3610 8365 3615
rect 8410 3610 8415 3615
rect 8360 3590 8415 3610
rect 8360 3585 8365 3590
rect 8410 3585 8415 3590
rect 8445 3585 8450 3615
rect 8730 3615 9130 3620
rect 8730 3585 8735 3615
rect 8765 3585 9095 3615
rect 9125 3585 9130 3615
rect 9145 3605 9150 3635
rect 9180 3605 10690 3635
rect 10720 3605 10725 3635
rect 10970 3630 10975 3660
rect 11005 3630 12095 3660
rect 10970 3625 12095 3630
rect 9145 3600 10725 3605
rect 7615 3580 7655 3585
rect 8730 3580 9130 3585
rect 9200 3580 10140 3585
rect 6505 3560 8965 3565
rect 6505 3530 6630 3560
rect 6660 3530 7000 3560
rect 7030 3530 7080 3560
rect 7110 3530 7450 3560
rect 7480 3530 7575 3560
rect 7605 3530 7670 3560
rect 7700 3530 7710 3560
rect 7740 3530 7815 3560
rect 7845 3530 7980 3560
rect 8010 3530 8200 3560
rect 8230 3530 8395 3560
rect 8425 3530 8500 3560
rect 8530 3530 8590 3560
rect 8620 3530 8930 3560
rect 8960 3530 8965 3560
rect 9200 3550 9205 3580
rect 9235 3550 10105 3580
rect 10135 3550 10140 3580
rect 9200 3545 10140 3550
rect 6505 3525 8965 3530
rect 10685 3535 10725 3540
rect 9990 3520 10470 3525
rect 7625 3475 7630 3505
rect 7660 3475 7665 3505
rect 9990 3490 9995 3520
rect 10025 3490 10215 3520
rect 10245 3490 10435 3520
rect 10465 3490 10470 3520
rect 10685 3505 10690 3535
rect 10720 3505 10725 3535
rect 11035 3535 11425 3540
rect 10685 3500 10725 3505
rect 10750 3520 11010 3525
rect 9990 3485 10470 3490
rect 10750 3490 10755 3520
rect 10785 3490 10975 3520
rect 11005 3490 11010 3520
rect 11035 3505 11040 3535
rect 11070 3530 11425 3535
rect 11070 3505 11380 3530
rect 11035 3500 11380 3505
rect 10750 3485 11010 3490
rect 11370 3495 11380 3500
rect 11415 3495 11425 3530
rect 11370 3485 11425 3495
rect 7625 3470 7665 3475
rect 8845 3235 8885 3240
rect 8060 3220 8100 3225
rect 6505 3215 6605 3220
rect 6505 3185 6570 3215
rect 6600 3185 6605 3215
rect 6505 3180 6605 3185
rect 7515 3200 7555 3205
rect 7515 3170 7520 3200
rect 7550 3170 7555 3200
rect 8060 3190 8065 3220
rect 8095 3190 8100 3220
rect 8845 3205 8850 3235
rect 8880 3205 8885 3235
rect 8845 3200 8885 3205
rect 8060 3185 8100 3190
rect 9000 3195 9185 3200
rect 7515 3165 7555 3170
rect 9000 3165 9005 3195
rect 9035 3165 9150 3195
rect 9180 3165 9185 3195
rect 9000 3160 9185 3165
rect 9770 3195 11230 3200
rect 9770 3165 9775 3195
rect 9805 3165 9885 3195
rect 9915 3165 10105 3195
rect 10135 3165 10325 3195
rect 10355 3165 10485 3195
rect 10515 3165 10645 3195
rect 10675 3165 10865 3195
rect 10895 3165 11085 3195
rect 11115 3165 11195 3195
rect 11225 3165 11230 3195
rect 9770 3160 11230 3165
rect 8115 3035 8155 3040
rect 8115 3030 8120 3035
rect 6830 3025 8120 3030
rect 6830 2995 6835 3025
rect 6865 3010 7695 3025
rect 6865 2995 6870 3010
rect 6830 2990 6870 2995
rect 7690 2995 7695 3010
rect 7725 3010 8120 3025
rect 7725 2995 7730 3010
rect 8115 3005 8120 3010
rect 8150 3005 8155 3035
rect 8115 3000 8155 3005
rect 8730 3025 9240 3030
rect 7690 2990 7730 2995
rect 8730 2995 8735 3025
rect 8765 2995 9205 3025
rect 9235 2995 9240 3025
rect 8730 2990 9240 2995
rect 6505 2970 8625 2975
rect 6505 2940 6630 2970
rect 6660 2940 6740 2970
rect 6770 2940 6890 2970
rect 6920 2940 7000 2970
rect 7030 2940 7080 2970
rect 7110 2940 7190 2970
rect 7220 2940 7340 2970
rect 7370 2940 7450 2970
rect 7480 2940 7600 2970
rect 7630 2940 7820 2970
rect 7850 2940 7985 2970
rect 8015 2940 8200 2970
rect 8230 2940 8395 2970
rect 8425 2940 8590 2970
rect 8620 2940 8625 2970
rect 11490 2945 11545 2950
rect 6505 2935 8625 2940
rect 8845 2940 11545 2945
rect 8845 2910 8850 2940
rect 8880 2910 11500 2940
rect 8845 2905 11500 2910
rect 11535 2905 11545 2940
rect 11490 2895 11545 2905
<< via2 >>
rect 11555 4155 11590 4190
rect 11380 3760 11415 3795
rect 11380 3495 11415 3530
rect 11500 2905 11535 2940
<< metal3 >>
rect 11545 4190 11600 4200
rect 11545 4155 11555 4190
rect 11590 4155 11600 4190
rect 11545 4145 11600 4155
rect 11370 3795 11425 3805
rect 11370 3760 11380 3795
rect 11415 3760 11425 3795
rect 11370 3750 11425 3760
rect 11545 3735 11845 4145
rect 11370 3530 11425 3540
rect 11370 3495 11380 3530
rect 11415 3495 11425 3530
rect 11370 3485 11425 3495
rect 11545 2950 12095 3555
rect 11490 2940 12095 2950
rect 11490 2905 11500 2940
rect 11535 2905 12095 2940
rect 11490 2895 12095 2905
<< via3 >>
rect 11380 3760 11415 3795
rect 11380 3495 11415 3530
<< mimcap >>
rect 11560 3795 11830 4130
rect 11560 3760 11570 3795
rect 11605 3760 11830 3795
rect 11560 3750 11830 3760
rect 11560 3530 12080 3540
rect 11560 3495 11570 3530
rect 11605 3495 12080 3530
rect 11560 2910 12080 3495
<< mimcapcontact >>
rect 11570 3760 11605 3795
rect 11570 3495 11605 3530
<< metal4 >>
rect 11370 3795 11615 3805
rect 11370 3760 11380 3795
rect 11415 3760 11570 3795
rect 11605 3760 11615 3795
rect 11370 3750 11615 3760
rect 11370 3530 11615 3540
rect 11370 3495 11380 3530
rect 11415 3495 11570 3530
rect 11605 3495 11615 3530
rect 11370 3485 11615 3495
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
