MACRO divide_by_120
  CLASS BLOCK ;
  FOREIGN divide_by_120 ;
  ORIGIN -210.650 -14.450 ;
  SIZE 53.400 BY 4.300 ;
  OBS
      LAYER nwell ;
        RECT 211.300 16.950 263.850 18.000 ;
      LAYER li1 ;
        RECT 213.300 18.350 213.700 18.750 ;
        RECT 215.400 18.350 215.800 18.750 ;
        RECT 218.750 18.350 219.150 18.750 ;
        RECT 221.600 18.350 222.000 18.750 ;
        RECT 225.350 18.350 225.750 18.750 ;
        RECT 227.500 18.350 227.900 18.750 ;
        RECT 229.700 18.350 230.100 18.750 ;
        RECT 230.950 18.350 231.350 18.750 ;
        RECT 232.050 18.350 232.450 18.750 ;
        RECT 234.400 18.350 234.800 18.750 ;
        RECT 236.600 18.350 237.000 18.750 ;
        RECT 239.700 18.350 240.100 18.750 ;
        RECT 241.400 18.350 241.800 18.750 ;
        RECT 243.200 18.350 243.600 18.750 ;
        RECT 246.200 18.350 246.600 18.750 ;
        RECT 247.900 18.350 248.300 18.750 ;
        RECT 249.700 18.350 250.100 18.750 ;
        RECT 252.700 18.350 253.100 18.750 ;
        RECT 254.400 18.350 254.800 18.750 ;
        RECT 256.200 18.350 256.600 18.750 ;
        RECT 259.200 18.350 259.600 18.750 ;
        RECT 260.900 18.350 261.300 18.750 ;
        RECT 262.700 18.350 263.100 18.750 ;
        RECT 213.400 17.600 213.600 18.350 ;
        RECT 214.900 17.800 215.300 18.200 ;
        RECT 215.500 17.600 215.700 18.350 ;
        RECT 215.900 17.800 216.250 18.200 ;
        RECT 216.050 17.600 216.250 17.800 ;
        RECT 216.450 17.700 216.850 18.100 ;
        RECT 218.850 17.600 219.050 18.350 ;
        RECT 220.500 17.800 220.900 18.200 ;
        RECT 221.200 17.800 221.500 18.200 ;
        RECT 221.700 17.600 221.900 18.350 ;
        RECT 225.450 17.600 225.650 18.350 ;
        RECT 227.000 17.800 227.400 18.200 ;
        RECT 227.600 17.600 227.800 18.350 ;
        RECT 228.100 17.800 228.500 18.200 ;
        RECT 228.100 17.600 228.300 17.800 ;
        RECT 229.800 17.600 230.000 18.350 ;
        RECT 231.050 17.600 231.250 18.350 ;
        RECT 232.150 17.600 232.350 18.350 ;
        RECT 233.750 17.850 234.150 18.200 ;
        RECT 233.950 17.600 234.150 17.850 ;
        RECT 234.500 17.600 234.700 18.350 ;
        RECT 235.800 17.850 236.200 18.200 ;
        RECT 236.700 17.600 236.900 18.350 ;
        RECT 239.800 17.600 240.000 18.350 ;
        RECT 241.500 17.600 241.700 18.350 ;
        RECT 243.300 17.600 243.500 18.350 ;
        RECT 245.550 17.800 245.950 18.200 ;
        RECT 245.750 17.600 245.950 17.800 ;
        RECT 246.300 17.600 246.500 18.350 ;
        RECT 248.000 17.600 248.200 18.350 ;
        RECT 248.450 17.800 248.850 18.200 ;
        RECT 249.800 17.600 250.000 18.350 ;
        RECT 252.050 17.800 252.450 18.200 ;
        RECT 252.250 17.600 252.450 17.800 ;
        RECT 252.800 17.600 253.000 18.350 ;
        RECT 254.500 17.600 254.700 18.350 ;
        RECT 254.950 17.800 255.350 18.200 ;
        RECT 256.300 17.600 256.500 18.350 ;
        RECT 258.550 17.800 258.950 18.200 ;
        RECT 258.750 17.600 258.950 17.800 ;
        RECT 259.300 17.600 259.500 18.350 ;
        RECT 261.000 17.600 261.200 18.350 ;
        RECT 261.450 17.800 261.850 18.200 ;
        RECT 262.800 17.600 263.000 18.350 ;
        RECT 211.500 17.500 211.900 17.600 ;
        RECT 212.800 17.500 213.100 17.600 ;
        RECT 211.500 17.300 213.100 17.500 ;
        RECT 211.500 17.200 211.900 17.300 ;
        RECT 212.800 17.200 213.100 17.300 ;
        RECT 213.350 17.200 214.050 17.600 ;
        RECT 214.900 17.500 215.200 17.600 ;
        RECT 214.250 17.300 215.200 17.500 ;
        RECT 211.600 16.750 211.800 17.200 ;
        RECT 211.200 16.350 211.800 16.750 ;
        RECT 211.600 16.000 211.800 16.350 ;
        RECT 212.250 16.400 212.650 16.600 ;
        RECT 214.250 16.400 214.450 17.300 ;
        RECT 214.900 17.200 215.200 17.300 ;
        RECT 215.450 17.200 215.750 17.600 ;
        RECT 216.000 17.200 216.300 17.600 ;
        RECT 218.250 17.500 218.550 17.600 ;
        RECT 217.150 17.300 218.550 17.500 ;
        RECT 216.050 17.000 216.250 17.200 ;
        RECT 212.250 16.200 214.450 16.400 ;
        RECT 213.150 16.000 213.350 16.200 ;
        RECT 214.250 16.000 214.450 16.200 ;
        RECT 214.700 16.800 216.250 17.000 ;
        RECT 214.700 16.000 214.900 16.800 ;
        RECT 217.150 16.600 217.350 17.300 ;
        RECT 218.250 17.200 218.550 17.300 ;
        RECT 218.800 17.200 219.100 17.600 ;
        RECT 219.350 17.200 219.650 17.600 ;
        RECT 220.450 17.200 220.750 17.600 ;
        RECT 221.000 17.200 221.300 17.600 ;
        RECT 221.550 17.200 221.900 17.600 ;
        RECT 222.100 17.200 222.400 17.600 ;
        RECT 223.650 17.500 224.050 17.600 ;
        RECT 224.850 17.500 225.150 17.600 ;
        RECT 223.650 17.300 225.150 17.500 ;
        RECT 223.650 17.200 224.050 17.300 ;
        RECT 224.850 17.200 225.150 17.300 ;
        RECT 225.400 17.200 226.100 17.600 ;
        RECT 226.950 17.500 227.250 17.600 ;
        RECT 226.300 17.300 227.250 17.500 ;
        RECT 217.850 16.600 218.250 17.000 ;
        RECT 215.150 16.500 215.550 16.600 ;
        RECT 216.850 16.500 217.350 16.600 ;
        RECT 215.150 16.300 217.350 16.500 ;
        RECT 215.150 16.200 215.550 16.300 ;
        RECT 216.850 16.200 217.350 16.300 ;
        RECT 218.050 16.400 218.250 16.600 ;
        RECT 219.350 16.400 219.550 17.200 ;
        RECT 219.850 17.000 220.250 17.200 ;
        RECT 220.500 17.000 220.700 17.200 ;
        RECT 222.150 17.000 222.350 17.200 ;
        RECT 219.850 16.800 223.150 17.000 ;
        RECT 218.050 16.200 219.550 16.400 ;
        RECT 219.750 16.200 220.150 16.550 ;
        RECT 220.500 16.200 221.800 16.400 ;
        RECT 222.350 16.200 222.750 16.550 ;
        RECT 217.150 16.000 217.350 16.200 ;
        RECT 218.250 16.000 218.450 16.200 ;
        RECT 219.350 16.000 219.550 16.200 ;
        RECT 220.500 16.000 220.700 16.200 ;
        RECT 221.600 16.000 221.800 16.200 ;
        RECT 222.950 16.000 223.150 16.800 ;
        RECT 211.600 15.600 212.300 16.000 ;
        RECT 212.550 15.600 212.850 16.000 ;
        RECT 213.100 15.600 213.400 16.000 ;
        RECT 213.650 15.600 213.950 16.000 ;
        RECT 214.200 15.600 214.500 16.000 ;
        RECT 214.700 15.700 215.200 16.000 ;
        RECT 214.900 15.600 215.200 15.700 ;
        RECT 215.450 15.600 215.750 16.000 ;
        RECT 216.000 15.600 216.300 16.000 ;
        RECT 217.150 15.600 217.450 16.000 ;
        RECT 217.700 15.600 218.000 16.000 ;
        RECT 218.250 15.600 218.550 16.000 ;
        RECT 218.800 15.600 219.100 16.000 ;
        RECT 219.350 15.600 219.650 16.000 ;
        RECT 220.450 15.600 220.750 16.000 ;
        RECT 221.000 15.600 221.300 16.000 ;
        RECT 221.550 15.600 221.850 16.000 ;
        RECT 222.100 15.600 222.400 16.000 ;
        RECT 222.650 15.700 223.150 16.000 ;
        RECT 223.850 16.000 224.050 17.200 ;
        RECT 224.300 16.400 224.700 16.550 ;
        RECT 226.300 16.400 226.500 17.300 ;
        RECT 226.950 17.200 227.250 17.300 ;
        RECT 227.500 17.200 227.800 17.600 ;
        RECT 228.050 17.200 228.350 17.600 ;
        RECT 229.200 17.200 229.500 17.600 ;
        RECT 229.750 17.200 230.050 17.600 ;
        RECT 230.300 17.200 230.600 17.600 ;
        RECT 231.000 17.200 231.300 17.600 ;
        RECT 231.550 17.200 231.850 17.600 ;
        RECT 232.100 17.200 232.400 17.600 ;
        RECT 233.900 17.500 234.200 17.600 ;
        RECT 232.800 17.300 234.200 17.500 ;
        RECT 228.100 17.000 228.300 17.200 ;
        RECT 224.300 16.200 226.500 16.400 ;
        RECT 225.200 16.000 225.400 16.200 ;
        RECT 226.300 16.000 226.500 16.200 ;
        RECT 226.750 16.800 228.300 17.000 ;
        RECT 228.550 17.000 228.950 17.200 ;
        RECT 229.250 17.000 229.450 17.200 ;
        RECT 230.350 17.000 230.550 17.200 ;
        RECT 228.550 16.800 230.550 17.000 ;
        RECT 226.750 16.000 226.950 16.800 ;
        RECT 227.200 16.500 227.600 16.600 ;
        RECT 228.250 16.500 228.650 16.550 ;
        RECT 227.200 16.300 228.650 16.500 ;
        RECT 227.200 16.200 227.600 16.300 ;
        RECT 228.250 16.200 228.650 16.300 ;
        RECT 223.850 15.700 224.350 16.000 ;
        RECT 222.650 15.600 222.950 15.700 ;
        RECT 224.050 15.600 224.350 15.700 ;
        RECT 224.600 15.600 224.900 16.000 ;
        RECT 225.150 15.600 225.450 16.000 ;
        RECT 225.700 15.600 226.000 16.000 ;
        RECT 226.250 15.600 226.550 16.000 ;
        RECT 226.750 15.700 227.250 16.000 ;
        RECT 226.950 15.600 227.250 15.700 ;
        RECT 227.500 15.600 227.800 16.000 ;
        RECT 228.050 15.600 228.750 16.000 ;
        RECT 228.950 15.900 229.150 16.800 ;
        RECT 231.600 16.650 231.800 17.200 ;
        RECT 232.800 16.850 233.000 17.300 ;
        RECT 233.900 17.200 234.200 17.300 ;
        RECT 234.450 17.200 234.750 17.600 ;
        RECT 235.000 17.200 235.300 17.600 ;
        RECT 236.100 17.200 236.400 17.600 ;
        RECT 236.650 17.200 236.950 17.600 ;
        RECT 237.200 17.500 237.500 17.600 ;
        RECT 238.450 17.500 238.850 17.600 ;
        RECT 239.200 17.500 239.500 17.600 ;
        RECT 237.200 17.300 238.250 17.500 ;
        RECT 237.200 17.200 237.500 17.300 ;
        RECT 231.150 16.600 231.800 16.650 ;
        RECT 229.450 16.400 231.800 16.600 ;
        RECT 232.500 16.450 233.000 16.850 ;
        RECT 233.500 16.600 233.900 17.000 ;
        RECT 229.450 16.200 229.850 16.400 ;
        RECT 231.150 16.250 231.800 16.400 ;
        RECT 231.600 16.000 231.800 16.250 ;
        RECT 232.800 16.000 233.000 16.450 ;
        RECT 233.700 16.400 233.900 16.600 ;
        RECT 235.000 16.400 235.200 17.200 ;
        RECT 235.500 17.000 235.900 17.200 ;
        RECT 236.150 17.000 236.350 17.200 ;
        RECT 237.250 17.000 237.450 17.200 ;
        RECT 235.500 16.800 237.450 17.000 ;
        RECT 233.700 16.200 235.200 16.400 ;
        RECT 235.650 16.500 236.050 16.550 ;
        RECT 237.450 16.500 237.850 16.550 ;
        RECT 235.650 16.300 237.850 16.500 ;
        RECT 235.650 16.200 236.050 16.300 ;
        RECT 237.450 16.200 237.850 16.300 ;
        RECT 233.900 16.000 234.100 16.200 ;
        RECT 235.000 16.000 235.200 16.200 ;
        RECT 238.050 16.000 238.250 17.300 ;
        RECT 238.450 17.300 239.500 17.500 ;
        RECT 238.450 17.200 238.850 17.300 ;
        RECT 239.200 17.200 239.500 17.300 ;
        RECT 239.750 17.200 240.450 17.600 ;
        RECT 240.750 17.200 241.200 17.600 ;
        RECT 241.450 17.200 241.750 17.600 ;
        RECT 242.000 17.200 242.300 17.600 ;
        RECT 242.700 17.200 243.000 17.600 ;
        RECT 243.250 17.200 243.550 17.600 ;
        RECT 243.800 17.200 244.100 17.600 ;
        RECT 245.700 17.500 246.000 17.600 ;
        RECT 245.150 17.300 246.000 17.500 ;
        RECT 229.750 15.900 230.050 16.000 ;
        RECT 228.950 15.700 230.050 15.900 ;
        RECT 229.750 15.600 230.050 15.700 ;
        RECT 230.300 15.600 230.600 16.000 ;
        RECT 231.550 15.600 231.850 16.000 ;
        RECT 232.100 15.600 232.400 16.000 ;
        RECT 232.800 15.600 233.100 16.000 ;
        RECT 233.350 15.600 233.650 16.000 ;
        RECT 233.900 15.600 234.200 16.000 ;
        RECT 234.450 15.600 234.750 16.000 ;
        RECT 235.000 15.600 235.300 16.000 ;
        RECT 235.700 15.600 236.400 16.000 ;
        RECT 236.650 15.600 236.950 16.000 ;
        RECT 237.200 15.600 237.500 16.000 ;
        RECT 237.750 15.700 238.250 16.000 ;
        RECT 238.650 16.000 238.850 17.200 ;
        RECT 239.100 16.400 239.500 16.550 ;
        RECT 240.750 16.400 240.950 17.200 ;
        RECT 242.050 17.000 242.250 17.200 ;
        RECT 241.150 16.800 242.250 17.000 ;
        RECT 241.150 16.600 241.750 16.800 ;
        RECT 239.100 16.200 241.300 16.400 ;
        RECT 240.000 16.000 240.200 16.200 ;
        RECT 241.100 16.000 241.300 16.200 ;
        RECT 241.550 16.000 241.750 16.600 ;
        RECT 242.000 16.400 242.400 16.600 ;
        RECT 242.750 16.400 242.950 17.200 ;
        RECT 243.850 16.400 244.050 17.200 ;
        RECT 245.150 16.700 245.350 17.300 ;
        RECT 245.700 17.200 246.000 17.300 ;
        RECT 246.250 17.200 246.950 17.600 ;
        RECT 247.250 17.200 247.700 17.600 ;
        RECT 247.950 17.200 248.250 17.600 ;
        RECT 248.500 17.200 248.800 17.600 ;
        RECT 249.200 17.200 249.500 17.600 ;
        RECT 249.750 17.200 250.050 17.600 ;
        RECT 250.300 17.200 250.600 17.600 ;
        RECT 252.200 17.500 252.500 17.600 ;
        RECT 251.650 17.300 252.500 17.500 ;
        RECT 242.000 16.200 244.050 16.400 ;
        RECT 244.350 16.500 245.350 16.700 ;
        RECT 244.350 16.300 244.750 16.500 ;
        RECT 243.850 16.000 244.050 16.200 ;
        RECT 238.650 15.700 239.150 16.000 ;
        RECT 237.750 15.600 238.050 15.700 ;
        RECT 238.850 15.600 239.150 15.700 ;
        RECT 239.400 15.600 239.700 16.000 ;
        RECT 239.950 15.600 240.250 16.000 ;
        RECT 240.500 15.600 240.800 16.000 ;
        RECT 241.050 15.600 241.350 16.000 ;
        RECT 241.550 15.800 242.450 16.000 ;
        RECT 242.150 15.600 242.450 15.800 ;
        RECT 242.700 15.600 243.000 16.000 ;
        RECT 243.250 15.600 243.600 16.000 ;
        RECT 243.800 15.600 244.100 16.000 ;
        RECT 211.600 15.400 211.800 15.600 ;
        RECT 211.500 15.000 211.900 15.400 ;
        RECT 212.600 14.850 212.800 15.600 ;
        RECT 213.700 14.850 213.900 15.600 ;
        RECT 216.050 14.850 216.250 15.600 ;
        RECT 216.450 15.100 216.850 15.500 ;
        RECT 217.200 15.400 217.400 15.600 ;
        RECT 217.100 15.050 217.500 15.400 ;
        RECT 217.750 14.850 217.950 15.600 ;
        RECT 218.850 14.850 219.050 15.600 ;
        RECT 221.050 14.850 221.250 15.600 ;
        RECT 221.800 15.050 222.200 15.400 ;
        RECT 223.350 15.150 223.650 15.550 ;
        RECT 223.400 14.850 223.600 15.150 ;
        RECT 224.650 14.850 224.850 15.600 ;
        RECT 225.750 14.850 225.950 15.600 ;
        RECT 228.100 14.850 228.300 15.600 ;
        RECT 229.800 15.050 230.200 15.400 ;
        RECT 230.400 14.850 230.600 15.600 ;
        RECT 232.150 14.850 232.350 15.600 ;
        RECT 233.400 14.850 233.600 15.600 ;
        RECT 234.500 14.850 234.700 15.600 ;
        RECT 236.150 14.850 236.350 15.600 ;
        RECT 239.450 14.850 239.650 15.600 ;
        RECT 240.550 14.850 240.750 15.600 ;
        RECT 242.870 15.000 243.200 15.400 ;
        RECT 243.400 14.850 243.600 15.600 ;
        RECT 245.150 15.550 245.350 16.500 ;
        RECT 245.600 15.950 246.000 16.150 ;
        RECT 247.250 15.950 247.450 17.200 ;
        RECT 248.550 17.000 248.750 17.200 ;
        RECT 247.650 16.800 248.750 17.000 ;
        RECT 247.650 16.600 248.250 16.800 ;
        RECT 245.600 15.750 247.800 15.950 ;
        RECT 246.500 15.550 246.700 15.750 ;
        RECT 247.600 15.550 247.800 15.750 ;
        RECT 248.050 15.550 248.250 16.600 ;
        RECT 248.500 15.950 248.900 16.150 ;
        RECT 249.250 15.950 249.450 17.200 ;
        RECT 250.350 15.950 250.550 17.200 ;
        RECT 251.650 16.700 251.850 17.300 ;
        RECT 252.200 17.200 252.500 17.300 ;
        RECT 252.750 17.200 253.450 17.600 ;
        RECT 253.750 17.200 254.200 17.600 ;
        RECT 254.450 17.200 254.750 17.600 ;
        RECT 255.000 17.200 255.300 17.600 ;
        RECT 255.700 17.200 256.000 17.600 ;
        RECT 256.250 17.200 256.550 17.600 ;
        RECT 256.800 17.200 257.100 17.600 ;
        RECT 258.700 17.500 259.000 17.600 ;
        RECT 258.150 17.300 259.000 17.500 ;
        RECT 250.850 16.500 251.850 16.700 ;
        RECT 250.850 16.300 251.250 16.500 ;
        RECT 248.500 15.750 250.550 15.950 ;
        RECT 250.350 15.550 250.550 15.750 ;
        RECT 251.650 15.550 251.850 16.500 ;
        RECT 252.100 15.950 252.500 16.150 ;
        RECT 253.750 15.950 253.950 17.200 ;
        RECT 255.050 17.000 255.250 17.200 ;
        RECT 254.150 16.800 255.250 17.000 ;
        RECT 254.150 16.600 254.750 16.800 ;
        RECT 252.100 15.750 254.300 15.950 ;
        RECT 253.000 15.550 253.200 15.750 ;
        RECT 254.100 15.550 254.300 15.750 ;
        RECT 254.550 15.550 254.750 16.600 ;
        RECT 255.000 15.950 255.400 16.150 ;
        RECT 255.750 15.950 255.950 17.200 ;
        RECT 256.850 15.950 257.050 17.200 ;
        RECT 258.150 16.700 258.350 17.300 ;
        RECT 258.700 17.200 259.000 17.300 ;
        RECT 259.250 17.200 259.950 17.600 ;
        RECT 260.250 17.200 260.700 17.600 ;
        RECT 260.950 17.200 261.250 17.600 ;
        RECT 261.500 17.200 261.800 17.600 ;
        RECT 262.200 17.200 262.500 17.600 ;
        RECT 262.750 17.200 263.050 17.600 ;
        RECT 263.300 17.200 263.600 17.600 ;
        RECT 257.350 16.500 258.350 16.700 ;
        RECT 257.350 16.300 257.750 16.500 ;
        RECT 255.000 15.750 257.050 15.950 ;
        RECT 256.850 15.550 257.050 15.750 ;
        RECT 258.150 15.550 258.350 16.500 ;
        RECT 258.600 15.950 259.000 16.150 ;
        RECT 260.250 15.950 260.450 17.200 ;
        RECT 261.550 17.000 261.750 17.200 ;
        RECT 260.650 16.800 261.750 17.000 ;
        RECT 260.650 16.600 261.250 16.800 ;
        RECT 258.600 15.750 260.800 15.950 ;
        RECT 259.500 15.550 259.700 15.750 ;
        RECT 260.600 15.550 260.800 15.750 ;
        RECT 261.050 15.550 261.250 16.600 ;
        RECT 261.500 15.950 261.900 16.150 ;
        RECT 262.250 15.950 262.450 17.200 ;
        RECT 263.350 15.950 263.550 17.200 ;
        RECT 263.760 16.300 264.050 16.700 ;
        RECT 261.500 15.750 263.550 15.950 ;
        RECT 263.350 15.550 263.550 15.750 ;
        RECT 244.650 15.150 244.950 15.550 ;
        RECT 245.150 15.250 245.650 15.550 ;
        RECT 245.350 15.150 245.650 15.250 ;
        RECT 245.900 15.150 246.200 15.550 ;
        RECT 246.450 15.150 246.750 15.550 ;
        RECT 247.000 15.150 247.300 15.550 ;
        RECT 247.550 15.150 247.850 15.550 ;
        RECT 248.050 15.350 248.950 15.550 ;
        RECT 248.650 15.150 248.950 15.350 ;
        RECT 249.200 15.150 249.500 15.550 ;
        RECT 249.750 15.150 250.050 15.550 ;
        RECT 250.300 15.150 250.600 15.550 ;
        RECT 251.150 15.150 251.450 15.550 ;
        RECT 251.650 15.250 252.150 15.550 ;
        RECT 251.850 15.150 252.150 15.250 ;
        RECT 252.400 15.150 252.700 15.550 ;
        RECT 252.950 15.150 253.250 15.550 ;
        RECT 253.500 15.150 253.800 15.550 ;
        RECT 254.050 15.150 254.350 15.550 ;
        RECT 254.550 15.350 255.450 15.550 ;
        RECT 255.150 15.150 255.450 15.350 ;
        RECT 255.700 15.150 256.000 15.550 ;
        RECT 256.250 15.150 256.550 15.550 ;
        RECT 256.800 15.150 257.100 15.550 ;
        RECT 257.650 15.150 257.950 15.550 ;
        RECT 258.150 15.250 258.650 15.550 ;
        RECT 258.350 15.150 258.650 15.250 ;
        RECT 258.900 15.150 259.200 15.550 ;
        RECT 259.450 15.150 259.750 15.550 ;
        RECT 260.000 15.150 260.300 15.550 ;
        RECT 260.550 15.150 260.850 15.550 ;
        RECT 261.050 15.350 261.950 15.550 ;
        RECT 261.650 15.150 261.950 15.350 ;
        RECT 262.200 15.150 262.500 15.550 ;
        RECT 262.750 15.150 263.050 15.550 ;
        RECT 263.300 15.150 263.600 15.550 ;
        RECT 244.700 14.850 244.900 15.150 ;
        RECT 245.950 14.850 246.150 15.150 ;
        RECT 247.050 14.850 247.250 15.150 ;
        RECT 249.800 14.850 250.000 15.150 ;
        RECT 251.200 14.850 251.400 15.150 ;
        RECT 252.450 14.850 252.650 15.150 ;
        RECT 253.550 14.850 253.750 15.150 ;
        RECT 256.300 14.850 256.500 15.150 ;
        RECT 257.700 14.850 257.900 15.150 ;
        RECT 258.950 14.850 259.150 15.150 ;
        RECT 260.050 14.850 260.250 15.150 ;
        RECT 262.800 14.850 263.000 15.150 ;
        RECT 212.500 14.450 212.900 14.850 ;
        RECT 213.600 14.450 214.000 14.850 ;
        RECT 215.950 14.450 216.350 14.850 ;
        RECT 217.650 14.450 218.050 14.850 ;
        RECT 218.750 14.450 219.150 14.850 ;
        RECT 220.950 14.450 221.350 14.850 ;
        RECT 223.300 14.450 223.700 14.850 ;
        RECT 224.550 14.450 224.950 14.850 ;
        RECT 225.650 14.450 226.050 14.850 ;
        RECT 228.000 14.450 228.400 14.850 ;
        RECT 230.300 14.450 230.700 14.850 ;
        RECT 232.050 14.450 232.450 14.850 ;
        RECT 233.300 14.450 233.700 14.850 ;
        RECT 234.400 14.450 234.800 14.850 ;
        RECT 236.050 14.450 236.450 14.850 ;
        RECT 239.350 14.450 239.750 14.850 ;
        RECT 240.450 14.450 240.850 14.850 ;
        RECT 243.300 14.450 243.700 14.850 ;
        RECT 244.600 14.450 245.000 14.850 ;
        RECT 245.850 14.450 246.250 14.850 ;
        RECT 246.950 14.450 247.350 14.850 ;
        RECT 249.700 14.450 250.100 14.850 ;
        RECT 251.100 14.450 251.500 14.850 ;
        RECT 252.350 14.450 252.750 14.850 ;
        RECT 253.450 14.450 253.850 14.850 ;
        RECT 256.200 14.450 256.600 14.850 ;
        RECT 257.600 14.450 258.000 14.850 ;
        RECT 258.850 14.450 259.250 14.850 ;
        RECT 259.950 14.450 260.350 14.850 ;
        RECT 262.700 14.450 263.100 14.850 ;
      LAYER met1 ;
        RECT 213.300 18.350 213.700 18.750 ;
        RECT 215.400 18.350 215.800 18.750 ;
        RECT 218.750 18.350 219.150 18.750 ;
        RECT 221.600 18.350 222.000 18.750 ;
        RECT 225.350 18.350 225.750 18.750 ;
        RECT 227.500 18.350 227.900 18.750 ;
        RECT 229.700 18.350 230.100 18.750 ;
        RECT 230.950 18.350 231.350 18.750 ;
        RECT 232.050 18.350 232.450 18.750 ;
        RECT 234.400 18.350 234.800 18.750 ;
        RECT 236.600 18.350 237.000 18.750 ;
        RECT 239.700 18.350 240.100 18.750 ;
        RECT 241.400 18.350 241.800 18.750 ;
        RECT 243.200 18.350 243.600 18.750 ;
        RECT 246.200 18.350 246.600 18.750 ;
        RECT 247.900 18.350 248.300 18.750 ;
        RECT 249.700 18.350 250.100 18.750 ;
        RECT 252.700 18.350 253.100 18.750 ;
        RECT 254.400 18.350 254.800 18.750 ;
        RECT 256.200 18.350 256.600 18.750 ;
        RECT 259.200 18.350 259.600 18.750 ;
        RECT 260.900 18.350 261.300 18.750 ;
        RECT 262.700 18.350 263.100 18.750 ;
        RECT 214.900 18.000 215.300 18.200 ;
        RECT 215.900 18.000 216.250 18.200 ;
        RECT 214.900 17.800 216.250 18.000 ;
        RECT 216.450 18.000 216.850 18.100 ;
        RECT 220.500 18.000 220.900 18.200 ;
        RECT 216.450 17.800 220.900 18.000 ;
        RECT 221.200 18.000 221.500 18.200 ;
        RECT 227.000 18.000 227.400 18.200 ;
        RECT 228.100 18.000 228.500 18.200 ;
        RECT 221.200 17.800 223.850 18.000 ;
        RECT 227.000 17.800 228.500 18.000 ;
        RECT 233.750 18.050 234.150 18.200 ;
        RECT 235.800 18.050 236.200 18.200 ;
        RECT 233.750 17.850 236.200 18.050 ;
        RECT 245.550 18.000 245.950 18.200 ;
        RECT 248.450 18.000 248.850 18.200 ;
        RECT 245.550 17.800 248.850 18.000 ;
        RECT 252.050 18.000 252.450 18.200 ;
        RECT 254.950 18.000 255.350 18.200 ;
        RECT 252.050 17.800 255.350 18.000 ;
        RECT 258.550 18.000 258.950 18.200 ;
        RECT 261.450 18.000 261.850 18.200 ;
        RECT 258.550 17.800 261.850 18.000 ;
        RECT 216.450 17.700 216.850 17.800 ;
        RECT 223.650 17.600 223.850 17.800 ;
        RECT 245.750 17.600 245.950 17.800 ;
        RECT 252.250 17.600 252.450 17.800 ;
        RECT 258.750 17.600 258.950 17.800 ;
        RECT 223.650 17.200 224.050 17.600 ;
        RECT 211.200 16.350 211.600 16.750 ;
        RECT 219.750 16.350 222.750 16.550 ;
        RECT 219.750 16.200 220.150 16.350 ;
        RECT 222.350 16.200 222.750 16.350 ;
        RECT 231.150 16.250 231.550 16.650 ;
        RECT 263.760 16.300 264.050 16.700 ;
        RECT 211.500 15.300 211.900 15.400 ;
        RECT 216.450 15.300 216.850 15.500 ;
        RECT 231.150 15.400 231.350 16.250 ;
        RECT 211.500 15.100 216.850 15.300 ;
        RECT 217.100 15.250 217.500 15.400 ;
        RECT 221.800 15.250 222.200 15.400 ;
        RECT 229.800 15.250 230.200 15.400 ;
        RECT 211.500 15.000 211.900 15.100 ;
        RECT 217.100 15.050 230.200 15.250 ;
        RECT 231.150 15.200 243.200 15.400 ;
        RECT 242.870 15.000 243.200 15.200 ;
        RECT 212.500 14.450 212.900 14.850 ;
        RECT 213.600 14.450 214.000 14.850 ;
        RECT 215.950 14.450 216.350 14.850 ;
        RECT 217.650 14.450 218.050 14.850 ;
        RECT 218.750 14.450 219.150 14.850 ;
        RECT 220.950 14.450 221.350 14.850 ;
        RECT 223.300 14.450 223.700 14.850 ;
        RECT 224.550 14.450 224.950 14.850 ;
        RECT 225.650 14.450 226.050 14.850 ;
        RECT 228.000 14.450 228.400 14.850 ;
        RECT 230.300 14.450 230.700 14.850 ;
        RECT 232.050 14.450 232.450 14.850 ;
        RECT 233.300 14.450 233.700 14.850 ;
        RECT 234.400 14.450 234.800 14.850 ;
        RECT 236.050 14.450 236.450 14.850 ;
        RECT 239.350 14.450 239.750 14.850 ;
        RECT 240.450 14.450 240.850 14.850 ;
        RECT 243.300 14.450 243.700 14.850 ;
        RECT 244.600 14.450 245.000 14.850 ;
        RECT 245.850 14.450 246.250 14.850 ;
        RECT 246.950 14.450 247.350 14.850 ;
        RECT 249.700 14.450 250.100 14.850 ;
        RECT 251.100 14.450 251.500 14.850 ;
        RECT 252.350 14.450 252.750 14.850 ;
        RECT 253.450 14.450 253.850 14.850 ;
        RECT 256.200 14.450 256.600 14.850 ;
        RECT 257.600 14.450 258.000 14.850 ;
        RECT 258.850 14.450 259.250 14.850 ;
        RECT 259.950 14.450 260.350 14.850 ;
        RECT 262.700 14.450 263.100 14.850 ;
      LAYER met2 ;
        RECT 211.300 18.350 263.100 18.750 ;
        RECT 210.650 16.350 211.600 16.750 ;
        RECT 263.760 16.300 264.050 16.700 ;
        RECT 211.300 14.450 263.100 14.850 ;
  END
END divide_by_120
END LIBRARY

